* NGSPICE file created from ExperiarCore.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

.subckt ExperiarCore addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6]
+ addr0[7] addr0[8] addr1[0] addr1[1] addr1[2] addr1[3] addr1[4] addr1[5] addr1[6]
+ addr1[7] addr1[8] clk0 clk1 coreIndex[0] coreIndex[1] coreIndex[2] coreIndex[3]
+ coreIndex[4] coreIndex[5] coreIndex[6] coreIndex[7] core_wb_ack_i core_wb_adr_o[0]
+ core_wb_adr_o[10] core_wb_adr_o[11] core_wb_adr_o[12] core_wb_adr_o[13] core_wb_adr_o[14]
+ core_wb_adr_o[15] core_wb_adr_o[16] core_wb_adr_o[17] core_wb_adr_o[18] core_wb_adr_o[19]
+ core_wb_adr_o[1] core_wb_adr_o[20] core_wb_adr_o[21] core_wb_adr_o[22] core_wb_adr_o[23]
+ core_wb_adr_o[24] core_wb_adr_o[25] core_wb_adr_o[26] core_wb_adr_o[27] core_wb_adr_o[2]
+ core_wb_adr_o[3] core_wb_adr_o[4] core_wb_adr_o[5] core_wb_adr_o[6] core_wb_adr_o[7]
+ core_wb_adr_o[8] core_wb_adr_o[9] core_wb_cyc_o core_wb_data_i[0] core_wb_data_i[10]
+ core_wb_data_i[11] core_wb_data_i[12] core_wb_data_i[13] core_wb_data_i[14] core_wb_data_i[15]
+ core_wb_data_i[16] core_wb_data_i[17] core_wb_data_i[18] core_wb_data_i[19] core_wb_data_i[1]
+ core_wb_data_i[20] core_wb_data_i[21] core_wb_data_i[22] core_wb_data_i[23] core_wb_data_i[24]
+ core_wb_data_i[25] core_wb_data_i[26] core_wb_data_i[27] core_wb_data_i[28] core_wb_data_i[29]
+ core_wb_data_i[2] core_wb_data_i[30] core_wb_data_i[31] core_wb_data_i[3] core_wb_data_i[4]
+ core_wb_data_i[5] core_wb_data_i[6] core_wb_data_i[7] core_wb_data_i[8] core_wb_data_i[9]
+ core_wb_data_o[0] core_wb_data_o[10] core_wb_data_o[11] core_wb_data_o[12] core_wb_data_o[13]
+ core_wb_data_o[14] core_wb_data_o[15] core_wb_data_o[16] core_wb_data_o[17] core_wb_data_o[18]
+ core_wb_data_o[19] core_wb_data_o[1] core_wb_data_o[20] core_wb_data_o[21] core_wb_data_o[22]
+ core_wb_data_o[23] core_wb_data_o[24] core_wb_data_o[25] core_wb_data_o[26] core_wb_data_o[27]
+ core_wb_data_o[28] core_wb_data_o[29] core_wb_data_o[2] core_wb_data_o[30] core_wb_data_o[31]
+ core_wb_data_o[3] core_wb_data_o[4] core_wb_data_o[5] core_wb_data_o[6] core_wb_data_o[7]
+ core_wb_data_o[8] core_wb_data_o[9] core_wb_error_i core_wb_sel_o[0] core_wb_sel_o[1]
+ core_wb_sel_o[2] core_wb_sel_o[3] core_wb_stall_i core_wb_stb_o core_wb_we_o csb0[0]
+ csb0[1] csb1[0] csb1[1] din0[0] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15]
+ din0[16] din0[17] din0[18] din0[19] din0[1] din0[20] din0[21] din0[22] din0[23]
+ din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[2] din0[30] din0[31]
+ din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] dout0[0] dout0[10] dout0[11]
+ dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19]
+ dout0[1] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27]
+ dout0[28] dout0[29] dout0[2] dout0[30] dout0[31] dout0[32] dout0[33] dout0[34] dout0[35]
+ dout0[36] dout0[37] dout0[38] dout0[39] dout0[3] dout0[40] dout0[41] dout0[42] dout0[43]
+ dout0[44] dout0[45] dout0[46] dout0[47] dout0[48] dout0[49] dout0[4] dout0[50] dout0[51]
+ dout0[52] dout0[53] dout0[54] dout0[55] dout0[56] dout0[57] dout0[58] dout0[59]
+ dout0[5] dout0[60] dout0[61] dout0[62] dout0[63] dout0[6] dout0[7] dout0[8] dout0[9]
+ dout1[0] dout1[10] dout1[11] dout1[12] dout1[13] dout1[14] dout1[15] dout1[16] dout1[17]
+ dout1[18] dout1[19] dout1[1] dout1[20] dout1[21] dout1[22] dout1[23] dout1[24] dout1[25]
+ dout1[26] dout1[27] dout1[28] dout1[29] dout1[2] dout1[30] dout1[31] dout1[32] dout1[33]
+ dout1[34] dout1[35] dout1[36] dout1[37] dout1[38] dout1[39] dout1[3] dout1[40] dout1[41]
+ dout1[42] dout1[43] dout1[44] dout1[45] dout1[46] dout1[47] dout1[48] dout1[49]
+ dout1[4] dout1[50] dout1[51] dout1[52] dout1[53] dout1[54] dout1[55] dout1[56] dout1[57]
+ dout1[58] dout1[59] dout1[5] dout1[60] dout1[61] dout1[62] dout1[63] dout1[6] dout1[7]
+ dout1[8] dout1[9] irq[0] irq[10] irq[11] irq[12] irq[13] irq[14] irq[15] irq[1]
+ irq[2] irq[3] irq[4] irq[5] irq[6] irq[7] irq[8] irq[9] jtag_tck jtag_tdi jtag_tdo
+ jtag_tms localMemory_wb_ack_o localMemory_wb_adr_i[0] localMemory_wb_adr_i[10] localMemory_wb_adr_i[11]
+ localMemory_wb_adr_i[12] localMemory_wb_adr_i[13] localMemory_wb_adr_i[14] localMemory_wb_adr_i[15]
+ localMemory_wb_adr_i[16] localMemory_wb_adr_i[17] localMemory_wb_adr_i[18] localMemory_wb_adr_i[19]
+ localMemory_wb_adr_i[1] localMemory_wb_adr_i[20] localMemory_wb_adr_i[21] localMemory_wb_adr_i[22]
+ localMemory_wb_adr_i[23] localMemory_wb_adr_i[2] localMemory_wb_adr_i[3] localMemory_wb_adr_i[4]
+ localMemory_wb_adr_i[5] localMemory_wb_adr_i[6] localMemory_wb_adr_i[7] localMemory_wb_adr_i[8]
+ localMemory_wb_adr_i[9] localMemory_wb_cyc_i localMemory_wb_data_i[0] localMemory_wb_data_i[10]
+ localMemory_wb_data_i[11] localMemory_wb_data_i[12] localMemory_wb_data_i[13] localMemory_wb_data_i[14]
+ localMemory_wb_data_i[15] localMemory_wb_data_i[16] localMemory_wb_data_i[17] localMemory_wb_data_i[18]
+ localMemory_wb_data_i[19] localMemory_wb_data_i[1] localMemory_wb_data_i[20] localMemory_wb_data_i[21]
+ localMemory_wb_data_i[22] localMemory_wb_data_i[23] localMemory_wb_data_i[24] localMemory_wb_data_i[25]
+ localMemory_wb_data_i[26] localMemory_wb_data_i[27] localMemory_wb_data_i[28] localMemory_wb_data_i[29]
+ localMemory_wb_data_i[2] localMemory_wb_data_i[30] localMemory_wb_data_i[31] localMemory_wb_data_i[3]
+ localMemory_wb_data_i[4] localMemory_wb_data_i[5] localMemory_wb_data_i[6] localMemory_wb_data_i[7]
+ localMemory_wb_data_i[8] localMemory_wb_data_i[9] localMemory_wb_data_o[0] localMemory_wb_data_o[10]
+ localMemory_wb_data_o[11] localMemory_wb_data_o[12] localMemory_wb_data_o[13] localMemory_wb_data_o[14]
+ localMemory_wb_data_o[15] localMemory_wb_data_o[16] localMemory_wb_data_o[17] localMemory_wb_data_o[18]
+ localMemory_wb_data_o[19] localMemory_wb_data_o[1] localMemory_wb_data_o[20] localMemory_wb_data_o[21]
+ localMemory_wb_data_o[22] localMemory_wb_data_o[23] localMemory_wb_data_o[24] localMemory_wb_data_o[25]
+ localMemory_wb_data_o[26] localMemory_wb_data_o[27] localMemory_wb_data_o[28] localMemory_wb_data_o[29]
+ localMemory_wb_data_o[2] localMemory_wb_data_o[30] localMemory_wb_data_o[31] localMemory_wb_data_o[3]
+ localMemory_wb_data_o[4] localMemory_wb_data_o[5] localMemory_wb_data_o[6] localMemory_wb_data_o[7]
+ localMemory_wb_data_o[8] localMemory_wb_data_o[9] localMemory_wb_error_o localMemory_wb_sel_i[0]
+ localMemory_wb_sel_i[1] localMemory_wb_sel_i[2] localMemory_wb_sel_i[3] localMemory_wb_stall_o
+ localMemory_wb_stb_i localMemory_wb_we_i manufacturerID[0] manufacturerID[10] manufacturerID[1]
+ manufacturerID[2] manufacturerID[3] manufacturerID[4] manufacturerID[5] manufacturerID[6]
+ manufacturerID[7] manufacturerID[8] manufacturerID[9] partID[0] partID[10] partID[11]
+ partID[12] partID[13] partID[14] partID[15] partID[1] partID[2] partID[3] partID[4]
+ partID[5] partID[6] partID[7] partID[8] partID[9] probe_env[0] probe_env[1] probe_errorCode[0]
+ probe_errorCode[1] probe_isBranch probe_isCompressed probe_isLoad probe_isStore
+ probe_jtagInstruction[0] probe_jtagInstruction[1] probe_jtagInstruction[2] probe_jtagInstruction[3]
+ probe_jtagInstruction[4] probe_opcode[0] probe_opcode[1] probe_opcode[2] probe_opcode[3]
+ probe_opcode[4] probe_opcode[5] probe_opcode[6] probe_programCounter[0] probe_programCounter[10]
+ probe_programCounter[11] probe_programCounter[12] probe_programCounter[13] probe_programCounter[14]
+ probe_programCounter[15] probe_programCounter[16] probe_programCounter[17] probe_programCounter[18]
+ probe_programCounter[19] probe_programCounter[1] probe_programCounter[20] probe_programCounter[21]
+ probe_programCounter[22] probe_programCounter[23] probe_programCounter[24] probe_programCounter[25]
+ probe_programCounter[26] probe_programCounter[27] probe_programCounter[28] probe_programCounter[29]
+ probe_programCounter[2] probe_programCounter[30] probe_programCounter[31] probe_programCounter[3]
+ probe_programCounter[4] probe_programCounter[5] probe_programCounter[6] probe_programCounter[7]
+ probe_programCounter[8] probe_programCounter[9] probe_state[0] probe_state[1] probe_takeBranch
+ vccd1 versionID[0] versionID[1] versionID[2] versionID[3] vssd1 wb_clk_i wb_rst_i
+ web0 wmask0[0] wmask0[1] wmask0[2] wmask0[3]
XFILLER_246_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18869_ _23139_/Q _18868_/X _18872_/S vssd1 vssd1 vccd1 vccd1 _18870_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20900_ _21317_/A _20894_/X _20779_/B _20897_/X vssd1 vssd1 vccd1 vccd1 _20900_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_255_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21880_ _21613_/X _21879_/Y _21683_/A _23799_/Q vssd1 vssd1 vccd1 vccd1 _21880_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_227_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20831_ _20843_/A _20831_/B vssd1 vssd1 vccd1 vccd1 _20832_/A sky130_fd_sc_hd__and2_1
XFILLER_70_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23550_ _23550_/CLK _23550_/D vssd1 vssd1 vccd1 vccd1 _23550_/Q sky130_fd_sc_hd__dfxtp_1
X_20762_ _20768_/A _20762_/B _20762_/C vssd1 vssd1 vccd1 vccd1 _20762_/X sky130_fd_sc_hd__or3_1
XFILLER_306_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_260 _17172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_271 _18827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_282 _15910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22501_ _23704_/CLK _22501_/D vssd1 vssd1 vccd1 vccd1 _22501_/Q sky130_fd_sc_hd__dfxtp_4
X_23481_ _23548_/CLK _23481_/D vssd1 vssd1 vccd1 vccd1 _23481_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_250_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_293 _18852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20693_ _11483_/X _20692_/X _20649_/X vssd1 vssd1 vccd1 vccd1 _20693_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_338_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22432_ _23503_/CLK _22432_/D vssd1 vssd1 vccd1 vccd1 _22432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_309_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_353_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22363_ _23563_/CLK _22363_/D vssd1 vssd1 vccd1 vccd1 _22363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_352_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_337_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21314_ _23782_/Q _21814_/B _21313_/X vssd1 vssd1 vccd1 vccd1 _21314_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_352_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22294_ _23558_/CLK _22294_/D vssd1 vssd1 vccd1 vccd1 _22294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_324_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_352_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_324_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21245_ _17149_/A _21242_/X _21244_/Y _21236_/X vssd1 vssd1 vccd1 vccd1 _23894_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_151_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_305_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21176_ _23873_/Q _21147_/X _21173_/Y _21174_/X _21175_/X vssd1 vssd1 vccd1 vccd1
+ _23873_/D sky130_fd_sc_hd__o221a_1
XFILLER_278_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_321_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_321_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20127_ _20137_/A _20127_/B _20127_/C vssd1 vssd1 vccd1 vccd1 _23648_/D sky130_fd_sc_hd__nor3_1
XFILLER_293_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20058_ _20067_/A vssd1 vssd1 vccd1 vccd1 _20058_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_133_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_292_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ _23309_/Q _23277_/Q _23245_/Q _23533_/Q _12070_/S _11163_/A vssd1 vssd1 vccd1
+ vccd1 _11901_/B sky130_fd_sc_hd__mux4_2
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ _12700_/X _12871_/Y _12875_/Y _12877_/Y _12879_/Y vssd1 vssd1 vccd1 vccd1
+ _12880_/X sky130_fd_sc_hd__o32a_1
XFILLER_234_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23817_ _23818_/CLK _23817_/D vssd1 vssd1 vccd1 vccd1 _23817_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _22366_/Q _22398_/Q _22687_/Q _23054_/Q _11719_/A _12246_/A vssd1 vssd1 vccd1
+ vccd1 _11832_/B sky130_fd_sc_hd__mux4_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _14550_/A _14550_/B _14550_/C vssd1 vssd1 vccd1 vccd1 _14551_/C sky130_fd_sc_hd__or3_1
XFILLER_198_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11762_ _23922_/Q vssd1 vssd1 vccd1 vccd1 _21652_/A sky130_fd_sc_hd__inv_4
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23748_ _23866_/CLK _23748_/D vssd1 vssd1 vccd1 vccd1 _23748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13501_/A vssd1 vssd1 vccd1 vccd1 _13621_/A sky130_fd_sc_hd__inv_2
XFILLER_199_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _15595_/A vssd1 vssd1 vccd1 vccd1 _15215_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_202_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11693_ _12523_/A vssd1 vssd1 vccd1 vccd1 _12196_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23679_ _23684_/CLK _23679_/D vssd1 vssd1 vccd1 vccd1 _23679_/Q sky130_fd_sc_hd__dfxtp_1
X_16220_ _18785_/A vssd1 vssd1 vccd1 vccd1 _16220_/X sky130_fd_sc_hd__buf_2
X_13432_ _13432_/A _13432_/B vssd1 vssd1 vccd1 vccd1 _13433_/A sky130_fd_sc_hd__and2_2
XFILLER_329_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16151_ _22216_/A _22219_/A _16151_/C vssd1 vssd1 vccd1 vccd1 _16165_/B sky130_fd_sc_hd__and3_2
XFILLER_344_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13363_ _13464_/B _13363_/B vssd1 vssd1 vccd1 vccd1 _13367_/C sky130_fd_sc_hd__nor2_8
XFILLER_343_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_315_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15102_ _12283_/X _15048_/X _15100_/X _21500_/B _15041_/X vssd1 vssd1 vccd1 vccd1
+ _18792_/A sky130_fd_sc_hd__a32o_4
XFILLER_355_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12314_ _12324_/A vssd1 vssd1 vccd1 vccd1 _12314_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16082_ _21550_/A vssd1 vssd1 vccd1 vccd1 _21605_/A sky130_fd_sc_hd__buf_8
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13294_ _13287_/Y _13289_/Y _13291_/Y _13293_/Y _11483_/A vssd1 vssd1 vccd1 vccd1
+ _13295_/C sky130_fd_sc_hd__o221a_1
XFILLER_331_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15033_ input137/X input162/X _15033_/S vssd1 vssd1 vccd1 vccd1 _15033_/X sky130_fd_sc_hd__mux2_8
X_19910_ _19910_/A vssd1 vssd1 vccd1 vccd1 _23586_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12245_ _22299_/Q _23435_/Q _12245_/S vssd1 vssd1 vccd1 vccd1 _12246_/B sky130_fd_sc_hd__mux2_1
XFILLER_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19841_ _23556_/Q _19264_/A _19841_/S vssd1 vssd1 vccd1 vccd1 _19842_/A sky130_fd_sc_hd__mux2_1
X_12176_ _12291_/A _12176_/B vssd1 vssd1 vccd1 vccd1 _12176_/Y sky130_fd_sc_hd__nor2_1
XFILLER_150_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_311_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11127_ _11127_/A vssd1 vssd1 vccd1 vccd1 _11780_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_324_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16984_ _21294_/B _16984_/B vssd1 vssd1 vccd1 vccd1 _17224_/B sky130_fd_sc_hd__nor2_1
X_19772_ _19828_/A vssd1 vssd1 vccd1 vccd1 _19841_/S sky130_fd_sc_hd__buf_6
XFILLER_296_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_296_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_288_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15935_ _18849_/A vssd1 vssd1 vccd1 vccd1 _19242_/A sky130_fd_sc_hd__clkbuf_4
X_18723_ _18723_/A vssd1 vssd1 vccd1 vccd1 _23087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_324_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23414_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18654_ _23057_/Q _17585_/X _18658_/S vssd1 vssd1 vccd1 vccd1 _18655_/A sky130_fd_sc_hd__mux2_1
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ _15674_/A _15865_/Y _15676_/X vssd1 vssd1 vccd1 vccd1 _15866_/Y sky130_fd_sc_hd__a21oi_2
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17605_ _22696_/Q _17604_/X _17608_/S vssd1 vssd1 vccd1 vccd1 _17606_/A sky130_fd_sc_hd__mux2_1
XFILLER_291_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14817_ _20493_/B vssd1 vssd1 vccd1 vccd1 _16079_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_236_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18585_ _18585_/A vssd1 vssd1 vccd1 vccd1 _23026_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_251_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15797_ _15797_/A _15797_/B vssd1 vssd1 vccd1 vccd1 _15797_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_340_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17536_ _22674_/Q _16297_/X _17538_/S vssd1 vssd1 vccd1 vccd1 _17537_/A sky130_fd_sc_hd__mux2_1
X_14748_ _14748_/A vssd1 vssd1 vccd1 vccd1 _14748_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17467_ _22644_/Q _16303_/X _17469_/S vssd1 vssd1 vccd1 vccd1 _17468_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_339_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14679_ _14836_/A vssd1 vssd1 vccd1 vccd1 _14682_/A sky130_fd_sc_hd__clkbuf_4
X_16418_ _15523_/X _22371_/Q _16418_/S vssd1 vssd1 vccd1 vccd1 _16419_/A sky130_fd_sc_hd__mux2_1
X_19206_ _19206_/A vssd1 vssd1 vccd1 vccd1 _23281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17398_ _19843_/B vssd1 vssd1 vccd1 vccd1 _19164_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_335_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19137_ _19148_/A vssd1 vssd1 vccd1 vccd1 _19146_/S sky130_fd_sc_hd__buf_2
XFILLER_353_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16349_ _15625_/X _22341_/Q _16355_/S vssd1 vssd1 vccd1 vccd1 _16350_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19068_ _19068_/A vssd1 vssd1 vccd1 vccd1 _23226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput401 _14018_/X vssd1 vssd1 vccd1 vccd1 din0[5] sky130_fd_sc_hd__buf_2
XFILLER_334_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18019_ _18098_/A vssd1 vssd1 vccd1 vccd1 _18053_/A sky130_fd_sc_hd__buf_2
Xoutput412 _22566_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[13] sky130_fd_sc_hd__buf_2
XFILLER_218_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput423 _22576_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[23] sky130_fd_sc_hd__buf_2
XFILLER_322_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_350_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput434 _22557_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[4] sky130_fd_sc_hd__buf_2
XFILLER_303_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput445 _13432_/A vssd1 vssd1 vccd1 vccd1 probe_isBranch sky130_fd_sc_hd__buf_2
XFILLER_321_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput456 _23881_/Q vssd1 vssd1 vccd1 vccd1 probe_opcode[2] sky130_fd_sc_hd__buf_2
X_21030_ _21051_/A vssd1 vssd1 vccd1 vccd1 _21048_/B sky130_fd_sc_hd__clkbuf_2
Xoutput467 _23926_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[15] sky130_fd_sc_hd__buf_2
XFILLER_271_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput478 _23936_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[25] sky130_fd_sc_hd__buf_2
Xoutput489 _23917_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[6] sky130_fd_sc_hd__buf_2
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_302_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22981_ _23552_/CLK _22981_/D vssd1 vssd1 vccd1 vccd1 _22981_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_274_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21932_ _21932_/A _21932_/B vssd1 vssd1 vccd1 vccd1 _22038_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21863_ _21379_/X _21855_/X _21862_/X _21984_/A vssd1 vssd1 vccd1 vccd1 _21863_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23602_ _23602_/CLK _23602_/D vssd1 vssd1 vccd1 vccd1 _23602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_270_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20814_ _20814_/A vssd1 vssd1 vccd1 vccd1 _23758_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21794_ _21790_/B _21793_/Y _22171_/B vssd1 vssd1 vccd1 vccd1 _21794_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23533_ _23534_/CLK _23533_/D vssd1 vssd1 vccd1 vccd1 _23533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20745_ _21077_/A _20724_/X _20733_/X vssd1 vssd1 vccd1 vccd1 _20745_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_195_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23464_ _23558_/CLK _23464_/D vssd1 vssd1 vccd1 vccd1 _23464_/Q sky130_fd_sc_hd__dfxtp_4
X_20676_ _17159_/A _20617_/X _20662_/X vssd1 vssd1 vccd1 vccd1 _20676_/X sky130_fd_sc_hd__a21o_1
XFILLER_183_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22415_ _23583_/CLK _22415_/D vssd1 vssd1 vccd1 vccd1 _22415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_311_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23395_ _23555_/CLK _23395_/D vssd1 vssd1 vccd1 vccd1 _23395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_337_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22346_ _23546_/CLK _22346_/D vssd1 vssd1 vccd1 vccd1 _22346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_345_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_313_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22277_ _23541_/CLK _22277_/D vssd1 vssd1 vccd1 vccd1 _22277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12030_ _22371_/Q _22403_/Q _22692_/Q _23059_/Q _12029_/X _12717_/A vssd1 vssd1 vccd1
+ vccd1 _12030_/X sky130_fd_sc_hd__mux4_1
X_21228_ _14541_/X _21202_/X _21227_/Y _21218_/X vssd1 vssd1 vccd1 vccd1 _23888_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21159_ _20708_/A _21158_/X _21142_/X _20520_/A _21135_/X vssd1 vssd1 vccd1 vccd1
+ _21159_/X sky130_fd_sc_hd__a221o_1
XFILLER_278_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13981_ _13981_/A _13985_/B vssd1 vssd1 vccd1 vccd1 _13982_/A sky130_fd_sc_hd__and2_2
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15720_ _12741_/Y _15460_/B _14259_/A _12743_/B vssd1 vssd1 vccd1 vccd1 _15720_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ _23417_/Q _23033_/Q _23385_/Q _23353_/Q _12825_/X _12672_/A vssd1 vssd1 vccd1
+ vccd1 _12932_/X sky130_fd_sc_hd__mux4_2
XFILLER_219_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _23702_/Q _14905_/X _15650_/X vssd1 vssd1 vccd1 vccd1 _15651_/Y sky130_fd_sc_hd__o21ai_4
X_12863_ _12856_/X _12858_/X _12860_/X _12862_/X _11276_/A vssd1 vssd1 vccd1 vccd1
+ _12864_/C sky130_fd_sc_hd__a221o_1
XFILLER_74_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _20160_/A _15068_/C vssd1 vssd1 vccd1 vccd1 _14603_/A sky130_fd_sc_hd__nor2_2
XFILLER_73_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ _18403_/A _18375_/C vssd1 vssd1 vccd1 vccd1 _18370_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _12324_/A vssd1 vssd1 vccd1 vccd1 _11814_/X sky130_fd_sc_hd__buf_8
X_15582_ _15582_/A _15582_/B vssd1 vssd1 vccd1 vccd1 _15582_/Y sky130_fd_sc_hd__nand2_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _22795_/Q _22763_/Q _22664_/Q _22731_/Q _12792_/X _12793_/X vssd1 vssd1 vccd1
+ vccd1 _12795_/B sky130_fd_sc_hd__mux4_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _22584_/Q _17091_/A _17028_/A _17320_/X vssd1 vssd1 vccd1 vccd1 _22584_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _18769_/A vssd1 vssd1 vccd1 vccd1 _19163_/A sky130_fd_sc_hd__buf_2
X_11745_ _11745_/A vssd1 vssd1 vccd1 vccd1 _11745_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_159_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ _17245_/X _17251_/X _17195_/X _17215_/X vssd1 vssd1 vccd1 vccd1 _17252_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_187_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_348_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14464_ _15211_/A vssd1 vssd1 vccd1 vccd1 _14464_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11676_ _11676_/A vssd1 vssd1 vccd1 vccd1 _12844_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_202_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16203_ _16457_/C _16203_/B vssd1 vssd1 vccd1 vccd1 _16310_/A sky130_fd_sc_hd__nand2_1
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13415_ _13410_/A _13410_/B _13410_/C _13410_/D _14343_/S vssd1 vssd1 vccd1 vccd1
+ _13415_/X sky130_fd_sc_hd__o41a_1
X_17183_ _23479_/Q _17113_/X _17114_/X _17181_/X _17182_/Y vssd1 vssd1 vccd1 vccd1
+ _17183_/X sky130_fd_sc_hd__a32o_1
X_14395_ _22897_/Q _14394_/X _14164_/X _22590_/Q vssd1 vssd1 vccd1 vccd1 _16936_/C
+ sky130_fd_sc_hd__a22o_4
XFILLER_128_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16134_ _22944_/Q _14509_/A _14513_/A _22976_/Q vssd1 vssd1 vccd1 vccd1 _16134_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_343_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13346_ _12162_/Y _13345_/X _12167_/Y vssd1 vssd1 vccd1 vccd1 _13351_/B sky130_fd_sc_hd__a21bo_1
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_317_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_332_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16065_ _23809_/Q _14742_/X _14606_/A vssd1 vssd1 vccd1 vccd1 _16065_/X sky130_fd_sc_hd__a21o_1
XFILLER_331_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13277_ _23329_/Q _23297_/Q _23265_/Q _23553_/Q _13275_/X _13276_/X vssd1 vssd1 vccd1
+ vccd1 _13278_/B sky130_fd_sc_hd__mux4_2
XFILLER_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15016_ _14658_/X _14636_/X _15133_/A vssd1 vssd1 vccd1 vccd1 _15456_/B sky130_fd_sc_hd__mux2_2
X_12228_ _12221_/X _12223_/X _12225_/X _12227_/X _11272_/A vssd1 vssd1 vccd1 vccd1
+ _12229_/C sky130_fd_sc_hd__a221o_1
XFILLER_300_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19824_ _23548_/Q _19239_/A _19826_/S vssd1 vssd1 vccd1 vccd1 _19825_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12159_ _12159_/A _12163_/A vssd1 vssd1 vccd1 vccd1 _13497_/A sky130_fd_sc_hd__nor2_2
XFILLER_111_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_300_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19755_ _19755_/A vssd1 vssd1 vccd1 vccd1 _23517_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16967_ _17262_/A vssd1 vssd1 vccd1 vccd1 _16996_/A sky130_fd_sc_hd__buf_2
XFILLER_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18706_ _16825_/X _23080_/Q _18708_/S vssd1 vssd1 vccd1 vccd1 _18707_/A sky130_fd_sc_hd__mux2_1
XFILLER_265_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15918_ _13399_/Y _13581_/B _15918_/S vssd1 vssd1 vccd1 vccd1 _15918_/X sky130_fd_sc_hd__mux2_1
X_16898_ _16898_/A vssd1 vssd1 vccd1 vccd1 _22546_/D sky130_fd_sc_hd__clkbuf_1
X_19686_ _19686_/A vssd1 vssd1 vccd1 vccd1 _23486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15849_ _13015_/B _15996_/B _15082_/X _13015_/A vssd1 vssd1 vccd1 vccd1 _15849_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_18637_ _18637_/A vssd1 vssd1 vccd1 vccd1 _23049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_280_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18568_ _18568_/A vssd1 vssd1 vccd1 vccd1 _23018_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_339_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17519_ _22666_/Q _16271_/X _17527_/S vssd1 vssd1 vccd1 vccd1 _17520_/A sky130_fd_sc_hd__mux2_1
XFILLER_342_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18499_ _18494_/X _18498_/Y _18490_/X vssd1 vssd1 vccd1 vccd1 _22994_/D sky130_fd_sc_hd__a21oi_1
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_339_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20530_ _21285_/A _20530_/B vssd1 vssd1 vccd1 vccd1 _20536_/B sky130_fd_sc_hd__nor2_2
XFILLER_220_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_327_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_308_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20461_ _21149_/A _20463_/B vssd1 vssd1 vccd1 vccd1 _20461_/Y sky130_fd_sc_hd__nand2_1
XFILLER_229_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22200_ _22193_/A _21366_/X _22199_/Y _22122_/X vssd1 vssd1 vccd1 vccd1 _23940_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_335_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23180_ _23950_/A _23180_/D vssd1 vssd1 vccd1 vccd1 _23180_/Q sky130_fd_sc_hd__dfxtp_1
X_20392_ _20445_/A vssd1 vssd1 vccd1 vccd1 _20392_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_173_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_350_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22131_ _22129_/X _22130_/Y _21379_/A vssd1 vssd1 vccd1 vccd1 _22146_/A sky130_fd_sc_hd__a21oi_1
XFILLER_134_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_335_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_307_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22062_ _22031_/A _22031_/B _22030_/A vssd1 vssd1 vccd1 vccd1 _22085_/A sky130_fd_sc_hd__a21o_2
XTAP_6619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21013_ _21013_/A _21043_/B vssd1 vssd1 vccd1 vccd1 _21013_/Y sky130_fd_sc_hd__nand2_1
Xoutput286 _14086_/X vssd1 vssd1 vccd1 vccd1 addr0[1] sky130_fd_sc_hd__buf_2
XFILLER_142_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput297 _13992_/X vssd1 vssd1 vccd1 vccd1 addr1[3] sky130_fd_sc_hd__buf_2
XTAP_5918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_4 _22139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_287_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22964_ _23846_/CLK _22964_/D vssd1 vssd1 vccd1 vccd1 _22964_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21915_ _21892_/A _21892_/B _21889_/A vssd1 vssd1 vccd1 vccd1 _21919_/A sky130_fd_sc_hd__o21ai_1
XFILLER_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22895_ _23424_/CLK _22895_/D vssd1 vssd1 vccd1 vccd1 _22895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21846_ _21846_/A _22044_/A vssd1 vssd1 vccd1 vccd1 _21846_/Y sky130_fd_sc_hd__nor2_1
XPHY_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21777_ _21775_/Y _21772_/Y _21771_/X _21721_/X vssd1 vssd1 vccd1 vccd1 _21778_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_358_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23516_ _23546_/CLK _23516_/D vssd1 vssd1 vccd1 vccd1 _23516_/Q sky130_fd_sc_hd__dfxtp_1
X_11530_ _23330_/Q _23298_/Q _23266_/Q _23554_/Q _11517_/X _11519_/X vssd1 vssd1 vccd1
+ vccd1 _11530_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20728_ _23741_/Q _20697_/X _20727_/X _20706_/X vssd1 vssd1 vccd1 vccd1 _23741_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_345_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23447_ _23544_/CLK _23447_/D vssd1 vssd1 vccd1 vccd1 _23447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11461_ _11461_/A vssd1 vssd1 vccd1 vccd1 _11461_/X sky130_fd_sc_hd__buf_2
XFILLER_109_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20659_ _23730_/Q _20628_/X _20658_/X _20637_/X vssd1 vssd1 vccd1 vccd1 _23730_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_356_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13200_ _12816_/X _13197_/X _13199_/X _11246_/A vssd1 vssd1 vccd1 vccd1 _13200_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14180_ _21925_/A _14180_/B _16118_/A _14180_/D vssd1 vssd1 vccd1 vccd1 _20533_/A
+ sky130_fd_sc_hd__or4_4
X_11392_ _11270_/Y _20400_/A _15565_/A vssd1 vssd1 vccd1 vccd1 _14356_/B sky130_fd_sc_hd__mux2_4
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_353_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23378_ _23535_/CLK _23378_/D vssd1 vssd1 vccd1 vccd1 _23378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_341_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_326_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13131_ _13131_/A _13131_/B vssd1 vssd1 vccd1 vccd1 _13131_/Y sky130_fd_sc_hd__nor2_1
XFILLER_136_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22329_ _23525_/CLK _22329_/D vssd1 vssd1 vccd1 vccd1 _22329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_314_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_297_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13062_ _13131_/A _13062_/B vssd1 vssd1 vccd1 vccd1 _13062_/Y sky130_fd_sc_hd__nor2_1
XFILLER_279_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12013_ _12029_/A vssd1 vssd1 vccd1 vccd1 _12013_/X sky130_fd_sc_hd__buf_4
XFILLER_155_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17870_ _22806_/Q _17639_/X _17870_/S vssd1 vssd1 vccd1 vccd1 _17871_/A sky130_fd_sc_hd__mux2_1
XFILLER_340_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_321_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_305_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_305_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16821_ _16821_/A vssd1 vssd1 vccd1 vccd1 _22522_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19540_ _19540_/A vssd1 vssd1 vccd1 vccd1 _19549_/S sky130_fd_sc_hd__buf_4
X_16752_ _22503_/Q _16747_/X _16748_/X input17/X vssd1 vssd1 vccd1 vccd1 _16753_/B
+ sky130_fd_sc_hd__o22a_1
X_13964_ _13964_/A _13965_/B vssd1 vssd1 vccd1 vccd1 _13964_/Y sky130_fd_sc_hd__nor2_1
XFILLER_219_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15703_ _21868_/B _21868_/C _15891_/A vssd1 vssd1 vccd1 vccd1 _15703_/Y sky130_fd_sc_hd__o21ai_4
X_12915_ _13493_/A _13493_/B vssd1 vssd1 vccd1 vccd1 _12916_/B sky130_fd_sc_hd__nor2_2
XFILLER_111_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19471_ _23391_/Q _18856_/X _19477_/S vssd1 vssd1 vccd1 vccd1 _19472_/A sky130_fd_sc_hd__mux2_1
X_16683_ _22486_/Q _16679_/Y _16810_/B _16808_/B vssd1 vssd1 vccd1 vccd1 _22486_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13895_ _13895_/A vssd1 vssd1 vccd1 vccd1 _21351_/A sky130_fd_sc_hd__buf_4
XFILLER_235_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18422_ _22968_/Q _18420_/B _18421_/Y vssd1 vssd1 vccd1 vccd1 _22968_/D sky130_fd_sc_hd__o21a_1
XFILLER_222_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15634_ _15633_/X _15244_/Y _15674_/A vssd1 vssd1 vccd1 vccd1 _15634_/X sky130_fd_sc_hd__a21bo_2
X_12846_ _12904_/A _12846_/B vssd1 vssd1 vccd1 vccd1 _12846_/X sky130_fd_sc_hd__or2_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _22944_/Q _18351_/B _18352_/Y vssd1 vssd1 vccd1 vccd1 _22944_/D sky130_fd_sc_hd__o21a_1
XFILLER_221_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _15565_/A vssd1 vssd1 vccd1 vccd1 _15818_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12777_ _12777_/A vssd1 vssd1 vccd1 vccd1 _12777_/X sky130_fd_sc_hd__buf_4
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17304_ _22582_/Q _17255_/X _17028_/A _17303_/X vssd1 vssd1 vccd1 vccd1 _22582_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14516_/A vssd1 vssd1 vccd1 vccd1 _14936_/A sky130_fd_sc_hd__buf_8
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18284_ _18286_/A _18286_/C _18283_/Y vssd1 vssd1 vccd1 vccd1 _22921_/D sky130_fd_sc_hd__o21a_1
XFILLER_202_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11728_ _23910_/Q _13803_/A _12135_/A vssd1 vssd1 vccd1 vccd1 _13500_/B sky130_fd_sc_hd__mux2_2
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15496_ _15479_/B _15718_/B _15636_/A vssd1 vssd1 vccd1 vccd1 _15496_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_308_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17235_ _22029_/A _17234_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17235_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14447_ _14447_/A _14506_/B _20770_/A vssd1 vssd1 vccd1 vccd1 _14731_/A sky130_fd_sc_hd__or3_4
XFILLER_317_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11659_ _11659_/A vssd1 vssd1 vccd1 vccd1 _12334_/A sky130_fd_sc_hd__buf_2
XFILLER_266_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17166_ _22569_/Q _17141_/X _17131_/X _17165_/X vssd1 vssd1 vccd1 vccd1 _22569_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_190_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14378_ _15130_/S _14381_/B vssd1 vssd1 vccd1 vccd1 _14767_/A sky130_fd_sc_hd__or2_1
XFILLER_7_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16117_ _15564_/A _13549_/B _15574_/X _16116_/X vssd1 vssd1 vccd1 vccd1 _16117_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_317_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13329_ _13329_/A _13632_/A vssd1 vssd1 vccd1 vccd1 _13395_/B sky130_fd_sc_hd__xnor2_4
X_17097_ _17250_/A vssd1 vssd1 vccd1 vccd1 _17137_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_304_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16048_ _18859_/A vssd1 vssd1 vccd1 vccd1 _19252_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_320_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19807_ _23540_/Q _19213_/A _19815_/S vssd1 vssd1 vccd1 vccd1 _19808_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17999_ _22841_/Q _17990_/X _17986_/X _17998_/X _17983_/X vssd1 vssd1 vccd1 vccd1
+ _17999_/X sky130_fd_sc_hd__a221o_1
XFILLER_215_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19738_ _19738_/A vssd1 vssd1 vccd1 vccd1 _23509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19669_ _19223_/X _23479_/Q _19671_/S vssd1 vssd1 vccd1 vccd1 _19670_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21700_ _22093_/A vssd1 vssd1 vccd1 vccd1 _21714_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22680_ _23047_/CLK _22680_/D vssd1 vssd1 vccd1 vccd1 _22680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21631_ _21585_/A _21587_/B _21630_/X vssd1 vssd1 vccd1 vccd1 _21632_/B sky130_fd_sc_hd__a21oi_2
XFILLER_339_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21562_ _23821_/Q _23755_/Q vssd1 vssd1 vccd1 vccd1 _21564_/A sky130_fd_sc_hd__nor2_1
XFILLER_327_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23301_ _23397_/CLK _23301_/D vssd1 vssd1 vccd1 vccd1 _23301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_339_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20513_ _23716_/Q _20523_/B _20513_/C vssd1 vssd1 vccd1 vccd1 _20515_/C sky130_fd_sc_hd__and3_1
XFILLER_193_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21493_ _23819_/Q _23753_/Q vssd1 vssd1 vccd1 vccd1 _21494_/B sky130_fd_sc_hd__nand2_1
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23232_ _23264_/CLK _23232_/D vssd1 vssd1 vccd1 vccd1 _23232_/Q sky130_fd_sc_hd__dfxtp_1
X_20444_ _21025_/A _20463_/B vssd1 vssd1 vccd1 vccd1 _20444_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_335_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23163_ _23549_/CLK _23163_/D vssd1 vssd1 vccd1 vccd1 _23163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20375_ _17279_/A _20295_/X _20376_/B vssd1 vssd1 vccd1 vccd1 _20375_/X sky130_fd_sc_hd__o21a_1
XTAP_7106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_311_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22114_ _22114_/A _22119_/A vssd1 vssd1 vccd1 vccd1 _22114_/Y sky130_fd_sc_hd__nand2_1
XTAP_7139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23094_ _23510_/CLK _23094_/D vssd1 vssd1 vccd1 vccd1 _23094_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_304_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22045_ _22045_/A vssd1 vssd1 vccd1 vccd1 _22045_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_288_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_291_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_188_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23903_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_275_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_117_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23600_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_228_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22947_ _22947_/CLK _22947_/D vssd1 vssd1 vccd1 vccd1 _22947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12700_ _12700_/A vssd1 vssd1 vccd1 vccd1 _12700_/X sky130_fd_sc_hd__buf_2
X_13680_ _13882_/A vssd1 vssd1 vccd1 vccd1 _13890_/B sky130_fd_sc_hd__clkbuf_2
X_22878_ _23584_/CLK _22878_/D vssd1 vssd1 vccd1 vccd1 _22878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12631_ _22470_/Q _22630_/Q _22309_/Q _23445_/Q _12029_/X _12717_/A vssd1 vssd1 vccd1
+ vccd1 _12631_/X sky130_fd_sc_hd__mux4_1
XPHY_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21829_ _21829_/A _21829_/B vssd1 vssd1 vccd1 vccd1 _21829_/Y sky130_fd_sc_hd__nor2_1
XFILLER_358_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15350_ _16177_/S vssd1 vssd1 vccd1 vccd1 _16070_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_180_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_346_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12562_ _12196_/X _12559_/X _12561_/X _11706_/A vssd1 vssd1 vccd1 vccd1 _12562_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14301_ _12163_/Y _12807_/Y _14329_/S vssd1 vssd1 vccd1 vccd1 _14301_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11513_ _11403_/X _11511_/Y _14179_/A _11486_/B vssd1 vssd1 vccd1 vccd1 _11557_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_12_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15281_ _11884_/Y _15048_/X _15278_/X _21594_/A _15041_/X vssd1 vssd1 vccd1 vccd1
+ _18801_/A sky130_fd_sc_hd__a32o_4
X_12493_ _12519_/A _12493_/B _12493_/C vssd1 vssd1 vccd1 vccd1 _12493_/X sky130_fd_sc_hd__and3_4
X_17020_ _17020_/A _17033_/B vssd1 vssd1 vccd1 vccd1 _17020_/Y sky130_fd_sc_hd__nand2_1
X_14232_ _14232_/A vssd1 vssd1 vccd1 vccd1 _14232_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_345_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11444_ _14393_/A _11438_/X _11443_/X vssd1 vssd1 vccd1 vccd1 _11444_/X sky130_fd_sc_hd__a21o_1
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_314_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14163_ _22908_/Q _14160_/X _16929_/A _22601_/Q vssd1 vssd1 vccd1 vccd1 _14553_/A
+ sky130_fd_sc_hd__a22oi_2
X_11375_ _11375_/A vssd1 vssd1 vccd1 vccd1 _11826_/A sky130_fd_sc_hd__buf_4
XFILLER_180_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13114_ _13114_/A vssd1 vssd1 vccd1 vccd1 _13114_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14094_ _22594_/Q _14081_/A _14093_/Y _14083_/X vssd1 vssd1 vccd1 vccd1 _14094_/X
+ sky130_fd_sc_hd__a22o_4
X_18971_ _16847_/X _23183_/Q _18979_/S vssd1 vssd1 vccd1 vccd1 _18972_/A sky130_fd_sc_hd__mux2_1
XFILLER_332_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_316_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17922_ _17956_/A vssd1 vssd1 vccd1 vccd1 _17922_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_279_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13045_ _23328_/Q _23296_/Q _23264_/Q _23552_/Q _11432_/A _13037_/X vssd1 vssd1 vccd1
+ vccd1 _13046_/B sky130_fd_sc_hd__mux4_1
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17853_ _22798_/Q _17614_/X _17859_/S vssd1 vssd1 vccd1 vccd1 _17854_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16804_ _16804_/A _16804_/B vssd1 vssd1 vccd1 vccd1 _16805_/A sky130_fd_sc_hd__or2_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17784_ _17784_/A vssd1 vssd1 vccd1 vccd1 _22767_/D sky130_fd_sc_hd__clkbuf_1
X_14996_ _23818_/Q _14907_/X _14992_/X _14995_/X _14923_/X vssd1 vssd1 vccd1 vccd1
+ _14996_/X sky130_fd_sc_hd__a221o_4
XFILLER_82_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19523_ _19220_/X _23414_/Q _19527_/S vssd1 vssd1 vccd1 vccd1 _19524_/A sky130_fd_sc_hd__mux2_1
XFILLER_281_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16735_ _16741_/A _16735_/B vssd1 vssd1 vccd1 vccd1 _16736_/A sky130_fd_sc_hd__or2_1
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13947_ _16679_/B _14097_/A vssd1 vssd1 vccd1 vccd1 _13947_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16666_ _16666_/A vssd1 vssd1 vccd1 vccd1 _22479_/D sky130_fd_sc_hd__clkbuf_1
X_19454_ _19454_/A vssd1 vssd1 vccd1 vccd1 _23383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13878_ _13892_/A _14069_/C vssd1 vssd1 vccd1 vccd1 _13878_/Y sky130_fd_sc_hd__nor2_1
XFILLER_262_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18405_ _15644_/A _18409_/C _18380_/X vssd1 vssd1 vccd1 vccd1 _18405_/Y sky130_fd_sc_hd__a21oi_1
X_15617_ _15672_/A vssd1 vssd1 vccd1 vccd1 _15617_/X sky130_fd_sc_hd__clkbuf_2
X_12829_ _23324_/Q _23292_/Q _23260_/Q _23548_/Q _12825_/X _12672_/A vssd1 vssd1 vccd1
+ vccd1 _12830_/B sky130_fd_sc_hd__mux4_2
XFILLER_201_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19385_ _19396_/A vssd1 vssd1 vccd1 vccd1 _19394_/S sky130_fd_sc_hd__buf_2
X_16597_ _16049_/X _22449_/Q _16601_/S vssd1 vssd1 vccd1 vccd1 _16598_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18336_ _22938_/Q _18334_/B _18335_/Y vssd1 vssd1 vccd1 vccd1 _22938_/D sky130_fd_sc_hd__o21a_1
XFILLER_231_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15548_ _22961_/Q _16177_/S vssd1 vssd1 vccd1 vccd1 _15548_/X sky130_fd_sc_hd__or2_1
XFILLER_348_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18267_ _18279_/D vssd1 vssd1 vccd1 vccd1 _18275_/C sky130_fd_sc_hd__clkbuf_2
X_15479_ _15479_/A _15479_/B vssd1 vssd1 vccd1 vccd1 _15479_/Y sky130_fd_sc_hd__nand2_2
XFILLER_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17218_ _22574_/Q _17199_/X _17190_/X _17217_/X vssd1 vssd1 vccd1 vccd1 _22574_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_190_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18198_ _18198_/A _18198_/B _18164_/B vssd1 vssd1 vccd1 vccd1 _18203_/B sky130_fd_sc_hd__or3b_4
XFILLER_352_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17149_ _17149_/A _17172_/B vssd1 vssd1 vccd1 vccd1 _17149_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20160_ _20160_/A _21084_/B vssd1 vssd1 vccd1 vccd1 _21097_/B sky130_fd_sc_hd__or2_4
XFILLER_157_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20091_ _20098_/C _20098_/D _18012_/X vssd1 vssd1 vccd1 vccd1 _20091_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_301_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23850_ _23851_/CLK _23850_/D vssd1 vssd1 vccd1 vccd1 _23850_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22801_ _22801_/CLK _22801_/D vssd1 vssd1 vccd1 vccd1 _22801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23781_ _23946_/CLK _23781_/D vssd1 vssd1 vccd1 vccd1 _23781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20993_ _21064_/B vssd1 vssd1 vccd1 vccd1 _20993_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22732_ _23450_/CLK _22732_/D vssd1 vssd1 vccd1 vccd1 _22732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_2_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_309_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22663_ _22695_/CLK _22663_/D vssd1 vssd1 vccd1 vccd1 _22663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21614_ _21604_/A _21614_/B vssd1 vssd1 vccd1 vccd1 _21624_/C sky130_fd_sc_hd__and2b_1
XFILLER_240_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22594_ _22977_/CLK _22594_/D vssd1 vssd1 vccd1 vccd1 _22594_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_205_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21545_ _21451_/A _21544_/X _21546_/B _21542_/C _21542_/A vssd1 vssd1 vccd1 vccd1
+ _21545_/X sky130_fd_sc_hd__o2111a_1
XFILLER_224_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21476_ _21981_/A _21476_/B vssd1 vssd1 vccd1 vccd1 _21476_/Y sky130_fd_sc_hd__nand2_1
XFILLER_308_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23215_ _23535_/CLK _23215_/D vssd1 vssd1 vccd1 vccd1 _23215_/Q sky130_fd_sc_hd__dfxtp_1
X_20427_ _20595_/A _20408_/X _20426_/X _20420_/X vssd1 vssd1 vccd1 vccd1 _23690_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_355_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_335_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23146_ _23370_/CLK _23146_/D vssd1 vssd1 vccd1 vccd1 _23146_/Q sky130_fd_sc_hd__dfxtp_1
X_11160_ _12538_/A vssd1 vssd1 vccd1 vccd1 _12425_/A sky130_fd_sc_hd__buf_6
X_20358_ _20808_/A vssd1 vssd1 vccd1 vccd1 _20963_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_353_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_351_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_310_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11091_ _12544_/B vssd1 vssd1 vccd1 vccd1 _13472_/A sky130_fd_sc_hd__buf_2
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23077_ _23493_/CLK _23077_/D vssd1 vssd1 vccd1 vccd1 _23077_/Q sky130_fd_sc_hd__dfxtp_1
X_20289_ _20376_/A _20289_/B vssd1 vssd1 vccd1 vccd1 _20289_/Y sky130_fd_sc_hd__nor2_1
XTAP_6246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22028_ _22029_/A _22032_/A vssd1 vssd1 vccd1 vccd1 _22030_/A sky130_fd_sc_hd__and2_1
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14850_ _14634_/X _14637_/X _14850_/S vssd1 vssd1 vccd1 vccd1 _14850_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _13855_/A _13801_/B vssd1 vssd1 vccd1 vccd1 _13802_/A sky130_fd_sc_hd__and2_1
XFILLER_264_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14781_ _14323_/A _14328_/X _14841_/S vssd1 vssd1 vccd1 vccd1 _14781_/X sky130_fd_sc_hd__mux2_1
X_11993_ _12909_/A _11993_/B vssd1 vssd1 vccd1 vccd1 _11993_/X sky130_fd_sc_hd__or2_1
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_290_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16520_ _16049_/X _22416_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _16521_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13732_ _15176_/A _21191_/A vssd1 vssd1 vccd1 vccd1 _13777_/B sky130_fd_sc_hd__nor2_2
XFILLER_217_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16451_ _16124_/X _22386_/Q _16451_/S vssd1 vssd1 vccd1 vccd1 _16452_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13663_ _22607_/Q _22608_/Q _22609_/Q _22610_/Q vssd1 vssd1 vccd1 vccd1 _13670_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_16_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15402_ _23825_/Q _14906_/A _15398_/X _15401_/X _14610_/A vssd1 vssd1 vccd1 vccd1
+ _15402_/X sky130_fd_sc_hd__a221o_2
XFILLER_232_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19170_ _19169_/X _23270_/Q _19179_/S vssd1 vssd1 vccd1 vccd1 _19171_/A sky130_fd_sc_hd__mux2_1
X_12614_ _12233_/X _15122_/A _12613_/X _12161_/X vssd1 vssd1 vccd1 vccd1 _13349_/B
+ sky130_fd_sc_hd__a211o_4
X_16382_ _16382_/A vssd1 vssd1 vccd1 vccd1 _22356_/D sky130_fd_sc_hd__clkbuf_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13594_ _13594_/A vssd1 vssd1 vccd1 vccd1 _14198_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_346_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18121_ _18245_/A vssd1 vssd1 vccd1 vccd1 _18121_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_85_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23449_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_197_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15333_ _13738_/A _15331_/Y _15332_/Y _13834_/A vssd1 vssd1 vccd1 vccd1 _15333_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_61_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12545_ _11404_/A _13695_/B _12544_/X _12344_/X vssd1 vssd1 vccd1 vccd1 _13361_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23535_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18052_ _18052_/A vssd1 vssd1 vccd1 vccd1 _18052_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15264_ _23790_/Q _14605_/X _14606_/X vssd1 vssd1 vccd1 vccd1 _15264_/X sky130_fd_sc_hd__a21o_1
X_12476_ _12476_/A vssd1 vssd1 vccd1 vccd1 _12476_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_333_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17003_ _20517_/B vssd1 vssd1 vccd1 vccd1 _20524_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14215_ _14215_/A vssd1 vssd1 vccd1 vccd1 _14215_/X sky130_fd_sc_hd__clkbuf_2
X_11427_ _11420_/Y _11422_/Y _11424_/Y _11426_/Y _11247_/X vssd1 vssd1 vccd1 vccd1
+ _11451_/B sky130_fd_sc_hd__o221ai_1
X_15195_ _15020_/S _15131_/Y _14630_/X vssd1 vssd1 vccd1 vccd1 _15195_/X sky130_fd_sc_hd__a21o_1
XFILLER_126_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_298_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14146_ _14211_/B _16945_/A vssd1 vssd1 vccd1 vccd1 _14159_/A sky130_fd_sc_hd__nand2_1
XFILLER_113_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ _11659_/A _12329_/A _11821_/A _11457_/D vssd1 vssd1 vccd1 vccd1 _12519_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_287_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_302_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_301_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14077_ _14241_/A _15112_/A _13890_/Y vssd1 vssd1 vccd1 vccd1 _15056_/A sky130_fd_sc_hd__a21oi_4
X_18954_ _18954_/A vssd1 vssd1 vccd1 vccd1 _23175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11289_ _23896_/Q vssd1 vssd1 vccd1 vccd1 _12511_/A sky130_fd_sc_hd__inv_2
XFILLER_98_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17905_ _22814_/Q _17891_/X _17904_/X _17657_/X vssd1 vssd1 vccd1 vccd1 _22814_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_267_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13028_ _13028_/A vssd1 vssd1 vccd1 vccd1 _13029_/B sky130_fd_sc_hd__inv_2
XFILLER_112_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18885_ _23145_/Q _18785_/X _18885_/S vssd1 vssd1 vccd1 vccd1 _18886_/A sky130_fd_sc_hd__mux2_1
XTAP_6780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17836_ _17836_/A vssd1 vssd1 vccd1 vccd1 _22790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17767_ _17789_/A vssd1 vssd1 vccd1 vccd1 _17776_/S sky130_fd_sc_hd__buf_4
XFILLER_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14979_ _14819_/X _14971_/X _14978_/Y _14698_/X vssd1 vssd1 vccd1 vccd1 _14979_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_281_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19506_ _19506_/A vssd1 vssd1 vccd1 vccd1 _23406_/D sky130_fd_sc_hd__clkbuf_1
X_16718_ _16718_/A vssd1 vssd1 vccd1 vccd1 _22493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17698_ _22729_/Q _17598_/X _17704_/S vssd1 vssd1 vccd1 vccd1 _17699_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_420 _14062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_431 _23880_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19437_ _19437_/A vssd1 vssd1 vccd1 vccd1 _23375_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_442 _23917_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16649_ _22472_/Q _16265_/X _16651_/S vssd1 vssd1 vccd1 vccd1 _16650_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_453 _22602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_288_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_464 _21281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_475 _21716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_486 _13970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19368_ _23345_/Q _18811_/X _19372_/S vssd1 vssd1 vccd1 vccd1 _19369_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_497 _14574_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18319_ _15724_/X _18323_/C _18292_/X vssd1 vssd1 vccd1 vccd1 _18319_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19299_ _19299_/A vssd1 vssd1 vccd1 vccd1 _23314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_337_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_309_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21330_ _21307_/X _21314_/Y _21325_/X _21327_/X _21329_/X vssd1 vssd1 vccd1 vccd1
+ _21330_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_337_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_318_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21261_ _22254_/A _21261_/B vssd1 vssd1 vccd1 vccd1 _21262_/A sky130_fd_sc_hd__and2_1
XFILLER_317_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23000_ _23592_/CLK _23000_/D vssd1 vssd1 vccd1 vccd1 _23000_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_351_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_5_0_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_20212_ _20146_/X _20595_/A _20211_/X _20203_/X vssd1 vssd1 vccd1 vccd1 _23658_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_150_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21192_ _21192_/A vssd1 vssd1 vccd1 vccd1 _21193_/C sky130_fd_sc_hd__inv_2
XFILLER_144_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_289_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20143_ _20143_/A vssd1 vssd1 vccd1 vccd1 _20890_/B sky130_fd_sc_hd__buf_2
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20074_ _23633_/Q _20072_/B _18268_/A vssd1 vssd1 vccd1 vccd1 _20074_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_106_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23902_ _23902_/CLK _23902_/D vssd1 vssd1 vccd1 vccd1 _23902_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23833_ _23871_/CLK _23833_/D vssd1 vssd1 vccd1 vccd1 _23833_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23764_ _23804_/CLK _23764_/D vssd1 vssd1 vccd1 vccd1 _23764_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20976_ _23808_/Q _20969_/X _20975_/X _20964_/X vssd1 vssd1 vccd1 vccd1 _23808_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22715_ _23054_/CLK _22715_/D vssd1 vssd1 vccd1 vccd1 _22715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_281_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23695_ _23696_/CLK _23695_/D vssd1 vssd1 vccd1 vccd1 _23695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22646_ _23896_/CLK _22646_/D vssd1 vssd1 vccd1 vccd1 _22646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_327_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22577_ _23643_/CLK _22577_/D vssd1 vssd1 vccd1 vccd1 _22577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12330_ _23466_/Q _23562_/Q _22526_/Q _22330_/Q _11799_/A _12329_/X vssd1 vssd1 vccd1
+ vccd1 _12331_/B sky130_fd_sc_hd__mux4_1
XFILLER_343_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21528_ _21528_/A _21528_/B vssd1 vssd1 vccd1 vccd1 _21528_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_342_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12261_ _23905_/Q _11911_/B _11935_/B vssd1 vssd1 vccd1 vccd1 _12261_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_181_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21459_ _23818_/Q _23752_/Q vssd1 vssd1 vccd1 vccd1 _21459_/Y sky130_fd_sc_hd__nand2_1
X_14000_ _14000_/A _14099_/A vssd1 vssd1 vccd1 vccd1 _14000_/Y sky130_fd_sc_hd__nor2_8
X_11212_ _23903_/Q vssd1 vssd1 vccd1 vccd1 _11240_/A sky130_fd_sc_hd__buf_4
XFILLER_330_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12192_ _12535_/S vssd1 vssd1 vccd1 vccd1 _12244_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_351_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_351_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23129_ _23545_/CLK _23129_/D vssd1 vssd1 vccd1 vccd1 _23129_/Q sky130_fd_sc_hd__dfxtp_1
X_11143_ _13084_/A vssd1 vssd1 vccd1 vccd1 _13199_/A sky130_fd_sc_hd__clkbuf_2
XTAP_6010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_296_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_132_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _22971_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15951_ _15950_/X _14509_/A _14513_/A _22971_/Q vssd1 vssd1 vccd1 vccd1 _15951_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_110_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11074_ _23884_/Q vssd1 vssd1 vccd1 vccd1 _14172_/B sky130_fd_sc_hd__clkbuf_2
XTAP_6076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput120 dout1[21] vssd1 vssd1 vccd1 vccd1 input120/X sky130_fd_sc_hd__clkbuf_1
XTAP_5331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput131 dout1[31] vssd1 vssd1 vccd1 vccd1 input131/X sky130_fd_sc_hd__clkbuf_1
XTAP_6087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput142 dout1[41] vssd1 vssd1 vccd1 vccd1 input142/X sky130_fd_sc_hd__buf_2
X_14902_ _14902_/A vssd1 vssd1 vccd1 vccd1 _14902_/X sky130_fd_sc_hd__clkbuf_2
XTAP_6098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput153 dout1[51] vssd1 vssd1 vccd1 vccd1 input153/X sky130_fd_sc_hd__buf_2
X_18670_ _18670_/A vssd1 vssd1 vccd1 vccd1 _23064_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15882_ _23836_/Q _14907_/X _15878_/X _15881_/X _15222_/X vssd1 vssd1 vccd1 vccd1
+ _15882_/X sky130_fd_sc_hd__a221o_1
Xinput164 dout1[61] vssd1 vssd1 vccd1 vccd1 input164/X sky130_fd_sc_hd__buf_2
XFILLER_264_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput175 irq[13] vssd1 vssd1 vccd1 vccd1 _20510_/C sky130_fd_sc_hd__clkbuf_4
XTAP_5397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput186 irq[9] vssd1 vssd1 vccd1 vccd1 _20507_/C sky130_fd_sc_hd__buf_2
XFILLER_313_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17621_ _22701_/Q _17620_/X _17624_/S vssd1 vssd1 vccd1 vccd1 _17622_/A sky130_fd_sc_hd__mux2_1
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput197 localMemory_wb_adr_i[16] vssd1 vssd1 vccd1 vccd1 input197/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_252_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14833_ _14833_/A vssd1 vssd1 vccd1 vccd1 _15865_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_264_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ _17552_/A vssd1 vssd1 vccd1 vccd1 _22679_/D sky130_fd_sc_hd__clkbuf_1
X_14764_ _15491_/S vssd1 vssd1 vccd1 vccd1 _15341_/S sky130_fd_sc_hd__clkbuf_2
X_11976_ _23476_/Q _23572_/Q _22536_/Q _22340_/Q _12675_/A _12746_/A vssd1 vssd1 vccd1
+ vccd1 _11976_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16503_ _16503_/A vssd1 vssd1 vccd1 vccd1 _22408_/D sky130_fd_sc_hd__clkbuf_1
X_13715_ _13715_/A _13728_/B _14015_/C vssd1 vssd1 vccd1 vccd1 _13716_/A sky130_fd_sc_hd__and3_4
XFILLER_205_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17483_ _22650_/Q _16220_/X _17483_/S vssd1 vssd1 vccd1 vccd1 _17484_/A sky130_fd_sc_hd__mux2_1
X_14695_ _15367_/A _14695_/B vssd1 vssd1 vccd1 vccd1 _14695_/Y sky130_fd_sc_hd__nor2_1
XFILLER_232_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19222_ _19222_/A vssd1 vssd1 vccd1 vccd1 _23286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16434_ _15823_/X _22378_/Q _16440_/S vssd1 vssd1 vccd1 vccd1 _16435_/A sky130_fd_sc_hd__mux2_1
X_13646_ _13646_/A _13646_/B vssd1 vssd1 vccd1 vccd1 _15335_/A sky130_fd_sc_hd__xnor2_4
XFILLER_176_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_347_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19153_ _23264_/Q _18859_/X _19157_/S vssd1 vssd1 vccd1 vccd1 _19154_/A sky130_fd_sc_hd__mux2_1
X_16365_ _16365_/A vssd1 vssd1 vccd1 vccd1 _22348_/D sky130_fd_sc_hd__clkbuf_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ _23935_/Q vssd1 vssd1 vccd1 vccd1 _17246_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_358_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_338_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18104_ _22872_/Q _18097_/X _18098_/X _23005_/Q _18099_/X vssd1 vssd1 vccd1 vccd1
+ _18104_/X sky130_fd_sc_hd__a221o_1
X_15316_ _21636_/A _15316_/B vssd1 vssd1 vccd1 vccd1 _15317_/B sky130_fd_sc_hd__nor2_1
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12528_ _23301_/Q _23269_/Q _23237_/Q _23525_/Q _12457_/S _12538_/A vssd1 vssd1 vccd1
+ vccd1 _12529_/B sky130_fd_sc_hd__mux4_2
X_16296_ _16296_/A vssd1 vssd1 vccd1 vccd1 _22320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_258_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19084_ _16908_/X _23234_/Q _19084_/S vssd1 vssd1 vccd1 vccd1 _19085_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_338_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18035_ _18051_/A vssd1 vssd1 vccd1 vccd1 _18035_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_184_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15247_ _13526_/A _14254_/X _14761_/X _13524_/Y _14682_/A vssd1 vssd1 vccd1 vccd1
+ _15247_/X sky130_fd_sc_hd__a221o_1
X_12459_ _22778_/Q _22746_/Q _22647_/Q _22714_/Q _12537_/S _12449_/X vssd1 vssd1 vccd1
+ vccd1 _12459_/X sky130_fd_sc_hd__mux4_2
XFILLER_274_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_315_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15178_ _15187_/B vssd1 vssd1 vccd1 vccd1 _15901_/B sky130_fd_sc_hd__clkinv_2
XFILLER_302_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_287_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_315_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14129_ _22712_/Q vssd1 vssd1 vccd1 vccd1 _14415_/S sky130_fd_sc_hd__inv_2
XFILLER_98_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19986_ _20008_/A _19986_/B _20003_/C vssd1 vssd1 vccd1 vccd1 _23608_/D sky130_fd_sc_hd__nor3_1
XFILLER_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_259_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18937_ _18937_/A vssd1 vssd1 vccd1 vccd1 _23168_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_274_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18868_ _18868_/A vssd1 vssd1 vccd1 vccd1 _18868_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_283_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17819_ _17819_/A vssd1 vssd1 vccd1 vccd1 _22782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_282_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18799_ _23117_/Q _18798_/X _18802_/S vssd1 vssd1 vccd1 vccd1 _18800_/A sky130_fd_sc_hd__mux2_1
XFILLER_255_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20830_ _20665_/B _20828_/X _20829_/X _23763_/Q vssd1 vssd1 vccd1 vccd1 _20831_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_345_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20761_ _22217_/A _20632_/A _20760_/X vssd1 vssd1 vccd1 vccd1 _20762_/C sky130_fd_sc_hd__o21a_1
XINSDIODE2_250 _21737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22500_ _23704_/CLK _22500_/D vssd1 vssd1 vccd1 vccd1 _22500_/Q sky130_fd_sc_hd__dfxtp_4
XINSDIODE2_261 _15651_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_272 _18827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_357_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23480_ _23480_/CLK _23480_/D vssd1 vssd1 vccd1 vccd1 _23480_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_167_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_283 _22067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_294 _15990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20692_ _20724_/A vssd1 vssd1 vccd1 vccd1 _20692_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_189_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22431_ _23502_/CLK _22431_/D vssd1 vssd1 vccd1 vccd1 _22431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22362_ _23564_/CLK _22362_/D vssd1 vssd1 vccd1 vccd1 _22362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_325_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_309_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_337_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21313_ _21346_/A _21313_/B vssd1 vssd1 vccd1 vccd1 _21313_/X sky130_fd_sc_hd__and2b_1
XFILLER_325_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22293_ _23527_/CLK _22293_/D vssd1 vssd1 vccd1 vccd1 _22293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_324_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_312_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21244_ _21244_/A _21274_/B vssd1 vssd1 vccd1 vccd1 _21244_/Y sky130_fd_sc_hd__nand2_1
XFILLER_321_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_352_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21175_ _21681_/A vssd1 vssd1 vccd1 vccd1 _21175_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_321_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20126_ _23648_/Q _23647_/Q _20126_/C _20126_/D vssd1 vssd1 vccd1 vccd1 _20127_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_89_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20057_ _20086_/A _20057_/B _20076_/C vssd1 vssd1 vccd1 vccd1 _23628_/D sky130_fd_sc_hd__nor3_1
XFILLER_274_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23816_ _23818_/CLK _23816_/D vssd1 vssd1 vccd1 vccd1 _23816_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_73_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _11939_/A _11939_/B vssd1 vssd1 vccd1 vccd1 _13392_/A sky130_fd_sc_hd__and2b_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _12634_/A _11761_/B _11761_/C vssd1 vssd1 vccd1 vccd1 _21648_/A sky130_fd_sc_hd__nor3_4
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23747_ _23866_/CLK _23747_/D vssd1 vssd1 vccd1 vccd1 _23747_/Q sky130_fd_sc_hd__dfxtp_1
X_20959_ _23933_/Q vssd1 vssd1 vccd1 vccd1 _21999_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13500_/A _13500_/B _13521_/B vssd1 vssd1 vccd1 vccd1 _13501_/A sky130_fd_sc_hd__and3_1
XFILLER_214_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14910_/A vssd1 vssd1 vccd1 vccd1 _15595_/A sky130_fd_sc_hd__buf_4
XFILLER_158_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11692_ _13532_/A vssd1 vssd1 vccd1 vccd1 _13608_/A sky130_fd_sc_hd__clkinv_4
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23678_ _23714_/CLK _23678_/D vssd1 vssd1 vccd1 vccd1 _23678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_329_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13431_ _21336_/A vssd1 vssd1 vccd1 vccd1 _13432_/B sky130_fd_sc_hd__buf_2
X_22629_ _22632_/CLK _22629_/D vssd1 vssd1 vccd1 vccd1 _22629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_329_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16150_ _23940_/Q vssd1 vssd1 vccd1 vccd1 _22219_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13362_ _14290_/A _13362_/B vssd1 vssd1 vccd1 vccd1 _13363_/B sky130_fd_sc_hd__nor2_2
XFILLER_155_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15101_ _22984_/Q _14138_/A _15164_/A input243/X vssd1 vssd1 vccd1 vccd1 _21500_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_139_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12313_ _11911_/B _13764_/A _12312_/Y vssd1 vssd1 vccd1 vccd1 _13514_/A sky130_fd_sc_hd__a21oi_4
XFILLER_182_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16081_ _16005_/X _13566_/B _15478_/A vssd1 vssd1 vccd1 vccd1 _16081_/X sky130_fd_sc_hd__a21o_1
X_13293_ _11343_/A _13292_/X _11353_/A vssd1 vssd1 vccd1 vccd1 _13293_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_154_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_344_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_315_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15032_ _14218_/X _15432_/A _15433_/A _13829_/B _15031_/Y vssd1 vssd1 vccd1 vccd1
+ _15032_/Y sky130_fd_sc_hd__o221ai_1
X_12244_ _12244_/A vssd1 vssd1 vccd1 vccd1 _12245_/S sky130_fd_sc_hd__buf_4
XFILLER_343_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_331_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_308_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_330_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19840_ _19840_/A vssd1 vssd1 vccd1 vccd1 _23555_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12175_ _23212_/Q _23180_/Q _23148_/Q _23116_/Q _11700_/A _11565_/A vssd1 vssd1 vccd1
+ vccd1 _12176_/B sky130_fd_sc_hd__mux4_2
XFILLER_296_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11126_ _23902_/Q vssd1 vssd1 vccd1 vccd1 _11127_/A sky130_fd_sc_hd__clkbuf_4
X_19771_ _19771_/A _19771_/B vssd1 vssd1 vccd1 vccd1 _19828_/A sky130_fd_sc_hd__nor2_8
XFILLER_123_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16983_ _21317_/A _17163_/B vssd1 vssd1 vccd1 vccd1 _16983_/X sky130_fd_sc_hd__or2_1
XFILLER_150_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_311_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18722_ _16847_/X _23087_/Q _18730_/S vssd1 vssd1 vccd1 vccd1 _18723_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15934_ _15928_/X _15930_/Y _22067_/A _14210_/X vssd1 vssd1 vccd1 vccd1 _18849_/A
+ sky130_fd_sc_hd__o2bb2a_4
XTAP_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18653_ _18653_/A vssd1 vssd1 vccd1 vccd1 _23056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865_ _15865_/A _15865_/B vssd1 vssd1 vccd1 vccd1 _15865_/Y sky130_fd_sc_hd__nand2_2
XFILLER_49_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17604_ _18830_/A vssd1 vssd1 vccd1 vccd1 _17604_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_292_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14816_ _21382_/A _21482_/A vssd1 vssd1 vccd1 vccd1 _20493_/B sky130_fd_sc_hd__nor2_2
XFILLER_184_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18584_ _16857_/X _23026_/Q _18586_/S vssd1 vssd1 vccd1 vccd1 _18585_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_291_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ _13323_/A _13023_/X _13389_/X _15580_/B vssd1 vssd1 vccd1 vccd1 _15797_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_45_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_340_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17535_ _17535_/A vssd1 vssd1 vccd1 vccd1 _22673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11959_ _23220_/Q _23188_/Q _23156_/Q _23124_/Q _12680_/A _12041_/A vssd1 vssd1 vccd1
+ vccd1 _11960_/B sky130_fd_sc_hd__mux4_2
XFILLER_269_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14747_ _23845_/Q _14737_/X _14746_/X vssd1 vssd1 vccd1 vccd1 _14747_/X sky130_fd_sc_hd__o21a_2
XFILLER_33_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_339_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17466_ _17466_/A vssd1 vssd1 vccd1 vccd1 _22643_/D sky130_fd_sc_hd__clkbuf_1
X_14678_ _14815_/B vssd1 vssd1 vccd1 vccd1 _14836_/A sky130_fd_sc_hd__buf_2
XFILLER_220_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19205_ _19204_/X _23281_/Q _19211_/S vssd1 vssd1 vccd1 vccd1 _19206_/A sky130_fd_sc_hd__mux2_1
X_16417_ _16417_/A vssd1 vssd1 vccd1 vccd1 _22370_/D sky130_fd_sc_hd__clkbuf_1
X_13629_ _13629_/A _13629_/B vssd1 vssd1 vccd1 vccd1 _13629_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_158_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17397_ _17397_/A vssd1 vssd1 vccd1 vccd1 _22613_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_319_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_335_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19136_ _19136_/A vssd1 vssd1 vccd1 vccd1 _23256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_346_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16348_ _16348_/A vssd1 vssd1 vccd1 vccd1 _22340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19067_ _16883_/X _23226_/Q _19073_/S vssd1 vssd1 vccd1 vccd1 _19068_/A sky130_fd_sc_hd__mux2_1
X_16279_ _22315_/Q _16278_/X _16285_/S vssd1 vssd1 vccd1 vccd1 _16280_/A sky130_fd_sc_hd__mux2_1
XFILLER_334_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_350_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput402 _14020_/X vssd1 vssd1 vccd1 vccd1 din0[6] sky130_fd_sc_hd__buf_2
X_18018_ _18018_/A _18018_/B _18191_/A vssd1 vssd1 vccd1 vccd1 _18098_/A sky130_fd_sc_hd__and3_4
XFILLER_160_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput413 _22567_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[14] sky130_fd_sc_hd__buf_2
Xoutput424 _22577_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[24] sky130_fd_sc_hd__buf_2
XFILLER_334_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput435 _22558_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput446 _11068_/Y vssd1 vssd1 vccd1 vccd1 probe_isCompressed sky130_fd_sc_hd__buf_2
Xoutput457 _23882_/Q vssd1 vssd1 vccd1 vccd1 probe_opcode[3] sky130_fd_sc_hd__buf_2
XFILLER_330_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput468 _23927_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[16] sky130_fd_sc_hd__buf_2
XFILLER_299_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput479 _23937_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[26] sky130_fd_sc_hd__buf_2
XFILLER_271_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_302_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19969_ _17385_/B _19969_/B _19969_/C _19969_/D vssd1 vssd1 vccd1 vccd1 _19985_/C
+ sky130_fd_sc_hd__and4b_2
XFILLER_102_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22980_ _23424_/CLK _22980_/D vssd1 vssd1 vccd1 vccd1 _22980_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_256_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21931_ _22098_/A _22041_/A vssd1 vssd1 vccd1 vccd1 _21932_/B sky130_fd_sc_hd__nor2_1
XFILLER_41_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21862_ _21859_/Y _21860_/X _21861_/Y _21677_/X vssd1 vssd1 vccd1 vccd1 _21862_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_270_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23601_ _23602_/CLK _23601_/D vssd1 vssd1 vccd1 vccd1 _23601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20813_ _20825_/A _20813_/B vssd1 vssd1 vccd1 vccd1 _20814_/A sky130_fd_sc_hd__and2_1
XFILLER_270_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21793_ _21793_/A _21793_/B vssd1 vssd1 vccd1 vccd1 _21793_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23532_ _23950_/A _23532_/D vssd1 vssd1 vccd1 vccd1 _23532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_251_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20744_ _21177_/A _20744_/B vssd1 vssd1 vccd1 vccd1 _20747_/B sky130_fd_sc_hd__nor2_2
XFILLER_223_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23463_ _23555_/CLK _23463_/D vssd1 vssd1 vccd1 vccd1 _23463_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_357_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20675_ _20675_/A _21301_/C vssd1 vssd1 vccd1 vccd1 _20678_/B sky130_fd_sc_hd__and2_2
XFILLER_195_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22414_ _23583_/CLK _22414_/D vssd1 vssd1 vccd1 vccd1 _22414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_344_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23394_ _23489_/CLK _23394_/D vssd1 vssd1 vccd1 vccd1 _23394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22345_ _23100_/CLK _22345_/D vssd1 vssd1 vccd1 vccd1 _22345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_304_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22276_ _23510_/CLK _22276_/D vssd1 vssd1 vccd1 vccd1 _22276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21227_ _21227_/A _21227_/B vssd1 vssd1 vccd1 vccd1 _21227_/Y sky130_fd_sc_hd__nand2_1
XFILLER_278_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_321_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21158_ _21158_/A vssd1 vssd1 vccd1 vccd1 _21158_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_293_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20109_ _23643_/Q _20107_/C _20108_/Y vssd1 vssd1 vccd1 vccd1 _23643_/D sky130_fd_sc_hd__a21oi_1
XFILLER_144_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13980_ _13980_/A vssd1 vssd1 vccd1 vccd1 _13980_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21089_ _21083_/X _20894_/X _20613_/B _21085_/Y vssd1 vssd1 vccd1 vccd1 _21091_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_247_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12931_ _12968_/A _12931_/B vssd1 vssd1 vccd1 vccd1 _12931_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _12953_/A _12861_/X _12797_/X vssd1 vssd1 vccd1 vccd1 _12862_/X sky130_fd_sc_hd__o21a_1
XFILLER_248_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _23830_/Q _14907_/X _15646_/X _15649_/X _14923_/X vssd1 vssd1 vccd1 vccd1
+ _15650_/X sky130_fd_sc_hd__a221o_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _23471_/Q _23567_/Q _22531_/Q _22335_/Q _12094_/A _11754_/A vssd1 vssd1 vccd1
+ vccd1 _11813_/X sky130_fd_sc_hd__mux4_1
X_14601_ _14601_/A vssd1 vssd1 vccd1 vccd1 _20160_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _13612_/X _15867_/S _15580_/Y _14866_/A vssd1 vssd1 vccd1 vccd1 _15581_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _12793_/A vssd1 vssd1 vccd1 vccd1 _12793_/X sky130_fd_sc_hd__buf_6
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _17242_/A _17314_/X _17319_/X _16997_/X vssd1 vssd1 vccd1 vccd1 _17320_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_214_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14210_/X _17655_/A _14522_/X _14531_/Y vssd1 vssd1 vccd1 vccd1 _18769_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_230_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11744_ _12780_/A _11744_/B vssd1 vssd1 vccd1 vccd1 _11744_/Y sky130_fd_sc_hd__nor2_1
XFILLER_202_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_348_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17251_ _22064_/A _17249_/X _17292_/S vssd1 vssd1 vccd1 vccd1 _17251_/X sky130_fd_sc_hd__mux2_1
X_14463_ _15593_/A vssd1 vssd1 vccd1 vccd1 _15211_/A sky130_fd_sc_hd__buf_2
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11675_ _12028_/A vssd1 vssd1 vccd1 vccd1 _12900_/A sky130_fd_sc_hd__buf_2
X_16202_ _17471_/A _17471_/B _18770_/B vssd1 vssd1 vccd1 vccd1 _19555_/A sky130_fd_sc_hd__nand3_4
XFILLER_146_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13414_ _14288_/A vssd1 vssd1 vccd1 vccd1 _14343_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17182_ _17182_/A vssd1 vssd1 vccd1 vccd1 _17182_/Y sky130_fd_sc_hd__inv_2
XFILLER_316_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14394_ _14394_/A vssd1 vssd1 vccd1 vccd1 _14394_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_319_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_328_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16133_ _14682_/A _16129_/Y _16130_/X _16132_/X vssd1 vssd1 vccd1 vccd1 _16133_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_128_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13345_ _13375_/A _13341_/X _13625_/A _13344_/X vssd1 vssd1 vccd1 vccd1 _13345_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_332_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16064_ _23745_/Q _23875_/Q _16103_/S vssd1 vssd1 vccd1 vccd1 _16064_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13276_ _13276_/A vssd1 vssd1 vccd1 vccd1 _13276_/X sky130_fd_sc_hd__buf_2
XFILLER_6_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_335_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_343_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15015_ _14766_/X _15014_/X _15084_/S vssd1 vssd1 vccd1 vccd1 _15293_/A sky130_fd_sc_hd__mux2_2
XFILLER_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12227_ _12378_/A _12226_/X _11346_/A vssd1 vssd1 vccd1 vccd1 _12227_/X sky130_fd_sc_hd__o21a_1
XFILLER_331_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_312_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19823_ _19823_/A vssd1 vssd1 vccd1 vccd1 _23547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_300_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12158_ _12159_/A _12163_/A vssd1 vssd1 vccd1 vccd1 _12160_/A sky130_fd_sc_hd__and2_1
XFILLER_312_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_12_0_wb_clk_i clkbuf_3_6_1_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _22899_/CLK
+ sky130_fd_sc_hd__clkbuf_4
X_11109_ _23910_/Q vssd1 vssd1 vccd1 vccd1 _14178_/A sky130_fd_sc_hd__buf_6
X_19754_ _19242_/X _23517_/Q _19754_/S vssd1 vssd1 vccd1 vccd1 _19755_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16966_ _16966_/A vssd1 vssd1 vccd1 vccd1 _17262_/A sky130_fd_sc_hd__clkbuf_2
X_12089_ _23924_/Q vssd1 vssd1 vccd1 vccd1 _21719_/A sky130_fd_sc_hd__inv_6
XFILLER_300_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18705_ _18705_/A vssd1 vssd1 vccd1 vccd1 _23079_/D sky130_fd_sc_hd__clkbuf_1
X_15917_ _13399_/B _14942_/A _15916_/Y _13237_/A vssd1 vssd1 vccd1 vccd1 _15920_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19685_ _19245_/X _23486_/Q _19693_/S vssd1 vssd1 vccd1 vccd1 _19686_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16897_ _16895_/X _22546_/Q _16909_/S vssd1 vssd1 vccd1 vccd1 _16898_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18636_ _23049_/Q _17559_/X _18636_/S vssd1 vssd1 vccd1 vccd1 _18637_/A sky130_fd_sc_hd__mux2_1
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _20138_/B _15848_/B vssd1 vssd1 vccd1 vccd1 _15848_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18567_ _16831_/X _23018_/Q _18575_/S vssd1 vssd1 vccd1 vccd1 _18568_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15779_ _13454_/A _15672_/X _15777_/X _15778_/X vssd1 vssd1 vccd1 vccd1 _15779_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_224_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17518_ _17529_/A vssd1 vssd1 vccd1 vccd1 _17527_/S sky130_fd_sc_hd__buf_2
XFILLER_303_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18498_ _22994_/Q _18505_/B vssd1 vssd1 vccd1 vccd1 _18498_/Y sky130_fd_sc_hd__nand2_1
XFILLER_205_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_296_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_296_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17449_ _17449_/A vssd1 vssd1 vccd1 vccd1 _22635_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_354_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20460_ _20680_/A _20447_/X _20457_/X _20459_/X vssd1 vssd1 vccd1 vccd1 _23702_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_335_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_307_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19119_ _19119_/A vssd1 vssd1 vccd1 vccd1 _23248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20391_ _23682_/Q _20391_/B vssd1 vssd1 vccd1 vccd1 _20391_/X sky130_fd_sc_hd__or2_1
XFILLER_335_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_334_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22130_ _23808_/Q _22130_/B vssd1 vssd1 vccd1 vccd1 _22130_/Y sky130_fd_sc_hd__nand2_1
XFILLER_160_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_350_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22061_ _22061_/A _22061_/B vssd1 vssd1 vccd1 vccd1 _22061_/Y sky130_fd_sc_hd__nand2_1
XTAP_6609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21012_ _21072_/B vssd1 vssd1 vccd1 vccd1 _21043_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput287 _14088_/X vssd1 vssd1 vccd1 vccd1 addr0[2] sky130_fd_sc_hd__buf_2
XFILLER_102_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput298 _13996_/Y vssd1 vssd1 vccd1 vccd1 addr1[4] sky130_fd_sc_hd__buf_2
XFILLER_142_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_5 _22166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22963_ _23846_/CLK _22963_/D vssd1 vssd1 vccd1 vccd1 _22963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21914_ _23832_/Q _21913_/X _21973_/S vssd1 vssd1 vccd1 vccd1 _21914_/X sky130_fd_sc_hd__mux2_2
XFILLER_215_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22894_ _23424_/CLK _22894_/D vssd1 vssd1 vccd1 vccd1 _22894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21845_ _21845_/A vssd1 vssd1 vccd1 vccd1 _22044_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_231_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21776_ _21721_/X _21771_/X _21772_/Y _21775_/Y vssd1 vssd1 vccd1 vccd1 _21799_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23515_ _23515_/CLK _23515_/D vssd1 vssd1 vccd1 vccd1 _23515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20727_ _20727_/A _20727_/B _20727_/C vssd1 vssd1 vccd1 vccd1 _20727_/X sky130_fd_sc_hd__or3_1
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23446_ _23446_/CLK _23446_/D vssd1 vssd1 vccd1 vccd1 _23446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_278_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11460_ _13278_/A vssd1 vssd1 vccd1 vccd1 _21848_/A sky130_fd_sc_hd__buf_6
XFILLER_345_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20658_ _20665_/A _20658_/B _20658_/C vssd1 vssd1 vccd1 vccd1 _20658_/X sky130_fd_sc_hd__or3_1
XFILLER_356_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_358_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23377_ _23537_/CLK _23377_/D vssd1 vssd1 vccd1 vccd1 _23377_/Q sky130_fd_sc_hd__dfxtp_1
X_11391_ _11486_/B vssd1 vssd1 vccd1 vccd1 _15565_/A sky130_fd_sc_hd__buf_4
X_20589_ _13440_/C _20773_/A _20574_/X vssd1 vssd1 vccd1 vccd1 _20589_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_99_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_319_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13130_ _22803_/Q _22771_/Q _22672_/Q _22739_/Q _13114_/X _13115_/X vssd1 vssd1 vccd1
+ vccd1 _13131_/B sky130_fd_sc_hd__mux4_2
XFILLER_152_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22328_ _23558_/CLK _22328_/D vssd1 vssd1 vccd1 vccd1 _22328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_341_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13061_ _23488_/Q _23584_/Q _22548_/Q _22352_/Q _13275_/A _11527_/X vssd1 vssd1 vccd1
+ vccd1 _13062_/B sky130_fd_sc_hd__mux4_1
X_22259_ _21327_/X _22258_/X _22257_/X _14556_/D vssd1 vssd1 vccd1 vccd1 _22260_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_322_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12012_ _12141_/A vssd1 vssd1 vccd1 vccd1 _12852_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_293_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23568_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16820_ _16819_/X _22522_/Q _16829_/S vssd1 vssd1 vccd1 vccd1 _16821_/A sky130_fd_sc_hd__mux2_1
XFILLER_305_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16751_ _16751_/A vssd1 vssd1 vccd1 vccd1 _22502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_281_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13963_ _13963_/A _13965_/B vssd1 vssd1 vccd1 vccd1 _13963_/Y sky130_fd_sc_hd__nor2_1
XFILLER_293_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15702_ _21856_/A _15701_/C _21888_/A vssd1 vssd1 vccd1 vccd1 _21868_/C sky130_fd_sc_hd__a21oi_2
X_19470_ _19470_/A vssd1 vssd1 vccd1 vccd1 _23390_/D sky130_fd_sc_hd__clkbuf_1
X_12914_ _13493_/A _13493_/B vssd1 vssd1 vccd1 vccd1 _12916_/A sky130_fd_sc_hd__and2_1
XFILLER_234_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16682_ input42/X _16680_/A _19987_/A vssd1 vssd1 vccd1 vccd1 _16808_/B sky130_fd_sc_hd__a21oi_1
X_13894_ _23913_/Q vssd1 vssd1 vccd1 vccd1 _13895_/A sky130_fd_sc_hd__inv_2
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18421_ _18441_/A _18427_/C vssd1 vssd1 vccd1 vccd1 _18421_/Y sky130_fd_sc_hd__nor2_1
X_12845_ _22284_/Q _23100_/Q _23516_/Q _22445_/Q _12843_/X _12844_/X vssd1 vssd1 vccd1
+ vccd1 _12846_/B sky130_fd_sc_hd__mux4_1
X_15633_ _15901_/A vssd1 vssd1 vccd1 vccd1 _15633_/X sky130_fd_sc_hd__buf_2
XFILLER_62_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _18360_/A _18357_/C vssd1 vssd1 vccd1 vccd1 _18352_/Y sky130_fd_sc_hd__nor2_1
XFILLER_203_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _12843_/A vssd1 vssd1 vccd1 vccd1 _12776_/X sky130_fd_sc_hd__buf_4
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _15564_/A _15564_/B vssd1 vssd1 vccd1 vccd1 _15564_/Y sky130_fd_sc_hd__nand2_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17242_/A _17296_/X _17302_/X _16997_/X vssd1 vssd1 vccd1 vccd1 _17303_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_202_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ _15440_/A vssd1 vssd1 vccd1 vccd1 _14516_/A sky130_fd_sc_hd__buf_2
X_11727_ _12260_/A _11727_/B _11727_/C vssd1 vssd1 vccd1 vccd1 _13803_/A sky130_fd_sc_hd__nor3_4
XFILLER_348_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18283_ _18286_/A _18286_/C _18175_/X vssd1 vssd1 vccd1 vccd1 _18283_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_148_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ _15495_/A vssd1 vssd1 vccd1 vccd1 _15718_/B sky130_fd_sc_hd__buf_2
XFILLER_187_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17234_ _15864_/X _17233_/X _17234_/S vssd1 vssd1 vccd1 vccd1 _17234_/X sky130_fd_sc_hd__mux2_1
XFILLER_317_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11658_ _11631_/X _11639_/X _11641_/X _11656_/X _11657_/X vssd1 vssd1 vccd1 vccd1
+ _11685_/B sky130_fd_sc_hd__a311o_1
X_14446_ _14467_/B _14446_/B _14467_/C vssd1 vssd1 vccd1 vccd1 _20770_/A sky130_fd_sc_hd__or3b_4
XFILLER_187_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17165_ _17167_/A _17156_/X _17164_/X _16996_/X _17109_/A vssd1 vssd1 vccd1 vccd1
+ _17165_/X sky130_fd_sc_hd__o221a_4
X_14377_ _14949_/S _14375_/Y _14376_/X vssd1 vssd1 vccd1 vccd1 _14377_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11589_ _12350_/A vssd1 vssd1 vccd1 vccd1 _11590_/A sky130_fd_sc_hd__buf_4
XFILLER_128_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_346_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13328_ _13328_/A _13604_/A vssd1 vssd1 vccd1 vccd1 _13632_/A sky130_fd_sc_hd__nor2_4
XFILLER_6_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16116_ _15752_/X _16113_/X _16115_/Y _16005_/X vssd1 vssd1 vccd1 vccd1 _16116_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_127_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_1_wb_clk_i clkbuf_2_2_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_6_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17096_ _14538_/X _17095_/X _17116_/S vssd1 vssd1 vccd1 vccd1 _17096_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_346_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_332_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16047_ _16045_/X _22139_/B _16047_/S vssd1 vssd1 vccd1 vccd1 _18859_/A sky130_fd_sc_hd__mux2_4
X_13259_ _13259_/A _13259_/B vssd1 vssd1 vccd1 vccd1 _13259_/Y sky130_fd_sc_hd__nor2_1
XFILLER_331_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19806_ _19828_/A vssd1 vssd1 vccd1 vccd1 _19815_/S sky130_fd_sc_hd__buf_4
X_17998_ input6/X input281/X _18005_/S vssd1 vssd1 vccd1 vccd1 _17998_/X sky130_fd_sc_hd__mux2_1
XFILLER_215_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19737_ _19217_/X _23509_/Q _19743_/S vssd1 vssd1 vccd1 vccd1 _19738_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16949_ _16949_/A vssd1 vssd1 vccd1 vccd1 _17244_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19668_ _19668_/A vssd1 vssd1 vccd1 vccd1 _23478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18619_ _16908_/X _23042_/Q _18619_/S vssd1 vssd1 vccd1 vccd1 _18620_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19599_ _23448_/Q _19226_/A _19599_/S vssd1 vssd1 vccd1 vccd1 _19600_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21630_ _21630_/A _23756_/Q vssd1 vssd1 vccd1 vccd1 _21630_/X sky130_fd_sc_hd__and2_1
XFILLER_178_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_339_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21561_ _21813_/A _21559_/Y _21560_/X _23789_/Q vssd1 vssd1 vccd1 vccd1 _21561_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_178_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23300_ _23556_/CLK _23300_/D vssd1 vssd1 vccd1 vccd1 _23300_/Q sky130_fd_sc_hd__dfxtp_1
X_20512_ _22710_/Q vssd1 vssd1 vccd1 vccd1 _20523_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_327_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_308_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21492_ _23819_/Q _23753_/Q vssd1 vssd1 vccd1 vccd1 _21494_/A sky130_fd_sc_hd__or2_1
XFILLER_193_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23231_ _23423_/CLK _23231_/D vssd1 vssd1 vccd1 vccd1 _23231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_308_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20443_ _20639_/A _20428_/X _20442_/X _20433_/X vssd1 vssd1 vccd1 vccd1 _23696_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23162_ _23420_/CLK _23162_/D vssd1 vssd1 vccd1 vccd1 _23162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_335_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20374_ _20374_/A _20400_/B vssd1 vssd1 vccd1 vccd1 _20376_/B sky130_fd_sc_hd__or2_1
XFILLER_133_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_7118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22113_ _22114_/A _22119_/A vssd1 vssd1 vccd1 vccd1 _22115_/A sky130_fd_sc_hd__nor2_1
XTAP_7129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23093_ _23349_/CLK _23093_/D vssd1 vssd1 vccd1 vccd1 _23093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_311_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_288_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22044_ _22044_/A vssd1 vssd1 vccd1 vccd1 _22044_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_350_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_304_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_349_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_291_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22946_ _23602_/CLK _22946_/D vssd1 vssd1 vccd1 vccd1 _22946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22877_ _23009_/CLK _22877_/D vssd1 vssd1 vccd1 vccd1 _22877_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_203_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12630_ _12998_/A _12630_/B vssd1 vssd1 vccd1 vccd1 _12630_/Y sky130_fd_sc_hd__nor2_1
XPHY_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_157_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23700_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21828_ _21828_/A _21828_/B vssd1 vssd1 vccd1 vccd1 _21828_/Y sky130_fd_sc_hd__xnor2_1
XPHY_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12561_ _12570_/A _12561_/B vssd1 vssd1 vccd1 vccd1 _12561_/X sky130_fd_sc_hd__or2_1
X_21759_ _23827_/Q _21758_/Y _22214_/S vssd1 vssd1 vccd1 vccd1 _21760_/B sky130_fd_sc_hd__mux2_1
XPHY_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_358_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_318_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11512_ _23908_/Q vssd1 vssd1 vccd1 vccd1 _14179_/A sky130_fd_sc_hd__buf_6
X_14300_ _12166_/X _12809_/B _14329_/S vssd1 vssd1 vccd1 vccd1 _14300_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15280_ _15280_/A vssd1 vssd1 vccd1 vccd1 _21594_/A sky130_fd_sc_hd__buf_6
XFILLER_211_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12492_ _12485_/X _12487_/X _12489_/X _12491_/X _11272_/A vssd1 vssd1 vccd1 vccd1
+ _12493_/C sky130_fd_sc_hd__a221o_1
XFILLER_345_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14231_ _14231_/A vssd1 vssd1 vccd1 vccd1 _14232_/A sky130_fd_sc_hd__clkbuf_2
X_11443_ _21077_/C _11440_/X _11502_/A vssd1 vssd1 vccd1 vccd1 _11443_/X sky130_fd_sc_hd__a21o_1
X_23429_ _23527_/CLK _23429_/D vssd1 vssd1 vccd1 vccd1 _23429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_314_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14162_ _14164_/A vssd1 vssd1 vccd1 vccd1 _16929_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_313_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11374_ _23898_/Q vssd1 vssd1 vccd1 vccd1 _11375_/A sky130_fd_sc_hd__buf_4
XFILLER_124_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_341_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_314_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13113_ _13225_/A vssd1 vssd1 vccd1 vccd1 _13117_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_180_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18970_ _19016_/S vssd1 vssd1 vccd1 vccd1 _18979_/S sky130_fd_sc_hd__buf_4
X_14093_ _14093_/A vssd1 vssd1 vccd1 vccd1 _14093_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_302_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17921_ _17971_/A vssd1 vssd1 vccd1 vccd1 _17956_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_301_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13044_ _12816_/X _13036_/Y _13039_/Y _13041_/Y _13043_/Y vssd1 vssd1 vccd1 vccd1
+ _13044_/X sky130_fd_sc_hd__o32a_1
XFILLER_332_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17852_ _17852_/A vssd1 vssd1 vccd1 vccd1 _22797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16803_ _22518_/Q _16729_/A _16730_/A input34/X vssd1 vssd1 vccd1 vccd1 _16804_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_208_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_293_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17783_ _22767_/Q _17617_/X _17787_/S vssd1 vssd1 vccd1 vccd1 _17784_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14995_ _23754_/Q _14911_/X _14913_/X _14993_/X _14994_/X vssd1 vssd1 vccd1 vccd1
+ _14995_/X sky130_fd_sc_hd__a221o_1
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19522_ _19522_/A vssd1 vssd1 vccd1 vccd1 _23413_/D sky130_fd_sc_hd__clkbuf_1
X_16734_ _22498_/Q _16729_/X _16730_/X input12/X vssd1 vssd1 vccd1 vccd1 _16735_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13946_ _13918_/X _15256_/A _13945_/Y _13924_/X vssd1 vssd1 vccd1 vccd1 _14097_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_235_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19453_ _23383_/Q _18830_/X _19455_/S vssd1 vssd1 vccd1 vccd1 _19454_/A sky130_fd_sc_hd__mux2_1
XFILLER_250_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16665_ _22479_/Q _16287_/X _16673_/S vssd1 vssd1 vccd1 vccd1 _16666_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13877_ _13874_/X _13875_/X _13876_/X vssd1 vssd1 vccd1 vccd1 _14069_/C sky130_fd_sc_hd__o21ai_4
XFILLER_223_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18404_ _22962_/Q _18402_/B _18403_/Y vssd1 vssd1 vccd1 vccd1 _22962_/D sky130_fd_sc_hd__o21a_1
X_15616_ _15616_/A vssd1 vssd1 vccd1 vccd1 _17159_/A sky130_fd_sc_hd__buf_6
X_19384_ _19384_/A vssd1 vssd1 vccd1 vccd1 _23352_/D sky130_fd_sc_hd__clkbuf_1
X_12828_ _12687_/X _12818_/Y _12822_/Y _12824_/Y _12827_/Y vssd1 vssd1 vccd1 vccd1
+ _12828_/X sky130_fd_sc_hd__o32a_1
X_16596_ _16596_/A vssd1 vssd1 vccd1 vccd1 _22448_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18335_ _18360_/A _18341_/C vssd1 vssd1 vccd1 vccd1 _18335_/Y sky130_fd_sc_hd__nor2_1
XFILLER_231_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15547_ _22929_/Q _15000_/A _15001_/A _22961_/Q vssd1 vssd1 vccd1 vccd1 _15547_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12759_ _12759_/A vssd1 vssd1 vccd1 vccd1 _12886_/A sky130_fd_sc_hd__buf_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_336_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18266_ _22914_/Q _22915_/Q _22916_/Q _22917_/Q vssd1 vssd1 vccd1 vccd1 _18279_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_202_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15478_ _15478_/A vssd1 vssd1 vccd1 vccd1 _15478_/X sky130_fd_sc_hd__buf_2
XFILLER_348_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17217_ _17167_/X _17210_/X _17216_/X _17176_/X vssd1 vssd1 vccd1 vccd1 _17217_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_352_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14429_ _15558_/A vssd1 vssd1 vccd1 vccd1 _14897_/A sky130_fd_sc_hd__clkbuf_2
X_18197_ _18188_/A _18118_/X _18186_/B _18196_/X _18192_/X vssd1 vssd1 vccd1 vccd1
+ _22893_/D sky130_fd_sc_hd__o221a_1
XFILLER_128_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_317_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_317_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_293_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17148_ _14167_/X _15560_/Y _17172_/B _17147_/Y vssd1 vssd1 vccd1 vccd1 _17148_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_305_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_289_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17079_ _17073_/X _17077_/X _16968_/X _17078_/X vssd1 vssd1 vccd1 vccd1 _17079_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20090_ _23637_/Q _23636_/Q _20090_/C _20090_/D vssd1 vssd1 vccd1 vccd1 _20098_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_131_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22800_ _23068_/CLK _22800_/D vssd1 vssd1 vccd1 vccd1 _22800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23780_ _23861_/CLK _23780_/D vssd1 vssd1 vccd1 vccd1 _23780_/Q sky130_fd_sc_hd__dfxtp_1
X_20992_ _20543_/A _20988_/X _20991_/X _20978_/X vssd1 vssd1 vccd1 vccd1 _23813_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22731_ _23575_/CLK _22731_/D vssd1 vssd1 vccd1 vccd1 _22731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_281_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22662_ _22695_/CLK _22662_/D vssd1 vssd1 vccd1 vccd1 _22662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21613_ _21613_/A vssd1 vssd1 vccd1 vccd1 _21613_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22593_ _22977_/CLK _22593_/D vssd1 vssd1 vccd1 vccd1 _22593_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_222_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21544_ _21485_/A _21485_/B _21452_/A _21452_/B vssd1 vssd1 vccd1 vccd1 _21544_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_328_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21475_ _21829_/B _21472_/X _21473_/Y _21474_/Y _21327_/A vssd1 vssd1 vccd1 vccd1
+ _21476_/B sky130_fd_sc_hd__a311o_1
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23214_ _23502_/CLK _23214_/D vssd1 vssd1 vccd1 vccd1 _23214_/Q sky130_fd_sc_hd__dfxtp_1
X_20426_ _23690_/Q _20429_/B vssd1 vssd1 vccd1 vccd1 _20426_/X sky130_fd_sc_hd__or2_1
XFILLER_181_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_323_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_351_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23145_ _23561_/CLK _23145_/D vssd1 vssd1 vccd1 vccd1 _23145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20357_ _23677_/Q _20391_/B vssd1 vssd1 vccd1 vccd1 _20357_/X sky130_fd_sc_hd__or2_1
XFILLER_135_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23076_ _23577_/CLK _23076_/D vssd1 vssd1 vccd1 vccd1 _23076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11090_ _13775_/B _20148_/A _11090_/C vssd1 vssd1 vccd1 vccd1 _12544_/B sky130_fd_sc_hd__nor3_2
XFILLER_311_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20288_ _15560_/Y _20215_/X _20289_/B vssd1 vssd1 vccd1 vccd1 _20288_/X sky130_fd_sc_hd__o21a_1
XTAP_5502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22027_ _22000_/B _22002_/B _22000_/A vssd1 vssd1 vccd1 vccd1 _22031_/A sky130_fd_sc_hd__a21bo_1
XTAP_6269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13800_ _13790_/X _13847_/A _13799_/X vssd1 vssd1 vccd1 vccd1 _13801_/B sky130_fd_sc_hd__a21oi_4
X_11992_ _23220_/Q _23188_/Q _23156_/Q _23124_/Q _12709_/A _11669_/X vssd1 vssd1 vccd1
+ vccd1 _11993_/B sky130_fd_sc_hd__mux4_2
XFILLER_290_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14780_ _14774_/Y _14779_/Y _14855_/A vssd1 vssd1 vccd1 vccd1 _14780_/X sky130_fd_sc_hd__mux2_1
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13731_ _13884_/A vssd1 vssd1 vccd1 vccd1 _21191_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_290_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22929_ _22929_/CLK _22929_/D vssd1 vssd1 vccd1 vccd1 _22929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16450_ _16450_/A vssd1 vssd1 vccd1 vccd1 _22385_/D sky130_fd_sc_hd__clkbuf_1
X_13662_ _22603_/Q _13662_/B _13662_/C vssd1 vssd1 vccd1 vccd1 _13670_/A sky130_fd_sc_hd__or3_1
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _23761_/Q _14910_/A _14912_/A _15399_/X _15400_/X vssd1 vssd1 vccd1 vccd1
+ _15401_/X sky130_fd_sc_hd__a221o_1
X_12613_ _13943_/A _13343_/B _13380_/A _13371_/A vssd1 vssd1 vccd1 vccd1 _12613_/X
+ sky130_fd_sc_hd__or4_2
X_16381_ _16197_/X _22356_/Q _16381_/S vssd1 vssd1 vccd1 vccd1 _16382_/A sky130_fd_sc_hd__mux2_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _13593_/A vssd1 vssd1 vccd1 vccd1 _13594_/A sky130_fd_sc_hd__clkbuf_2
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18120_ _21220_/A vssd1 vssd1 vccd1 vccd1 _18245_/A sky130_fd_sc_hd__clkbuf_4
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_346_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15332_ _15332_/A _15432_/B vssd1 vssd1 vccd1 vccd1 _15332_/Y sky130_fd_sc_hd__nand2_2
X_12544_ _23886_/Q _12544_/B vssd1 vssd1 vccd1 vccd1 _12544_/X sky130_fd_sc_hd__and2_1
XFILLER_345_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_346_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18051_ _18051_/A vssd1 vssd1 vccd1 vccd1 _18051_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_185_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15263_ _23726_/Q _23856_/Q _16022_/S vssd1 vssd1 vccd1 vccd1 _15263_/X sky130_fd_sc_hd__mux2_1
X_12475_ _12475_/A vssd1 vssd1 vccd1 vccd1 _12475_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17002_ _22710_/Q vssd1 vssd1 vccd1 vccd1 _20517_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_345_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11426_ _13259_/A _11425_/X _11135_/A vssd1 vssd1 vccd1 vccd1 _11426_/Y sky130_fd_sc_hd__o21ai_1
X_14214_ _14569_/A vssd1 vssd1 vccd1 vccd1 _14215_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_333_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15194_ _15192_/Y _15193_/X _15020_/S _15127_/Y vssd1 vssd1 vccd1 vccd1 _15194_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_138_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_54_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _22632_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14145_ _23012_/Q _14700_/C vssd1 vssd1 vccd1 vccd1 _14211_/B sky130_fd_sc_hd__nand2_1
XFILLER_126_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11357_ _23898_/Q _23897_/Q vssd1 vssd1 vccd1 vccd1 _11457_/D sky130_fd_sc_hd__or2_4
XFILLER_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_314_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14076_ _14049_/X _13888_/B _14009_/X _22811_/Q vssd1 vssd1 vccd1 vccd1 _14076_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_98_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18953_ _16822_/X _23175_/Q _18957_/S vssd1 vssd1 vccd1 vccd1 _18954_/A sky130_fd_sc_hd__mux2_1
XFILLER_302_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_298_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11288_ _11288_/A vssd1 vssd1 vccd1 vccd1 _11288_/X sky130_fd_sc_hd__buf_2
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17904_ _22813_/Q _17894_/X _17903_/X input253/X _17899_/X vssd1 vssd1 vccd1 vccd1
+ _17904_/X sky130_fd_sc_hd__a221o_1
X_13027_ _13601_/A _13323_/B _13026_/Y vssd1 vssd1 vccd1 vccd1 _13027_/X sky130_fd_sc_hd__o21a_1
XFILLER_295_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18884_ _18884_/A vssd1 vssd1 vccd1 vccd1 _23144_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_343_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17835_ _22790_/Q _17588_/X _17837_/S vssd1 vssd1 vccd1 vccd1 _17836_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17766_ _17766_/A vssd1 vssd1 vccd1 vccd1 _22759_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14978_ _15161_/A _21421_/B vssd1 vssd1 vccd1 vccd1 _14978_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19505_ _19194_/X _23406_/Q _19505_/S vssd1 vssd1 vccd1 vccd1 _19506_/A sky130_fd_sc_hd__mux2_1
XFILLER_263_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16717_ _16723_/A _16717_/B vssd1 vssd1 vccd1 vccd1 _16718_/A sky130_fd_sc_hd__or2_1
X_13929_ _23918_/Q vssd1 vssd1 vccd1 vccd1 _21522_/A sky130_fd_sc_hd__buf_2
X_17697_ _17697_/A vssd1 vssd1 vccd1 vccd1 _22728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_410 _14029_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_421 _14065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19436_ _23375_/Q _18804_/X _19444_/S vssd1 vssd1 vccd1 vccd1 _19437_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_432 _23881_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16648_ _16648_/A vssd1 vssd1 vccd1 vccd1 _22471_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_443 _23918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_454 wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_465 _21327_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_476 _21444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19367_ _19367_/A vssd1 vssd1 vccd1 vccd1 _23344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_487 _13964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16579_ _15749_/X _22441_/Q _16579_/S vssd1 vssd1 vccd1 vccd1 _16580_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_498 _14722_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_309_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18318_ _22932_/Q _18315_/C _18317_/Y vssd1 vssd1 vccd1 vccd1 _22932_/D sky130_fd_sc_hd__o21a_1
XFILLER_188_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_349_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19298_ _19207_/X _23314_/Q _19300_/S vssd1 vssd1 vccd1 vccd1 _19299_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_337_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18249_ _22911_/Q _18253_/B vssd1 vssd1 vccd1 vccd1 _18249_/X sky130_fd_sc_hd__or2_1
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_318_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21260_ _14393_/X _15794_/X _21260_/S vssd1 vssd1 vccd1 vccd1 _21261_/B sky130_fd_sc_hd__mux2_1
XFILLER_237_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_305_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20211_ _23658_/Q _20223_/B vssd1 vssd1 vccd1 vccd1 _20211_/X sky130_fd_sc_hd__or2_1
XFILLER_274_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21191_ _21191_/A _21191_/B vssd1 vssd1 vccd1 vccd1 _21192_/A sky130_fd_sc_hd__nand2_1
XFILLER_116_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20142_ _20160_/A _20986_/B vssd1 vssd1 vccd1 vccd1 _20143_/A sky130_fd_sc_hd__or2_2
XFILLER_277_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20073_ _23632_/Q _20069_/B _20072_/Y vssd1 vssd1 vccd1 vccd1 _23632_/D sky130_fd_sc_hd__o21a_1
XFILLER_253_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23901_ _23903_/CLK _23901_/D vssd1 vssd1 vccd1 vccd1 _23901_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23832_ _23832_/CLK _23832_/D vssd1 vssd1 vccd1 vccd1 _23832_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23763_ _23804_/CLK _23763_/D vssd1 vssd1 vccd1 vccd1 _23763_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_260_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20975_ _22139_/A _20966_/X _20747_/B _20970_/X vssd1 vssd1 vccd1 vccd1 _20975_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22714_ _23496_/CLK _22714_/D vssd1 vssd1 vccd1 vccd1 _22714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23694_ _23696_/CLK _23694_/D vssd1 vssd1 vccd1 vccd1 _23694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22645_ _23588_/CLK _22645_/D vssd1 vssd1 vccd1 vccd1 _22645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22576_ _23643_/CLK _22576_/D vssd1 vssd1 vccd1 vccd1 _22576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21527_ _21542_/A _21487_/B _21546_/A vssd1 vssd1 vccd1 vccd1 _21528_/B sky130_fd_sc_hd__a21oi_1
XFILLER_127_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12260_ _12260_/A _12260_/B _12260_/C vssd1 vssd1 vccd1 vccd1 _13724_/A sky130_fd_sc_hd__or3_4
X_21458_ _23818_/Q _23752_/Q vssd1 vssd1 vccd1 vccd1 _21460_/A sky130_fd_sc_hd__nor2_1
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_342_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ _13259_/A _11199_/Y _11202_/Y _11210_/Y vssd1 vssd1 vccd1 vccd1 _11211_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20409_ _20409_/A _21084_/B vssd1 vssd1 vccd1 vccd1 _20470_/A sky130_fd_sc_hd__nor2_4
XFILLER_294_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12191_ _23899_/Q vssd1 vssd1 vccd1 vccd1 _12535_/S sky130_fd_sc_hd__clkbuf_4
X_21389_ _21425_/A _21425_/B vssd1 vssd1 vccd1 vccd1 _21391_/A sky130_fd_sc_hd__nor2_1
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23128_ _23511_/CLK _23128_/D vssd1 vssd1 vccd1 vccd1 _23128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_311_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11142_ _12985_/A vssd1 vssd1 vccd1 vccd1 _13084_/A sky130_fd_sc_hd__clkbuf_2
XTAP_6000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_311_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_295_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15950_ _22939_/Q vssd1 vssd1 vccd1 vccd1 _15950_/X sky130_fd_sc_hd__buf_2
XTAP_5310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23059_ _23571_/CLK _23059_/D vssd1 vssd1 vccd1 vccd1 _23059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11073_ _14172_/C vssd1 vssd1 vccd1 vccd1 _13440_/C sky130_fd_sc_hd__buf_4
XFILLER_277_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput110 dout1[12] vssd1 vssd1 vccd1 vccd1 input110/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput121 dout1[22] vssd1 vssd1 vccd1 vccd1 input121/X sky130_fd_sc_hd__clkbuf_1
XTAP_5332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14901_ _14901_/A vssd1 vssd1 vccd1 vccd1 _14901_/X sky130_fd_sc_hd__clkbuf_2
Xinput132 dout1[32] vssd1 vssd1 vccd1 vccd1 input132/X sky130_fd_sc_hd__buf_2
XTAP_6088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput143 dout1[42] vssd1 vssd1 vccd1 vccd1 input143/X sky130_fd_sc_hd__buf_2
XTAP_6099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput154 dout1[52] vssd1 vssd1 vccd1 vccd1 input154/X sky130_fd_sc_hd__buf_2
XTAP_5365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15881_ _23772_/Q _14911_/X _14913_/X _15879_/X _15880_/X vssd1 vssd1 vccd1 vccd1
+ _15881_/X sky130_fd_sc_hd__a221o_2
XTAP_5376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput165 dout1[62] vssd1 vssd1 vccd1 vccd1 input165/X sky130_fd_sc_hd__buf_2
XFILLER_263_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ _18846_/A vssd1 vssd1 vccd1 vccd1 _17620_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput176 irq[14] vssd1 vssd1 vccd1 vccd1 _20518_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14832_ _22490_/Q _13692_/A _14247_/X _14831_/X _14072_/A vssd1 vssd1 vccd1 vccd1
+ _14832_/X sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_172_wb_clk_i _23917_/CLK vssd1 vssd1 vccd1 vccd1 _23776_/CLK sky130_fd_sc_hd__clkbuf_16
Xinput187 jtag_tck vssd1 vssd1 vccd1 vccd1 _18138_/A sky130_fd_sc_hd__buf_12
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput198 localMemory_wb_adr_i[17] vssd1 vssd1 vccd1 vccd1 input198/X sky130_fd_sc_hd__clkbuf_1
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_292_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_291_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_313_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_101_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23584_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_217_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _22679_/Q _17550_/X _17560_/S vssd1 vssd1 vccd1 vccd1 _17552_/A sky130_fd_sc_hd__mux2_1
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14763_ _14848_/A vssd1 vssd1 vccd1 vccd1 _15491_/S sky130_fd_sc_hd__clkbuf_2
X_11975_ _12056_/A _11975_/B vssd1 vssd1 vccd1 vccd1 _11975_/Y sky130_fd_sc_hd__nor2_1
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16502_ _15749_/X _22408_/Q _16502_/S vssd1 vssd1 vccd1 vccd1 _16503_/A sky130_fd_sc_hd__mux2_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13714_ _13718_/A _13714_/B _13718_/D vssd1 vssd1 vccd1 vccd1 _14015_/C sky130_fd_sc_hd__and3_4
XFILLER_44_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17482_ _17482_/A vssd1 vssd1 vccd1 vccd1 _22649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14694_ _14570_/X _21204_/A _14693_/Y _14521_/A vssd1 vssd1 vccd1 vccd1 _14695_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_205_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19221_ _19220_/X _23286_/Q _19227_/S vssd1 vssd1 vccd1 vccd1 _19222_/A sky130_fd_sc_hd__mux2_1
X_16433_ _16433_/A vssd1 vssd1 vccd1 vccd1 _22377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13645_ _13948_/A _13948_/B _11940_/A vssd1 vssd1 vccd1 vccd1 _13646_/B sky130_fd_sc_hd__a21oi_2
XFILLER_72_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19152_ _19152_/A vssd1 vssd1 vccd1 vccd1 _23263_/D sky130_fd_sc_hd__clkbuf_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_318_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16364_ _15898_/X _22348_/Q _16366_/S vssd1 vssd1 vccd1 vccd1 _16365_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_346_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13576_ _13581_/A _22087_/A _13490_/X _13575_/Y vssd1 vssd1 vccd1 vccd1 _13981_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_358_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _22872_/Q _18096_/X _18102_/X _18090_/X vssd1 vssd1 vccd1 vccd1 _22872_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_297_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15315_ _23921_/Q _15316_/B vssd1 vssd1 vccd1 vccd1 _15376_/C sky130_fd_sc_hd__and2_1
XFILLER_347_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19083_ _19083_/A vssd1 vssd1 vccd1 vccd1 _23233_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12527_ _12534_/A _12526_/X _11127_/A vssd1 vssd1 vccd1 vccd1 _12527_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_338_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16295_ _22320_/Q _16294_/X _16301_/S vssd1 vssd1 vccd1 vccd1 _16296_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18034_ _22850_/Q _18016_/X _18033_/X _18029_/X vssd1 vssd1 vccd1 vccd1 _22850_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_334_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15246_ _14580_/Y _15181_/X _15183_/X _15245_/Y vssd1 vssd1 vccd1 vccd1 _21227_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_338_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12458_ _12458_/A _12458_/B vssd1 vssd1 vccd1 vccd1 _12458_/Y sky130_fd_sc_hd__nand2_1
XFILLER_274_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_315_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11409_ _13212_/A vssd1 vssd1 vccd1 vccd1 _13273_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_315_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15177_ _14815_/B _15995_/A _15174_/X _15176_/X vssd1 vssd1 vccd1 vccd1 _15187_/B
+ sky130_fd_sc_hd__o211a_2
X_12389_ _12378_/A _12388_/X _11346_/A vssd1 vssd1 vccd1 vccd1 _12389_/X sky130_fd_sc_hd__o21a_1
XFILLER_342_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14128_ _15425_/A _20532_/C vssd1 vssd1 vccd1 vccd1 _14128_/Y sky130_fd_sc_hd__nor2_1
X_19985_ _23608_/Q _23607_/Q _19985_/C _19985_/D vssd1 vssd1 vccd1 vccd1 _20003_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_299_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18936_ _23168_/Q _18859_/X _18940_/S vssd1 vssd1 vccd1 vccd1 _18937_/A sky130_fd_sc_hd__mux2_1
X_14059_ _14064_/A _14066_/B _14059_/C vssd1 vssd1 vccd1 vccd1 _14059_/X sky130_fd_sc_hd__or3_1
XFILLER_97_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_290_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18867_ _18867_/A vssd1 vssd1 vccd1 vccd1 _23138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_294_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17818_ _22782_/Q _17562_/X _17826_/S vssd1 vssd1 vccd1 vccd1 _17819_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18798_ _18798_/A vssd1 vssd1 vccd1 vccd1 _18798_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_345_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17749_ _17749_/A vssd1 vssd1 vccd1 vccd1 _22751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_345_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20760_ _21079_/B _20642_/A _20662_/X vssd1 vssd1 vccd1 vccd1 _20760_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_240 _15230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_251 _17122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19419_ _19419_/A vssd1 vssd1 vccd1 vccd1 _23367_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_262 _15651_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_273 _15692_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20691_ _21153_/A _20744_/B vssd1 vssd1 vccd1 vccd1 _20695_/B sky130_fd_sc_hd__nor2_4
XINSDIODE2_284 _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_338_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_295 _15990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22430_ _23565_/CLK _22430_/D vssd1 vssd1 vccd1 vccd1 _22430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22361_ _23527_/CLK _22361_/D vssd1 vssd1 vccd1 vccd1 _22361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21312_ _21613_/A vssd1 vssd1 vccd1 vccd1 _21346_/A sky130_fd_sc_hd__buf_2
X_22292_ _23556_/CLK _22292_/D vssd1 vssd1 vccd1 vccd1 _22292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_324_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21243_ _21243_/A vssd1 vssd1 vccd1 vccd1 _21274_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21174_ _21083_/A _20509_/B _21150_/X vssd1 vssd1 vccd1 vccd1 _21174_/X sky130_fd_sc_hd__a21o_1
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_321_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20125_ _23648_/Q _20131_/D vssd1 vssd1 vccd1 vccd1 _20127_/B sky130_fd_sc_hd__nor2_1
XFILLER_259_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_293_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20056_ _20066_/A _23627_/Q _20056_/C _20056_/D vssd1 vssd1 vccd1 vccd1 _20076_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_292_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23815_ _23856_/CLK _23815_/D vssd1 vssd1 vccd1 vccd1 _23815_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11750_/Y _11752_/Y _11757_/Y _11759_/Y _11657_/A vssd1 vssd1 vccd1 vccd1
+ _11761_/C sky130_fd_sc_hd__o221a_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20958_ _23802_/Q _20953_/X _20957_/X _20948_/X vssd1 vssd1 vccd1 vccd1 _23802_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23746_ _23915_/CLK _23746_/D vssd1 vssd1 vccd1 vccd1 _23746_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11691_ _13536_/A _11691_/B vssd1 vssd1 vccd1 vccd1 _13532_/A sky130_fd_sc_hd__xnor2_4
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23677_ _23706_/CLK _23677_/D vssd1 vssd1 vccd1 vccd1 _23677_/Q sky130_fd_sc_hd__dfxtp_1
X_20889_ _23780_/Q _20786_/B _20888_/X _20788_/X vssd1 vssd1 vccd1 vccd1 _23780_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_201_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_329_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13430_ _21518_/A vssd1 vssd1 vccd1 vccd1 _21336_/A sky130_fd_sc_hd__buf_2
X_22628_ _23571_/CLK _22628_/D vssd1 vssd1 vccd1 vccd1 _22628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_325_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13361_ _12546_/A _13361_/B vssd1 vssd1 vccd1 vccd1 _14290_/A sky130_fd_sc_hd__and2b_4
X_22559_ _22977_/CLK _22559_/D vssd1 vssd1 vccd1 vccd1 _22559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_344_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15100_ _14804_/A _15051_/Y _15099_/Y _14698_/X vssd1 vssd1 vccd1 vccd1 _15100_/X
+ sky130_fd_sc_hd__a211o_1
X_12312_ _23904_/Q _11910_/A _12415_/S vssd1 vssd1 vccd1 vccd1 _12312_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_127_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13292_ _22482_/Q _22642_/Q _22321_/Q _23457_/Q _13275_/X _13276_/X vssd1 vssd1 vccd1
+ vccd1 _13292_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16080_ _15923_/A _16074_/X _16079_/X _15480_/A vssd1 vssd1 vccd1 vccd1 _16080_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_343_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15031_ _22500_/Q _14219_/X _14238_/X _15030_/X _14242_/X vssd1 vssd1 vccd1 vccd1
+ _15031_/Y sky130_fd_sc_hd__o221ai_4
X_12243_ _12423_/A _12243_/B vssd1 vssd1 vccd1 vccd1 _12243_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12174_ _12567_/A _12174_/B vssd1 vssd1 vccd1 vccd1 _12174_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_323_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11125_ _13210_/A vssd1 vssd1 vccd1 vccd1 _13765_/A sky130_fd_sc_hd__clkbuf_16
X_19770_ _19770_/A vssd1 vssd1 vccd1 vccd1 _23524_/D sky130_fd_sc_hd__clkbuf_1
X_16982_ _17250_/A vssd1 vssd1 vccd1 vccd1 _17163_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_150_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_296_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18721_ _18767_/S vssd1 vssd1 vccd1 vccd1 _18730_/S sky130_fd_sc_hd__buf_4
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15933_ _23002_/Q _16084_/A _16085_/A input231/X vssd1 vssd1 vccd1 vccd1 _22067_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18652_ _23056_/Q _17582_/X _18658_/S vssd1 vssd1 vccd1 vccd1 _18653_/A sky130_fd_sc_hd__mux2_1
XFILLER_329_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _15864_/A vssd1 vssd1 vccd1 vccd1 _15864_/X sky130_fd_sc_hd__buf_6
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17603_ _17603_/A vssd1 vssd1 vccd1 vccd1 _22695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ _21335_/B _14815_/B _14815_/C vssd1 vssd1 vccd1 vccd1 _21482_/A sky130_fd_sc_hd__and3_2
X_18583_ _18583_/A vssd1 vssd1 vccd1 vccd1 _23025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795_ _13605_/Y _15580_/B _15636_/X vssd1 vssd1 vccd1 vccd1 _15797_/A sky130_fd_sc_hd__a21oi_1
XFILLER_64_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ _22673_/Q _16294_/X _17538_/S vssd1 vssd1 vccd1 vccd1 _17535_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14746_ _23687_/Q _14738_/X _14739_/X _14744_/X _14745_/Y vssd1 vssd1 vccd1 vccd1
+ _14746_/X sky130_fd_sc_hd__a221o_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11958_ _12119_/S vssd1 vssd1 vccd1 vccd1 _12680_/A sky130_fd_sc_hd__buf_4
XFILLER_205_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17465_ _22643_/Q _16300_/X _17465_/S vssd1 vssd1 vccd1 vccd1 _17466_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14677_ _14676_/A _14674_/X _14676_/Y _14259_/X vssd1 vssd1 vccd1 vccd1 _14677_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_189_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11889_ _23213_/Q _23181_/Q _23149_/Q _23117_/Q _12120_/S _11696_/X vssd1 vssd1 vccd1
+ vccd1 _11890_/B sky130_fd_sc_hd__mux4_1
XFILLER_60_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19204_ _19204_/A vssd1 vssd1 vccd1 vccd1 _19204_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16416_ _15474_/X _22370_/Q _16418_/S vssd1 vssd1 vccd1 vccd1 _16417_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13628_ _13965_/A _13964_/A _13963_/A _13628_/D vssd1 vssd1 vccd1 vccd1 _13636_/C
+ sky130_fd_sc_hd__and4_1
X_17396_ _21681_/A _17396_/B _17396_/C vssd1 vssd1 vccd1 vccd1 _17397_/A sky130_fd_sc_hd__and3_1
XFILLER_347_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19135_ _23256_/Q _18833_/X _19135_/S vssd1 vssd1 vccd1 vccd1 _19136_/A sky130_fd_sc_hd__mux2_1
X_16347_ _15570_/X _22340_/Q _16355_/S vssd1 vssd1 vccd1 vccd1 _16348_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13559_ _13580_/A _13543_/Y _13188_/A vssd1 vssd1 vccd1 vccd1 _13569_/B sky130_fd_sc_hd__a21oi_4
XFILLER_347_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19066_ _19066_/A vssd1 vssd1 vccd1 vccd1 _23225_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16278_ _18843_/A vssd1 vssd1 vccd1 vccd1 _16278_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_334_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18017_ _18052_/A vssd1 vssd1 vccd1 vccd1 _18017_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_350_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15229_ _22922_/Q _14932_/X _14934_/X _15207_/X vssd1 vssd1 vccd1 vccd1 _15229_/X
+ sky130_fd_sc_hd__o22a_1
Xoutput403 _14022_/X vssd1 vssd1 vccd1 vccd1 din0[7] sky130_fd_sc_hd__buf_2
Xoutput414 _22568_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[15] sky130_fd_sc_hd__buf_2
XFILLER_172_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput425 _22578_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[25] sky130_fd_sc_hd__buf_2
XFILLER_321_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_315_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput436 _22559_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[6] sky130_fd_sc_hd__buf_2
XFILLER_287_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput447 _14521_/A vssd1 vssd1 vccd1 vccd1 probe_isLoad sky130_fd_sc_hd__buf_2
XFILLER_153_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput458 _23883_/Q vssd1 vssd1 vccd1 vccd1 probe_opcode[4] sky130_fd_sc_hd__buf_2
XFILLER_302_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_287_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput469 _23928_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[17] sky130_fd_sc_hd__buf_2
XFILLER_113_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_303_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_302_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19968_ _19968_/A _19971_/C _19971_/D vssd1 vssd1 vccd1 vccd1 _19969_/C sky130_fd_sc_hd__and3_1
XFILLER_234_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_330_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18919_ _18919_/A vssd1 vssd1 vccd1 vccd1 _23160_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_256_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19899_ _19899_/A vssd1 vssd1 vccd1 vccd1 _23581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21930_ _21987_/A vssd1 vssd1 vccd1 vccd1 _22098_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21861_ _21861_/A _22197_/B vssd1 vssd1 vccd1 vccd1 _21861_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23600_ _23600_/CLK _23600_/D vssd1 vssd1 vccd1 vccd1 _23600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20812_ _20626_/B _20810_/X _20811_/X _23758_/Q vssd1 vssd1 vccd1 vccd1 _20813_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21792_ _21792_/A _21792_/B vssd1 vssd1 vccd1 vccd1 _21793_/B sky130_fd_sc_hd__nor2_1
XFILLER_230_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20743_ _23743_/Q _20729_/X _20742_/X _20737_/X vssd1 vssd1 vccd1 vccd1 _23743_/D
+ sky130_fd_sc_hd__o211a_1
X_23531_ _23531_/CLK _23531_/D vssd1 vssd1 vccd1 vccd1 _23531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_357_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_329_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23462_ _23558_/CLK _23462_/D vssd1 vssd1 vccd1 vccd1 _23462_/Q sky130_fd_sc_hd__dfxtp_4
X_20674_ _23732_/Q _20667_/X _20672_/X _20673_/X vssd1 vssd1 vccd1 vccd1 _23732_/D
+ sky130_fd_sc_hd__o211a_1
X_22413_ _23451_/CLK _22413_/D vssd1 vssd1 vccd1 vccd1 _22413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23393_ _23451_/CLK _23393_/D vssd1 vssd1 vccd1 vccd1 _23393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22344_ _23480_/CLK _22344_/D vssd1 vssd1 vccd1 vccd1 _22344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22275_ _23505_/CLK _22275_/D vssd1 vssd1 vccd1 vccd1 _22275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_352_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21226_ _14546_/X _21202_/X _21225_/Y _21218_/X vssd1 vssd1 vccd1 vccd1 _23887_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_340_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21157_ _23867_/Q _21139_/X _21156_/X _21073_/X vssd1 vssd1 vccd1 vccd1 _23867_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_320_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20108_ _23643_/Q _20107_/C _20101_/X vssd1 vssd1 vccd1 vccd1 _20108_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_259_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21088_ _21075_/Y _21301_/D _21087_/Y _20137_/A vssd1 vssd1 vccd1 vccd1 _23845_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_101_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20039_ _20048_/B _20048_/C _23624_/Q vssd1 vssd1 vccd1 vccd1 _20041_/B sky130_fd_sc_hd__a21oi_1
X_12930_ _23321_/Q _23289_/Q _23257_/Q _23545_/Q _12680_/X _12637_/X vssd1 vssd1 vccd1
+ vccd1 _12931_/B sky130_fd_sc_hd__mux4_2
XFILLER_247_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_1_wb_clk_i clkbuf_3_4_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _22477_/Q _22637_/Q _22316_/Q _23452_/Q _12709_/X _12710_/X vssd1 vssd1 vccd1
+ vccd1 _12861_/X sky130_fd_sc_hd__mux4_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _23718_/Q _23848_/Q _15354_/S vssd1 vssd1 vccd1 vccd1 _14600_/X sky130_fd_sc_hd__mux2_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _11821_/A vssd1 vssd1 vccd1 vccd1 _12094_/A sky130_fd_sc_hd__buf_4
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _15580_/A _15580_/B vssd1 vssd1 vccd1 vccd1 _15580_/Y sky130_fd_sc_hd__nor2_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _12843_/A vssd1 vssd1 vccd1 vccd1 _12792_/X sky130_fd_sc_hd__buf_6
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _21300_/B _14192_/B _14530_/X vssd1 vssd1 vccd1 vccd1 _14531_/Y sky130_fd_sc_hd__o21ai_1
X_11743_ _23472_/Q _23568_/Q _22532_/Q _22336_/Q _11741_/X _12009_/A vssd1 vssd1 vccd1
+ vccd1 _11744_/B sky130_fd_sc_hd__mux4_1
XFILLER_159_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23729_ _23861_/CLK _23729_/D vssd1 vssd1 vccd1 vccd1 _23729_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17250_ _17250_/A vssd1 vssd1 vccd1 vccd1 _17292_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_169_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14462_ _14906_/A vssd1 vssd1 vccd1 vccd1 _15593_/A sky130_fd_sc_hd__clkbuf_4
X_11674_ _12909_/A _11674_/B vssd1 vssd1 vccd1 vccd1 _11674_/X sky130_fd_sc_hd__or2_1
XFILLER_175_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_329_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16201_ _14541_/X _14557_/A _14543_/X vssd1 vssd1 vccd1 vccd1 _18770_/B sky130_fd_sc_hd__o21a_1
X_13413_ _14675_/A _20214_/A vssd1 vssd1 vccd1 vccd1 _14288_/A sky130_fd_sc_hd__nor2_1
X_17181_ _17268_/A vssd1 vssd1 vccd1 vccd1 _17181_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14393_ _14393_/A vssd1 vssd1 vccd1 vccd1 _14393_/X sky130_fd_sc_hd__buf_8
XFILLER_329_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16132_ _13410_/B _15256_/B _16131_/Y _13439_/A vssd1 vssd1 vccd1 vccd1 _16132_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_344_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_319_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13344_ _13344_/A _13344_/B vssd1 vssd1 vccd1 vccd1 _13344_/X sky130_fd_sc_hd__or2_1
XFILLER_194_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_304_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16063_ _23681_/Q _16102_/B vssd1 vssd1 vccd1 vccd1 _16063_/X sky130_fd_sc_hd__or2_1
X_13275_ _13275_/A vssd1 vssd1 vccd1 vccd1 _13275_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_170_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_335_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_331_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15014_ _14640_/X _14645_/X _15129_/S vssd1 vssd1 vccd1 vccd1 _15014_/X sky130_fd_sc_hd__mux2_2
XFILLER_297_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12226_ _22461_/Q _22621_/Q _22300_/Q _23436_/Q _12215_/X _12216_/X vssd1 vssd1 vccd1
+ vccd1 _12226_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_331_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_335_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19822_ _23547_/Q _19236_/A _19826_/S vssd1 vssd1 vccd1 vccd1 _19823_/A sky130_fd_sc_hd__mux2_1
XFILLER_311_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12157_ _12137_/Y _20264_/A _12157_/S vssd1 vssd1 vccd1 vccd1 _12163_/A sky130_fd_sc_hd__mux2_2
XFILLER_69_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11108_ _14133_/B vssd1 vssd1 vccd1 vccd1 _14815_/B sky130_fd_sc_hd__buf_4
X_19753_ _19753_/A vssd1 vssd1 vccd1 vccd1 _23516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_284_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16965_ _21300_/B _16961_/X _17318_/S vssd1 vssd1 vccd1 vccd1 _16965_/X sky130_fd_sc_hd__mux2_1
X_12088_ _13421_/A _12157_/S _11400_/A _12087_/X vssd1 vssd1 vccd1 vccd1 _12112_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_351_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15916_ _13573_/A _15196_/X _14761_/A vssd1 vssd1 vccd1 vccd1 _15916_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_49_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18704_ _16822_/X _23079_/Q _18708_/S vssd1 vssd1 vccd1 vccd1 _18705_/A sky130_fd_sc_hd__mux2_1
X_19684_ _19684_/A vssd1 vssd1 vccd1 vccd1 _19693_/S sky130_fd_sc_hd__buf_6
XFILLER_49_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16896_ _16896_/A vssd1 vssd1 vccd1 vccd1 _16909_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_253_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18635_ _18635_/A vssd1 vssd1 vccd1 vccd1 _23048_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _13400_/A _13601_/Y _16031_/S vssd1 vssd1 vccd1 vccd1 _15848_/B sky130_fd_sc_hd__mux2_1
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18566_ _18623_/S vssd1 vssd1 vccd1 vccd1 _18575_/S sky130_fd_sc_hd__buf_6
XFILLER_224_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ _15479_/A _13633_/Y _14529_/A vssd1 vssd1 vccd1 vccd1 _15778_/X sky130_fd_sc_hd__a21o_1
XFILLER_212_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17517_ _17517_/A vssd1 vssd1 vccd1 vccd1 _22665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14729_ _22948_/Q vssd1 vssd1 vccd1 vccd1 _14729_/X sky130_fd_sc_hd__buf_2
XFILLER_342_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18497_ _18494_/X _18496_/Y _18490_/X vssd1 vssd1 vccd1 vccd1 _22993_/D sky130_fd_sc_hd__a21oi_1
XFILLER_178_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17448_ _22635_/Q _16275_/X _17454_/S vssd1 vssd1 vccd1 vccd1 _17449_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17379_ _17379_/A vssd1 vssd1 vccd1 vccd1 _22609_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_308_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_307_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23566_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_119_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19118_ _23248_/Q _18808_/X _19124_/S vssd1 vssd1 vccd1 vccd1 _19119_/A sky130_fd_sc_hd__mux2_1
XFILLER_307_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20390_ _20320_/X _20388_/Y _20389_/X _22197_/A _20294_/X vssd1 vssd1 vccd1 vccd1
+ _20754_/A sky130_fd_sc_hd__a32o_4
XFILLER_229_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_335_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19049_ _16857_/X _23218_/Q _19051_/S vssd1 vssd1 vccd1 vccd1 _19050_/A sky130_fd_sc_hd__mux2_1
XFILLER_334_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_350_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22060_ _23837_/Q _22059_/Y _22242_/B vssd1 vssd1 vccd1 vccd1 _22061_/B sky130_fd_sc_hd__mux2_1
XFILLER_133_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_204_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23500_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_350_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21011_ _20604_/A _21008_/X _21009_/X _21010_/X vssd1 vssd1 vccd1 vccd1 _23819_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput288 _14090_/X vssd1 vssd1 vccd1 vccd1 addr0[3] sky130_fd_sc_hd__buf_2
XFILLER_88_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput299 _13997_/Y vssd1 vssd1 vccd1 vccd1 addr1[5] sky130_fd_sc_hd__buf_2
XFILLER_99_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_303_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_6 _22166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22962_ _23846_/CLK _22962_/D vssd1 vssd1 vccd1 vccd1 _22962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21913_ _21913_/A _21913_/B vssd1 vssd1 vccd1 vccd1 _21913_/X sky130_fd_sc_hd__xor2_1
XFILLER_283_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22893_ _22893_/CLK _22893_/D vssd1 vssd1 vccd1 vccd1 _22893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21844_ _21847_/A _21844_/B vssd1 vssd1 vccd1 vccd1 _21844_/Y sky130_fd_sc_hd__nor2_1
XFILLER_270_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21775_ _21773_/X _21774_/X _21598_/X vssd1 vssd1 vccd1 vccd1 _21775_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_169_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23514_ _23546_/CLK _23514_/D vssd1 vssd1 vccd1 vccd1 _23514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20726_ _13214_/Y _20701_/X _20725_/Y vssd1 vssd1 vccd1 vccd1 _20727_/C sky130_fd_sc_hd__a21oi_2
XFILLER_357_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23445_ _23446_/CLK _23445_/D vssd1 vssd1 vccd1 vccd1 _23445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20657_ _21719_/A _20648_/X _20656_/Y vssd1 vssd1 vccd1 vccd1 _20658_/C sky130_fd_sc_hd__a21oi_1
XFILLER_183_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23376_ _23951_/A _23376_/D vssd1 vssd1 vccd1 vccd1 _23376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11390_ _13185_/S vssd1 vssd1 vccd1 vccd1 _11486_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_286_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20588_ _20588_/A _20966_/A vssd1 vssd1 vccd1 vccd1 _20591_/B sky130_fd_sc_hd__nor2_2
XFILLER_358_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22327_ _23555_/CLK _22327_/D vssd1 vssd1 vccd1 vccd1 _22327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_340_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13060_ _13121_/A _13060_/B vssd1 vssd1 vccd1 vccd1 _13060_/Y sky130_fd_sc_hd__nor2_1
XFILLER_191_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_313_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22258_ _21287_/A _22247_/X _22257_/X _21193_/C vssd1 vssd1 vccd1 vccd1 _22258_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_152_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12011_ _12949_/A _12011_/B vssd1 vssd1 vccd1 vccd1 _12011_/Y sky130_fd_sc_hd__nor2_1
X_21209_ _21215_/A _21209_/B vssd1 vssd1 vccd1 vccd1 _21210_/A sky130_fd_sc_hd__and2_1
X_22189_ _22189_/A _22189_/B vssd1 vssd1 vccd1 vccd1 _22189_/X sky130_fd_sc_hd__xor2_1
XFILLER_79_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16750_ _16759_/A _16750_/B vssd1 vssd1 vccd1 vccd1 _16751_/A sky130_fd_sc_hd__or2_1
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13962_ _13962_/A _13965_/B vssd1 vssd1 vccd1 vccd1 _13962_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15701_ _21888_/A _23928_/Q _15701_/C vssd1 vssd1 vccd1 vccd1 _21868_/B sky130_fd_sc_hd__and3_2
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_79_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23547_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12913_ _12893_/Y _20334_/A _12913_/S vssd1 vssd1 vccd1 vccd1 _13493_/B sky130_fd_sc_hd__mux2_4
X_16681_ _18277_/A vssd1 vssd1 vccd1 vccd1 _19987_/A sky130_fd_sc_hd__buf_12
XFILLER_219_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13893_ _13893_/A vssd1 vssd1 vccd1 vccd1 _13933_/A sky130_fd_sc_hd__buf_2
XFILLER_206_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18420_ _22968_/Q _18420_/B vssd1 vssd1 vccd1 vccd1 _18427_/C sky130_fd_sc_hd__and2_2
XFILLER_250_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15632_ _15673_/A vssd1 vssd1 vccd1 vccd1 _15923_/A sky130_fd_sc_hd__clkbuf_2
X_12844_ _12844_/A vssd1 vssd1 vccd1 vccd1 _12844_/X sky130_fd_sc_hd__buf_4
XFILLER_15_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _22944_/Q _18351_/B vssd1 vssd1 vccd1 vccd1 _18357_/C sky130_fd_sc_hd__and2_1
XFILLER_15_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _15531_/X _15562_/X _16154_/A vssd1 vssd1 vccd1 vccd1 _15564_/B sky130_fd_sc_hd__mux2_1
X_12775_ _12745_/X _12667_/X _11402_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13534_/A
+ sky130_fd_sc_hd__a22o_4
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17245_/A _17301_/X _17262_/X _17283_/X vssd1 vssd1 vccd1 vccd1 _17302_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_199_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _22914_/Q _14509_/X _14513_/X _22946_/Q vssd1 vssd1 vccd1 vccd1 _14514_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_199_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18282_ _22920_/Q _18276_/C _18281_/Y vssd1 vssd1 vccd1 vccd1 _22920_/D sky130_fd_sc_hd__o21a_1
X_11726_ _11718_/Y _11721_/Y _11723_/Y _11725_/Y _11243_/A vssd1 vssd1 vccd1 vccd1
+ _11727_/C sky130_fd_sc_hd__o221a_1
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _15090_/A _15491_/X _15493_/Y vssd1 vssd1 vccd1 vccd1 _15494_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_348_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17233_ _23484_/Q _17230_/X _17231_/X _17181_/X _17232_/Y vssd1 vssd1 vccd1 vccd1
+ _17233_/X sky130_fd_sc_hd__a32o_1
XFILLER_187_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14445_ _15346_/A vssd1 vssd1 vccd1 vccd1 _14755_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11657_ _11657_/A vssd1 vssd1 vccd1 vccd1 _11657_/X sky130_fd_sc_hd__buf_2
XFILLER_30_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_329_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_329_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17164_ _17160_/Y _17169_/A _17163_/X _17078_/A vssd1 vssd1 vccd1 vccd1 _17164_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_196_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_316_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14376_ _14381_/B _14952_/S vssd1 vssd1 vccd1 vccd1 _14376_/X sky130_fd_sc_hd__or2b_1
X_11588_ _12425_/A vssd1 vssd1 vccd1 vccd1 _12350_/A sky130_fd_sc_hd__buf_4
XFILLER_127_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16115_ _16154_/A _16115_/B vssd1 vssd1 vccd1 vccd1 _16115_/Y sky130_fd_sc_hd__nor2_1
X_13327_ _13599_/A _13327_/B vssd1 vssd1 vccd1 vccd1 _15718_/A sky130_fd_sc_hd__xnor2_4
XFILLER_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_346_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17095_ _23471_/Q _17061_/X _17062_/X _17094_/X _15312_/X vssd1 vssd1 vccd1 vccd1
+ _17095_/X sky130_fd_sc_hd__a32o_1
XFILLER_304_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16046_ _23005_/Q _16084_/A _16085_/A input234/X vssd1 vssd1 vccd1 vccd1 _22139_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_346_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13258_ _23233_/Q _23201_/Q _23169_/Q _23137_/Q _11206_/X _11208_/X vssd1 vssd1 vccd1
+ vccd1 _13259_/B sky130_fd_sc_hd__mux4_2
XFILLER_332_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_320_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_331_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12209_ _12475_/A vssd1 vssd1 vccd1 vccd1 _12209_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_142_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13189_ _22801_/Q _22769_/Q _22670_/Q _22737_/Q _13088_/S _11207_/A vssd1 vssd1 vccd1
+ vccd1 _13189_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_297_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19805_ _19805_/A vssd1 vssd1 vccd1 vccd1 _23539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17997_ _22841_/Q _17981_/X _17996_/X _17979_/X vssd1 vssd1 vccd1 vccd1 _22841_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19736_ _19736_/A vssd1 vssd1 vccd1 vccd1 _23508_/D sky130_fd_sc_hd__clkbuf_1
X_16948_ _16940_/X _16932_/A _16947_/X vssd1 vssd1 vccd1 vccd1 _16948_/X sky130_fd_sc_hd__a21o_1
XFILLER_78_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_293_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16879_ _19229_/A vssd1 vssd1 vccd1 vccd1 _16879_/X sky130_fd_sc_hd__clkbuf_2
X_19667_ _19220_/X _23478_/Q _19671_/S vssd1 vssd1 vccd1 vccd1 _19668_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18618_ _18618_/A vssd1 vssd1 vccd1 vccd1 _23041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19598_ _19598_/A vssd1 vssd1 vccd1 vccd1 _23447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_252_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18549_ _18549_/A _18549_/B vssd1 vssd1 vccd1 vccd1 _18550_/D sky130_fd_sc_hd__nor2_1
XFILLER_212_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21560_ _21560_/A vssd1 vssd1 vccd1 vccd1 _21560_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_221_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20511_ _23704_/Q _20517_/B _20511_/C vssd1 vssd1 vccd1 vccd1 _20515_/B sky130_fd_sc_hd__and3_1
XFILLER_166_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21491_ _22061_/A vssd1 vssd1 vccd1 vccd1 _21491_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_355_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23230_ _23550_/CLK _23230_/D vssd1 vssd1 vccd1 vccd1 _23230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_308_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20442_ _23696_/Q _20448_/B vssd1 vssd1 vccd1 vccd1 _20442_/X sky130_fd_sc_hd__or2_1
XFILLER_193_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23161_ _23545_/CLK _23161_/D vssd1 vssd1 vccd1 vccd1 _23161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20373_ _23679_/Q _20177_/A _20372_/Y _20360_/X vssd1 vssd1 vccd1 vccd1 _23679_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_335_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_323_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22112_ _21838_/A _22110_/Y _22111_/Y _21361_/A vssd1 vssd1 vccd1 vccd1 _22112_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_350_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23092_ _23510_/CLK _23092_/D vssd1 vssd1 vccd1 vccd1 _23092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_350_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_288_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22043_ _21812_/B _22039_/Y _22040_/Y _22042_/Y vssd1 vssd1 vccd1 vccd1 _22053_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_322_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_310_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_331_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_291_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_291_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22945_ _22947_/CLK _22945_/D vssd1 vssd1 vccd1 vccd1 _22945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22876_ _23009_/CLK _22876_/D vssd1 vssd1 vccd1 vccd1 _22876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21827_ _21827_/A _21826_/Y vssd1 vssd1 vccd1 vccd1 _21828_/B sky130_fd_sc_hd__or2b_1
XPHY_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12560_ _22361_/Q _22393_/Q _22682_/Q _23049_/Q _12244_/A _12292_/A vssd1 vssd1 vccd1
+ vccd1 _12561_/B sky130_fd_sc_hd__mux4_1
XPHY_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21758_ _21758_/A _21758_/B vssd1 vssd1 vccd1 vccd1 _21758_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_54_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11511_ _13273_/A _11511_/B vssd1 vssd1 vccd1 vccd1 _11511_/Y sky130_fd_sc_hd__nand2_1
XFILLER_358_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_197_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23560_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20709_ _14393_/X _20692_/X _20702_/X vssd1 vssd1 vccd1 vccd1 _20709_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_297_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12491_ _12321_/A _12490_/X _11678_/A vssd1 vssd1 vccd1 vccd1 _12491_/X sky130_fd_sc_hd__o21a_1
XFILLER_339_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21689_ _21689_/A _21689_/B _21689_/C _21694_/B vssd1 vssd1 vccd1 vccd1 _21690_/C
+ sky130_fd_sc_hd__nor4_1
XFILLER_11_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14230_ _14724_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _15189_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_126_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _23649_/CLK sky130_fd_sc_hd__clkbuf_16
X_11442_ _13107_/A vssd1 vssd1 vccd1 vccd1 _11502_/A sky130_fd_sc_hd__buf_4
X_23428_ _23556_/CLK _23428_/D vssd1 vssd1 vccd1 vccd1 _23428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14161_ _14161_/A vssd1 vssd1 vccd1 vccd1 _14164_/A sky130_fd_sc_hd__clkbuf_2
X_11373_ _13278_/A _11370_/X _11372_/X _11353_/A vssd1 vssd1 vccd1 vccd1 _11373_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23359_ _23423_/CLK _23359_/D vssd1 vssd1 vccd1 vccd1 _23359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_314_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_353_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_313_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13112_ _23937_/Q vssd1 vssd1 vccd1 vccd1 _16003_/A sky130_fd_sc_hd__inv_2
XFILLER_314_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14092_ _22593_/Q _14081_/X _14091_/Y _14083_/X vssd1 vssd1 vccd1 vccd1 _14092_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_166_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_341_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17920_ _22819_/Q _17914_/X _17919_/X _17912_/X vssd1 vssd1 vccd1 vccd1 _22819_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_313_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13043_ _13051_/A _13042_/X _12816_/X vssd1 vssd1 vccd1 vccd1 _13043_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17851_ _22797_/Q _17610_/X _17859_/S vssd1 vssd1 vccd1 vccd1 _17852_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16802_ _16802_/A vssd1 vssd1 vccd1 vccd1 _22517_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_310_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17782_ _17782_/A vssd1 vssd1 vccd1 vccd1 _22766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14994_ _23786_/Q _14917_/X _14919_/X vssd1 vssd1 vccd1 vccd1 _14994_/X sky130_fd_sc_hd__a21o_1
XFILLER_120_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19521_ _19217_/X _23413_/Q _19527_/S vssd1 vssd1 vccd1 vccd1 _19522_/A sky130_fd_sc_hd__mux2_1
XFILLER_282_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16733_ _16733_/A vssd1 vssd1 vccd1 vccd1 _22497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_281_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13945_ _13951_/A _13945_/B vssd1 vssd1 vccd1 vccd1 _13945_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19452_ _19452_/A vssd1 vssd1 vccd1 vccd1 _23382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16664_ _16664_/A vssd1 vssd1 vccd1 vccd1 _16673_/S sky130_fd_sc_hd__buf_6
XFILLER_207_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13876_ _11249_/Y _13798_/B _13709_/A vssd1 vssd1 vccd1 vccd1 _13876_/X sky130_fd_sc_hd__a21o_1
XFILLER_250_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18403_ _18403_/A _18409_/C vssd1 vssd1 vccd1 vccd1 _18403_/Y sky130_fd_sc_hd__nor2_1
X_15615_ _14987_/B _13612_/X _15574_/X _15614_/Y vssd1 vssd1 vccd1 vccd1 _15615_/X
+ sky130_fd_sc_hd__o211a_2
X_19383_ _23352_/Q _18833_/X _19383_/S vssd1 vssd1 vccd1 vccd1 _19384_/A sky130_fd_sc_hd__mux2_1
X_12827_ _12836_/A _12826_/X _12687_/X vssd1 vssd1 vccd1 vccd1 _12827_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_201_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16595_ _16013_/X _22448_/Q _16601_/S vssd1 vssd1 vccd1 vccd1 _16596_/A sky130_fd_sc_hd__mux2_1
XFILLER_250_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18334_ _22938_/Q _18334_/B vssd1 vssd1 vccd1 vccd1 _18341_/C sky130_fd_sc_hd__and2_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15546_ _14837_/X _15537_/X _15545_/X vssd1 vssd1 vccd1 vccd1 _15546_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_348_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12758_ _12871_/A _12758_/B vssd1 vssd1 vccd1 vccd1 _12758_/Y sky130_fd_sc_hd__nor2_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18265_ _19987_/A vssd1 vssd1 vccd1 vccd1 _18268_/A sky130_fd_sc_hd__clkbuf_16
X_11709_ _22304_/Q _23440_/Q _11894_/S vssd1 vssd1 vccd1 vccd1 _11709_/X sky130_fd_sc_hd__mux2_1
X_15477_ _22992_/Q _15620_/A _15621_/A input220/X vssd1 vssd1 vccd1 vccd1 _21766_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_187_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12689_ _11233_/A _12670_/Y _12678_/Y _12682_/Y _12688_/Y vssd1 vssd1 vccd1 vccd1
+ _12689_/X sky130_fd_sc_hd__o32a_1
XFILLER_336_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17216_ _17169_/X _17214_/X _17195_/X _17215_/X vssd1 vssd1 vccd1 vccd1 _17216_/X
+ sky130_fd_sc_hd__a211o_1
X_14428_ _14510_/A _15148_/A vssd1 vssd1 vccd1 vccd1 _15558_/A sky130_fd_sc_hd__and2b_1
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18196_ _18194_/X _18195_/Y _18191_/D vssd1 vssd1 vccd1 vccd1 _18196_/X sky130_fd_sc_hd__a21o_1
XFILLER_163_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17147_ _23476_/Q _17170_/B vssd1 vssd1 vccd1 vccd1 _17147_/Y sky130_fd_sc_hd__nand2_1
XFILLER_190_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14359_ _14358_/A _13306_/B _14358_/Y vssd1 vssd1 vccd1 vccd1 _14359_/X sky130_fd_sc_hd__o21a_1
XFILLER_345_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_317_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_332_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_305_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17078_ _17078_/A vssd1 vssd1 vccd1 vccd1 _17078_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16029_ _22941_/Q _15259_/B _16019_/X _16028_/Y _14727_/X vssd1 vssd1 vccd1 vccd1
+ _16029_/X sky130_fd_sc_hd__a221o_1
XFILLER_171_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_300_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_300_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19719_ _19191_/X _23501_/Q _19721_/S vssd1 vssd1 vccd1 vccd1 _19720_/A sky130_fd_sc_hd__mux2_1
X_20991_ _23813_/Q _21064_/B vssd1 vssd1 vccd1 vccd1 _20991_/X sky130_fd_sc_hd__or2_1
XFILLER_93_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22730_ _23574_/CLK _22730_/D vssd1 vssd1 vccd1 vccd1 _22730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22661_ _23444_/CLK _22661_/D vssd1 vssd1 vccd1 vccd1 _22661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21612_ _21984_/A vssd1 vssd1 vccd1 vccd1 _21612_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22592_ _22977_/CLK _22592_/D vssd1 vssd1 vccd1 vccd1 _22592_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_222_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21543_ _21451_/B _21543_/B _21543_/C vssd1 vssd1 vccd1 vccd1 _21543_/X sky130_fd_sc_hd__and3b_1
XFILLER_139_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_355_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21474_ _21474_/A _21712_/S vssd1 vssd1 vccd1 vccd1 _21474_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_354_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20425_ _20585_/A _20408_/X _20424_/X _20420_/X vssd1 vssd1 vccd1 vccd1 _23689_/D
+ sky130_fd_sc_hd__o211a_1
X_23213_ _23407_/CLK _23213_/D vssd1 vssd1 vccd1 vccd1 _23213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23144_ _23144_/CLK _23144_/D vssd1 vssd1 vccd1 vccd1 _23144_/Q sky130_fd_sc_hd__dfxtp_1
X_20356_ _20302_/X _20354_/X _20355_/Y _22067_/A _20307_/X vssd1 vssd1 vccd1 vccd1
+ _20723_/A sky130_fd_sc_hd__a32o_4
XFILLER_84_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_350_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_351_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23075_ _23491_/CLK _23075_/D vssd1 vssd1 vccd1 vccd1 _23075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20287_ _21773_/A _20368_/B vssd1 vssd1 vccd1 vccd1 _20289_/B sky130_fd_sc_hd__or2_1
XTAP_6226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22026_ _23836_/Q _22190_/B _22025_/Y _21377_/A vssd1 vssd1 vccd1 vccd1 _22026_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11991_ _11631_/X _11984_/X _11986_/X _11990_/X _11657_/X vssd1 vssd1 vccd1 vccd1
+ _12002_/B sky130_fd_sc_hd__a311o_1
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13730_ _15830_/A vssd1 vssd1 vccd1 vccd1 _13730_/X sky130_fd_sc_hd__buf_2
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22928_ _22961_/CLK _22928_/D vssd1 vssd1 vccd1 vccd1 _22928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13661_ _22601_/Q _22602_/Q _22599_/Q _22600_/Q vssd1 vssd1 vccd1 vccd1 _13662_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_216_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22859_ _22908_/CLK _22859_/D vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15400_ _23793_/Q _14603_/A _14918_/A vssd1 vssd1 vccd1 vccd1 _15400_/X sky130_fd_sc_hd__a21o_1
XFILLER_232_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _13942_/A _15198_/A vssd1 vssd1 vccd1 vccd1 _13371_/A sky130_fd_sc_hd__nor2_4
X_16380_ _16380_/A vssd1 vssd1 vccd1 vccd1 _22355_/D sky130_fd_sc_hd__clkbuf_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _13592_/A _13592_/B vssd1 vssd1 vccd1 vccd1 _13592_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_12_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15331_ _15331_/A _15433_/B vssd1 vssd1 vccd1 vccd1 _15331_/Y sky130_fd_sc_hd__nand2_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12543_ _11241_/A _12530_/X _12542_/X _12468_/B vssd1 vssd1 vccd1 vccd1 _13695_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_346_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_345_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18050_ _22855_/Q _18035_/X _18049_/X _18045_/X vssd1 vssd1 vccd1 vccd1 _22855_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15262_ _23662_/Q _15353_/B vssd1 vssd1 vccd1 vccd1 _15262_/X sky130_fd_sc_hd__or2_1
XFILLER_346_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12474_ _12485_/A _12474_/B vssd1 vssd1 vccd1 vccd1 _12474_/X sky130_fd_sc_hd__or2_1
XFILLER_185_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17001_ input70/X input65/X _17029_/S vssd1 vssd1 vccd1 vccd1 _17001_/X sky130_fd_sc_hd__mux2_8
XFILLER_184_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14213_ _14820_/A _14821_/B vssd1 vssd1 vccd1 vccd1 _14569_/A sky130_fd_sc_hd__or2_1
X_11425_ _23427_/Q _23043_/Q _23395_/Q _23363_/Q _11157_/X _11418_/X vssd1 vssd1 vccd1
+ vccd1 _11425_/X sky130_fd_sc_hd__mux4_2
XFILLER_144_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15193_ _15538_/A _14312_/X _14671_/S vssd1 vssd1 vccd1 vccd1 _15193_/X sky130_fd_sc_hd__o21a_1
XFILLER_354_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_327_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_314_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14144_ _15416_/A _17648_/A vssd1 vssd1 vccd1 vccd1 _16937_/A sky130_fd_sc_hd__or2_1
XFILLER_153_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11356_ _12476_/A vssd1 vssd1 vccd1 vccd1 _12329_/A sky130_fd_sc_hd__buf_4
XFILLER_180_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_342_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14075_ _22810_/Q _14013_/X _14074_/X vssd1 vssd1 vccd1 vccd1 _14075_/X sky130_fd_sc_hd__a21bo_4
X_18952_ _18952_/A vssd1 vssd1 vccd1 vccd1 _23174_/D sky130_fd_sc_hd__clkbuf_1
X_11287_ _12745_/A vssd1 vssd1 vccd1 vccd1 _11288_/A sky130_fd_sc_hd__buf_4
XFILLER_258_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_298_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17903_ _17959_/A vssd1 vssd1 vccd1 vccd1 _17903_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_94_wb_clk_i _22899_/CLK vssd1 vssd1 vccd1 vccd1 _23586_/CLK sky130_fd_sc_hd__clkbuf_16
X_13026_ _13026_/A _13026_/B vssd1 vssd1 vccd1 vccd1 _13026_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18883_ _23144_/Q _18782_/X _18885_/S vssd1 vssd1 vccd1 vccd1 _18884_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_23_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23902_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17834_ _17834_/A vssd1 vssd1 vccd1 vccd1 _22789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17765_ _22759_/Q _17591_/X _17765_/S vssd1 vssd1 vccd1 vccd1 _17766_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14977_ _15049_/C _14977_/B vssd1 vssd1 vccd1 vccd1 _21421_/B sky130_fd_sc_hd__or2_1
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19504_ _19504_/A vssd1 vssd1 vccd1 vccd1 _23405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16716_ _22493_/Q _16711_/X _16712_/X input38/X vssd1 vssd1 vccd1 vccd1 _16717_/B
+ sky130_fd_sc_hd__o22a_1
X_13928_ _13928_/A _13928_/B vssd1 vssd1 vccd1 vccd1 _15123_/A sky130_fd_sc_hd__xnor2_4
X_17696_ _22728_/Q _17594_/X _17704_/S vssd1 vssd1 vccd1 vccd1 _17697_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_400 _14098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_411 _14030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_422 _14067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16647_ _22471_/Q _16262_/X _16651_/S vssd1 vssd1 vccd1 vccd1 _16648_/A sky130_fd_sc_hd__mux2_1
X_19435_ _19481_/S vssd1 vssd1 vccd1 vccd1 _19444_/S sky130_fd_sc_hd__buf_4
X_13859_ _13273_/B _13808_/X _13709_/A vssd1 vssd1 vccd1 vccd1 _13859_/X sky130_fd_sc_hd__a21o_1
XINSDIODE2_433 _23881_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_288_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_444 _23918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_455 _23924_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_466 _22146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16578_ _16578_/A vssd1 vssd1 vccd1 vccd1 _22440_/D sky130_fd_sc_hd__clkbuf_1
X_19366_ _23344_/Q _18808_/X _19372_/S vssd1 vssd1 vccd1 vccd1 _19367_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_477 _21340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_488 _13963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_499 _14831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18317_ _18317_/A _18323_/C vssd1 vssd1 vccd1 vccd1 _18317_/Y sky130_fd_sc_hd__nor2_1
X_15529_ _21791_/A _23925_/Q _15529_/C vssd1 vssd1 vccd1 vccd1 _15611_/B sky130_fd_sc_hd__and3_1
X_19297_ _19297_/A vssd1 vssd1 vccd1 vccd1 _23313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_349_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_337_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18248_ _22862_/Q _18242_/X _18247_/X _18245_/X vssd1 vssd1 vccd1 vccd1 _22910_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_351_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18179_ _18179_/A _18195_/B vssd1 vssd1 vccd1 vccd1 _18179_/Y sky130_fd_sc_hd__nand2_1
XFILLER_190_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20210_ _20196_/X _20208_/X _20209_/Y _21474_/A _20200_/X vssd1 vssd1 vccd1 vccd1
+ _20595_/A sky130_fd_sc_hd__a32o_4
XFILLER_317_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_305_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21190_ _23944_/Q _23943_/Q vssd1 vssd1 vccd1 vccd1 _21191_/B sky130_fd_sc_hd__nor2_1
XFILLER_289_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_289_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20141_ _21285_/A _20186_/B _20139_/Y _20140_/X vssd1 vssd1 vccd1 vccd1 _20986_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_132_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_253_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20072_ _21122_/A _20072_/B vssd1 vssd1 vccd1 vccd1 _20072_/Y sky130_fd_sc_hd__nor2_1
XFILLER_298_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23900_ _23902_/CLK _23900_/D vssd1 vssd1 vccd1 vccd1 _23900_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23831_ _23832_/CLK _23831_/D vssd1 vssd1 vccd1 vccd1 _23831_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_245_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23762_ _23878_/CLK _23762_/D vssd1 vssd1 vccd1 vccd1 _23762_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_226_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20974_ _23807_/Q _20969_/X _20973_/X _20964_/X vssd1 vssd1 vccd1 vccd1 _23807_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22713_ _23896_/CLK _22713_/D vssd1 vssd1 vccd1 vccd1 _22713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23693_ _23693_/CLK _23693_/D vssd1 vssd1 vccd1 vccd1 _23693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22644_ _23893_/CLK _22644_/D vssd1 vssd1 vccd1 vccd1 _22644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_322_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_356_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_322_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22575_ _23646_/CLK _22575_/D vssd1 vssd1 vccd1 vccd1 _22575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_327_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21526_ _21526_/A _21549_/A _21526_/C vssd1 vssd1 vccd1 vccd1 _21546_/A sky130_fd_sc_hd__and3_1
XFILLER_139_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_342_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21457_ _22019_/A vssd1 vssd1 vccd1 vccd1 _21838_/A sky130_fd_sc_hd__buf_2
XFILLER_119_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_294_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11210_ _13253_/A _11209_/X _11135_/A vssd1 vssd1 vccd1 vccd1 _11210_/Y sky130_fd_sc_hd__o21ai_1
X_20408_ _20428_/A vssd1 vssd1 vccd1 vccd1 _20408_/X sky130_fd_sc_hd__clkbuf_2
X_12190_ _12421_/A vssd1 vssd1 vccd1 vccd1 _12565_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_324_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21388_ _15864_/X _15631_/A _21336_/X _14538_/X vssd1 vssd1 vccd1 vccd1 _21425_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_311_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23127_ _23543_/CLK _23127_/D vssd1 vssd1 vccd1 vccd1 _23127_/Q sky130_fd_sc_hd__dfxtp_1
X_11141_ _11141_/A vssd1 vssd1 vccd1 vccd1 _12985_/A sky130_fd_sc_hd__buf_2
XTAP_6001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20339_ _20333_/X _20708_/A _20338_/X _20324_/X vssd1 vssd1 vccd1 vccd1 _23674_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_6012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11072_ _12345_/B vssd1 vssd1 vccd1 vccd1 _14172_/C sky130_fd_sc_hd__buf_2
XFILLER_295_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23058_ _23058_/CLK _23058_/D vssd1 vssd1 vccd1 vccd1 _23058_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput100 dout0[61] vssd1 vssd1 vccd1 vccd1 input100/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput111 dout1[13] vssd1 vssd1 vccd1 vccd1 input111/X sky130_fd_sc_hd__clkbuf_1
XTAP_5322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput122 dout1[23] vssd1 vssd1 vccd1 vccd1 input122/X sky130_fd_sc_hd__clkbuf_1
X_14900_ _22918_/Q _14988_/B vssd1 vssd1 vccd1 vccd1 _14900_/X sky130_fd_sc_hd__and2_1
XTAP_5333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_292_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22009_ _22161_/A vssd1 vssd1 vccd1 vccd1 _22205_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput133 dout1[33] vssd1 vssd1 vccd1 vccd1 input133/X sky130_fd_sc_hd__buf_2
XTAP_6089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _23804_/Q _15219_/X _14919_/X vssd1 vssd1 vccd1 vccd1 _15880_/X sky130_fd_sc_hd__a21o_1
Xinput144 dout1[43] vssd1 vssd1 vccd1 vccd1 input144/X sky130_fd_sc_hd__buf_2
XTAP_5355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput155 dout1[53] vssd1 vssd1 vccd1 vccd1 input155/X sky130_fd_sc_hd__buf_2
XTAP_5366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput166 dout1[63] vssd1 vssd1 vccd1 vccd1 input166/X sky130_fd_sc_hd__buf_2
XTAP_5377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14831_ input135/X input140/X _15052_/S vssd1 vssd1 vccd1 vccd1 _14831_/X sky130_fd_sc_hd__mux2_8
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput177 irq[15] vssd1 vssd1 vccd1 vccd1 _20513_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput188 jtag_tdi vssd1 vssd1 vccd1 vccd1 _18009_/B sky130_fd_sc_hd__buf_12
Xinput199 localMemory_wb_adr_i[18] vssd1 vssd1 vccd1 vccd1 input199/X sky130_fd_sc_hd__clkbuf_1
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_291_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _18776_/A vssd1 vssd1 vccd1 vccd1 _17550_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14762_ _14762_/A vssd1 vssd1 vccd1 vccd1 _15801_/A sky130_fd_sc_hd__clkbuf_2
X_11974_ _22276_/Q _23092_/Q _23508_/Q _22437_/Q _11972_/X _11973_/X vssd1 vssd1 vccd1
+ vccd1 _11975_/B sky130_fd_sc_hd__mux4_1
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16501_ _16501_/A vssd1 vssd1 vccd1 vccd1 _22407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _13713_/A vssd1 vssd1 vccd1 vccd1 _13713_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17481_ _22649_/Q _16217_/X _17483_/S vssd1 vssd1 vccd1 vccd1 _17482_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14693_ _14587_/X _14619_/X _14692_/X vssd1 vssd1 vccd1 vccd1 _14693_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_189_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19220_ _19220_/A vssd1 vssd1 vccd1 vccd1 _19220_/X sky130_fd_sc_hd__clkbuf_2
X_16432_ _15785_/X _22377_/Q _16440_/S vssd1 vssd1 vccd1 vccd1 _16433_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_141_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _23856_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_177_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13644_ _13942_/B _13526_/X _13524_/Y vssd1 vssd1 vccd1 vccd1 _13948_/B sky130_fd_sc_hd__o21a_2
XFILLER_60_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19151_ _23263_/Q _18856_/X _19157_/S vssd1 vssd1 vccd1 vccd1 _19152_/A sky130_fd_sc_hd__mux2_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _16363_/A vssd1 vssd1 vccd1 vccd1 _22347_/D sky130_fd_sc_hd__clkbuf_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13581_/A _13575_/B vssd1 vssd1 vccd1 vccd1 _13575_/Y sky130_fd_sc_hd__nand2_1
XFILLER_346_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18102_ _22871_/Q _18097_/X _18098_/X _23004_/Q _18099_/X vssd1 vssd1 vccd1 vccd1
+ _18102_/X sky130_fd_sc_hd__a221o_1
XFILLER_318_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _14215_/X _21231_/A _15313_/X _14882_/X vssd1 vssd1 vccd1 vccd1 _15314_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_19082_ _16905_/X _23233_/Q _19084_/S vssd1 vssd1 vccd1 vccd1 _19083_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12526_ _23397_/Q _23013_/Q _23365_/Q _23333_/Q _11146_/A _11701_/A vssd1 vssd1 vccd1
+ vccd1 _12526_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_307_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16294_ _18859_/A vssd1 vssd1 vccd1 vccd1 _16294_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18033_ _22849_/Q _18017_/X _18020_/X _22982_/Q _18023_/X vssd1 vssd1 vccd1 vccd1
+ _18033_/X sky130_fd_sc_hd__a221o_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_318_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15245_ _13834_/A _15243_/Y _15244_/Y _13739_/A vssd1 vssd1 vccd1 vccd1 _15245_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_157_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12457_ _22294_/Q _23430_/Q _12457_/S vssd1 vssd1 vccd1 vccd1 _12458_/B sky130_fd_sc_hd__mux2_1
XFILLER_8_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11408_ _12891_/A vssd1 vssd1 vccd1 vccd1 _13212_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_299_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15176_ _15176_/A _15176_/B _15176_/C _15116_/Y vssd1 vssd1 vccd1 vccd1 _15176_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_153_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12388_ _22457_/Q _22617_/Q _22296_/Q _23432_/Q _11646_/A _11651_/A vssd1 vssd1 vccd1
+ vccd1 _12388_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_315_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14127_ _18126_/S _22882_/Q _14107_/X _14126_/X vssd1 vssd1 vccd1 vccd1 _14127_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_181_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11339_ _23236_/Q _23204_/Q _23172_/Q _23140_/Q _11468_/A _11469_/A vssd1 vssd1 vccd1
+ vccd1 _11340_/B sky130_fd_sc_hd__mux4_1
XFILLER_4_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19984_ _23606_/Q _23605_/Q vssd1 vssd1 vccd1 vccd1 _19985_/D sky130_fd_sc_hd__and2_1
XFILLER_287_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_330_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18935_ _18935_/A vssd1 vssd1 vccd1 vccd1 _23167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_286_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14058_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14058_/X sky130_fd_sc_hd__buf_2
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13009_ _13002_/X _13004_/X _13006_/X _13008_/X _11276_/A vssd1 vssd1 vccd1 vccd1
+ _13010_/C sky130_fd_sc_hd__a221o_1
X_18866_ _23138_/Q _18865_/X _18866_/S vssd1 vssd1 vccd1 vccd1 _18867_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17817_ _17874_/S vssd1 vssd1 vccd1 vccd1 _17826_/S sky130_fd_sc_hd__buf_6
X_18797_ _18797_/A vssd1 vssd1 vccd1 vccd1 _23116_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17748_ _22751_/Q _17566_/X _17754_/S vssd1 vssd1 vccd1 vccd1 _17749_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_230 _15114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17679_ _17679_/A vssd1 vssd1 vccd1 vccd1 _22720_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_241 _15312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19418_ _23367_/Q _18779_/X _19422_/S vssd1 vssd1 vccd1 vccd1 _19419_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_252 _15510_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_357_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20690_ _23735_/Q _20667_/X _20689_/X _20673_/X vssd1 vssd1 vccd1 vccd1 _23735_/D
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_263 _15651_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_274 _17182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_285 _15959_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_296 _15990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19349_ _19349_/A vssd1 vssd1 vccd1 vccd1 _23336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_349_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_309_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22360_ _23528_/CLK _22360_/D vssd1 vssd1 vccd1 vccd1 _22360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21311_ _20544_/A _21308_/C _22711_/Q vssd1 vssd1 vccd1 vccd1 _21613_/A sky130_fd_sc_hd__o21a_4
XFILLER_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22291_ _23491_/CLK _22291_/D vssd1 vssd1 vccd1 vccd1 _22291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_324_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21242_ _21242_/A vssd1 vssd1 vccd1 vccd1 _21242_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21173_ _21173_/A _21177_/B vssd1 vssd1 vccd1 vccd1 _21173_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_320_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20124_ _20137_/A _20124_/B _20131_/D vssd1 vssd1 vccd1 vccd1 _23647_/D sky130_fd_sc_hd__nor3_1
XFILLER_264_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20055_ _20066_/B _20063_/C _20066_/A vssd1 vssd1 vccd1 vccd1 _20057_/B sky130_fd_sc_hd__a21oi_1
XFILLER_58_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_292_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23814_ _23818_/CLK _23814_/D vssd1 vssd1 vccd1 vccd1 _23814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23745_ _23915_/CLK _23745_/D vssd1 vssd1 vccd1 vccd1 _23745_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ _21975_/A _20950_/X _20711_/B _20954_/X vssd1 vssd1 vccd1 vccd1 _20957_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_289_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11690_ _13536_/B vssd1 vssd1 vccd1 vccd1 _11691_/B sky130_fd_sc_hd__clkinv_2
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23676_ _23684_/CLK _23676_/D vssd1 vssd1 vccd1 vccd1 _23676_/Q sky130_fd_sc_hd__dfxtp_1
X_20888_ _21148_/A _20888_/B _20888_/C vssd1 vssd1 vccd1 vccd1 _20888_/X sky130_fd_sc_hd__or3_1
XFILLER_347_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22627_ _23567_/CLK _22627_/D vssd1 vssd1 vccd1 vccd1 _22627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_329_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13360_ _13360_/A vssd1 vssd1 vccd1 vccd1 _13464_/B sky130_fd_sc_hd__buf_4
XFILLER_328_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22558_ _22977_/CLK _22558_/D vssd1 vssd1 vccd1 vccd1 _22558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_318_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12311_ _12468_/B _12311_/B _12311_/C vssd1 vssd1 vccd1 vccd1 _13764_/A sky130_fd_sc_hd__or3_4
XFILLER_344_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21509_ _21522_/A _21515_/A vssd1 vssd1 vccd1 vccd1 _21509_/Y sky130_fd_sc_hd__nor2_1
X_13291_ _13291_/A _13291_/B vssd1 vssd1 vccd1 vccd1 _13291_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22489_ _23841_/CLK _22489_/D vssd1 vssd1 vccd1 vccd1 _22489_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15030_ input146/X input111/X _15030_/S vssd1 vssd1 vccd1 vccd1 _15030_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12242_ _22460_/Q _22620_/Q _12242_/S vssd1 vssd1 vccd1 vccd1 _12243_/B sky130_fd_sc_hd__mux2_1
XFILLER_257_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_312_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12173_ _22364_/Q _22396_/Q _22685_/Q _23052_/Q _11148_/A _11840_/X vssd1 vssd1 vccd1
+ vccd1 _12174_/B sky130_fd_sc_hd__mux4_2
XFILLER_269_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_351_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_323_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11124_ _11124_/A vssd1 vssd1 vccd1 vccd1 _13210_/A sky130_fd_sc_hd__buf_6
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16981_ _16981_/A vssd1 vssd1 vccd1 vccd1 _17250_/A sky130_fd_sc_hd__buf_2
XFILLER_96_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18720_ _18720_/A vssd1 vssd1 vccd1 vccd1 _23086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15932_ _15932_/A vssd1 vssd1 vccd1 vccd1 _16085_/A sky130_fd_sc_hd__buf_2
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15863_ _15863_/A vssd1 vssd1 vccd1 vccd1 _22283_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18651_ _18651_/A vssd1 vssd1 vccd1 vccd1 _23055_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17602_ _22695_/Q _17601_/X _17608_/S vssd1 vssd1 vccd1 vccd1 _17603_/A sky130_fd_sc_hd__mux2_1
XFILLER_292_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14814_ _23882_/Q _23881_/Q _14814_/C _21335_/B vssd1 vssd1 vccd1 vccd1 _21382_/A
+ sky130_fd_sc_hd__and4_1
X_18582_ _16854_/X _23025_/Q _18586_/S vssd1 vssd1 vccd1 vccd1 _18583_/A sky130_fd_sc_hd__mux2_1
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15794_ _15633_/X _15433_/Y _15674_/A vssd1 vssd1 vccd1 vccd1 _15794_/X sky130_fd_sc_hd__a21bo_2
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _17533_/A vssd1 vssd1 vccd1 vccd1 _22672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14745_ _14745_/A _21084_/A vssd1 vssd1 vccd1 vccd1 _14745_/Y sky130_fd_sc_hd__nor2_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11957_ _11957_/A vssd1 vssd1 vccd1 vccd1 _12047_/A sky130_fd_sc_hd__buf_2
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17464_ _17464_/A vssd1 vssd1 vccd1 vccd1 _22642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_339_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14676_ _14676_/A _14676_/B vssd1 vssd1 vccd1 vccd1 _14676_/Y sky130_fd_sc_hd__nor2_1
XFILLER_232_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11888_ _13522_/A _13525_/B vssd1 vssd1 vccd1 vccd1 _13518_/A sky130_fd_sc_hd__xnor2_2
XFILLER_349_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16415_ _16415_/A vssd1 vssd1 vccd1 vccd1 _22369_/D sky130_fd_sc_hd__clkbuf_1
X_19203_ _19203_/A vssd1 vssd1 vccd1 vccd1 _23280_/D sky130_fd_sc_hd__clkbuf_1
X_13627_ _21738_/A _13588_/A _15453_/A _13594_/A _13956_/A vssd1 vssd1 vccd1 vccd1
+ _13628_/D sky130_fd_sc_hd__a221oi_1
X_17395_ _17326_/A _17326_/B _17394_/Y _17325_/B vssd1 vssd1 vccd1 vccd1 _17396_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_319_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19134_ _19134_/A vssd1 vssd1 vccd1 vccd1 _23255_/D sky130_fd_sc_hd__clkbuf_1
X_16346_ _16368_/A vssd1 vssd1 vccd1 vccd1 _16355_/S sky130_fd_sc_hd__buf_6
XFILLER_201_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13558_ _13492_/X _13540_/A _13632_/B _13540_/X _13579_/A vssd1 vssd1 vccd1 vccd1
+ _13580_/A sky130_fd_sc_hd__o221ai_4
XFILLER_185_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_347_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19065_ _16879_/X _23225_/Q _19073_/S vssd1 vssd1 vccd1 vccd1 _19066_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12509_ _12500_/X _12504_/X _12506_/X _12508_/X _23898_/Q vssd1 vssd1 vccd1 vccd1
+ _12519_/B sky130_fd_sc_hd__a221o_1
XFILLER_335_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16277_ _16277_/A vssd1 vssd1 vccd1 vccd1 _22314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13489_ _14206_/A _13655_/A vssd1 vssd1 vccd1 vccd1 _13490_/A sky130_fd_sc_hd__nand2_2
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18016_ _18051_/A vssd1 vssd1 vccd1 vccd1 _18016_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15228_ _15207_/X _15225_/X _16028_/A vssd1 vssd1 vccd1 vccd1 _15228_/X sky130_fd_sc_hd__mux2_1
XFILLER_334_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_350_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput404 _14024_/X vssd1 vssd1 vccd1 vccd1 din0[8] sky130_fd_sc_hd__buf_2
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput415 _22569_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[16] sky130_fd_sc_hd__buf_2
XFILLER_126_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput426 _22579_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[26] sky130_fd_sc_hd__buf_2
XFILLER_172_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput437 _22560_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[7] sky130_fd_sc_hd__buf_2
Xoutput448 _13779_/A vssd1 vssd1 vccd1 vccd1 probe_isStore sky130_fd_sc_hd__buf_2
X_15159_ _21522_/A _15159_/B vssd1 vssd1 vccd1 vccd1 _15160_/B sky130_fd_sc_hd__nor2_1
XFILLER_314_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_303_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput459 _23884_/Q vssd1 vssd1 vccd1 vccd1 probe_opcode[5] sky130_fd_sc_hd__buf_2
XFILLER_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_302_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19967_ _23600_/Q _23599_/Q _23598_/Q _23597_/Q vssd1 vssd1 vccd1 vccd1 _19971_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_80_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_312_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18918_ _23160_/Q _18833_/X _18918_/S vssd1 vssd1 vccd1 vccd1 _18919_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19898_ _16284_/X _23581_/Q _19898_/S vssd1 vssd1 vccd1 vccd1 _19899_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18849_ _18849_/A vssd1 vssd1 vccd1 vccd1 _18849_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21860_ _21856_/Y _21857_/X _21858_/Y _21676_/B vssd1 vssd1 vccd1 vccd1 _21860_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_270_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20811_ _20811_/A vssd1 vssd1 vccd1 vccd1 _20811_/X sky130_fd_sc_hd__clkbuf_2
X_21791_ _21791_/A _21791_/B vssd1 vssd1 vccd1 vccd1 _21792_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23530_ _23530_/CLK _23530_/D vssd1 vssd1 vccd1 vccd1 _23530_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_20742_ _20757_/A _20742_/B _20742_/C vssd1 vssd1 vccd1 vccd1 _20742_/X sky130_fd_sc_hd__or3_1
XFILLER_169_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_357_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23461_ _23903_/CLK _23461_/D vssd1 vssd1 vccd1 vccd1 _23461_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20673_ _20763_/A vssd1 vssd1 vccd1 vccd1 _20673_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22412_ _23449_/CLK _22412_/D vssd1 vssd1 vccd1 vccd1 _22412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_338_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23392_ _23554_/CLK _23392_/D vssd1 vssd1 vccd1 vccd1 _23392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22343_ _23544_/CLK _22343_/D vssd1 vssd1 vccd1 vccd1 _22343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_313_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22274_ _23538_/CLK _22274_/D vssd1 vssd1 vccd1 vccd1 _22274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21225_ _21225_/A _21227_/B vssd1 vssd1 vccd1 vccd1 _21225_/Y sky130_fd_sc_hd__nand2_1
XFILLER_104_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_305_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21156_ _20700_/A _21140_/X _21142_/X _20509_/D _21135_/X vssd1 vssd1 vccd1 vccd1
+ _21156_/X sky130_fd_sc_hd__a221o_1
XFILLER_78_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_320_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20107_ _20120_/A _20107_/B _20107_/C vssd1 vssd1 vccd1 vccd1 _23642_/D sky130_fd_sc_hd__nor3_1
XFILLER_291_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21087_ _21083_/X _21085_/Y _21086_/X vssd1 vssd1 vccd1 vccd1 _21087_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_259_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20038_ _20048_/B _20048_/C _20037_/X vssd1 vssd1 vccd1 vccd1 _23623_/D sky130_fd_sc_hd__o21ba_1
XFILLER_246_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12860_ _12897_/A _12860_/B vssd1 vssd1 vccd1 vccd1 _12860_/X sky130_fd_sc_hd__or2_1
XFILLER_248_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11811_ _11630_/A _11802_/X _11806_/X _11808_/X _11810_/X vssd1 vssd1 vccd1 vccd1
+ _11811_/X sky130_fd_sc_hd__a32o_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _12784_/A _12790_/X _11631_/X vssd1 vssd1 vccd1 vccd1 _12791_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21989_ _21989_/A _21989_/B vssd1 vssd1 vccd1 vccd1 _21989_/Y sky130_fd_sc_hd__xnor2_4
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _15048_/A vssd1 vssd1 vccd1 vccd1 _14530_/X sky130_fd_sc_hd__clkbuf_4
X_11742_ _11742_/A vssd1 vssd1 vccd1 vccd1 _12009_/A sky130_fd_sc_hd__buf_4
XFILLER_214_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23728_ _23861_/CLK _23728_/D vssd1 vssd1 vccd1 vccd1 _23728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14609_/A _20986_/A vssd1 vssd1 vccd1 vccd1 _14906_/A sky130_fd_sc_hd__nor2_2
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _22794_/Q _22762_/Q _22663_/Q _22730_/Q _12709_/A _12793_/A vssd1 vssd1 vccd1
+ vccd1 _11674_/B sky130_fd_sc_hd__mux4_2
XFILLER_230_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23659_ _23818_/CLK _23659_/D vssd1 vssd1 vccd1 vccd1 _23659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16200_ _18769_/A vssd1 vssd1 vccd1 vccd1 _16200_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13412_ _13412_/A vssd1 vssd1 vccd1 vccd1 _20214_/A sky130_fd_sc_hd__buf_6
XFILLER_329_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17180_ _21888_/A vssd1 vssd1 vccd1 vccd1 _17180_/X sky130_fd_sc_hd__buf_12
XFILLER_328_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14392_ _14896_/A vssd1 vssd1 vccd1 vccd1 _14520_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_344_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16131_ _16131_/A _16131_/B vssd1 vssd1 vccd1 vccd1 _16131_/Y sky130_fd_sc_hd__nor2_1
X_13343_ _13518_/A _13343_/B _13380_/A vssd1 vssd1 vccd1 vccd1 _13344_/A sky130_fd_sc_hd__nor3_1
XFILLER_316_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_294_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_344_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16062_ _23617_/Q _14450_/A _14455_/A _23649_/Q vssd1 vssd1 vccd1 vccd1 _16062_/X
+ sky130_fd_sc_hd__o22a_2
X_13274_ _11403_/X _13273_/Y _23907_/Q _11486_/B vssd1 vssd1 vccd1 vccd1 _13319_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_108_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15013_ _15020_/S _15012_/Y _14630_/X vssd1 vssd1 vccd1 vccd1 _15013_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12225_ _12387_/A _12225_/B vssd1 vssd1 vccd1 vccd1 _12225_/X sky130_fd_sc_hd__or2_1
XFILLER_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_335_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19821_ _19821_/A vssd1 vssd1 vccd1 vccd1 _23546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_296_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12156_ _12156_/A _12156_/B _12156_/C vssd1 vssd1 vccd1 vccd1 _20264_/A sky130_fd_sc_hd__nand3_4
XFILLER_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_312_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_311_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_340_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_296_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11107_ _14176_/A _15176_/A vssd1 vssd1 vccd1 vccd1 _14133_/B sky130_fd_sc_hd__nor2_1
X_19752_ _19239_/X _23516_/Q _19754_/S vssd1 vssd1 vccd1 vccd1 _19753_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16964_ _16981_/A vssd1 vssd1 vccd1 vccd1 _17318_/S sky130_fd_sc_hd__buf_2
X_12087_ _12087_/A _12134_/A _13765_/B vssd1 vssd1 vccd1 vccd1 _12087_/X sky130_fd_sc_hd__or3_1
XFILLER_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18703_ _18703_/A vssd1 vssd1 vccd1 vccd1 _23078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_351_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15915_ _16034_/A _15915_/B vssd1 vssd1 vccd1 vccd1 _15920_/A sky130_fd_sc_hd__or2_1
X_19683_ _19683_/A vssd1 vssd1 vccd1 vccd1 _23485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16895_ _19245_/A vssd1 vssd1 vccd1 vccd1 _16895_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_264_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18634_ _23048_/Q _17556_/X _18636_/S vssd1 vssd1 vccd1 vccd1 _18635_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15846_ _14755_/X _15834_/X _15845_/X vssd1 vssd1 vccd1 vccd1 _15846_/Y sky130_fd_sc_hd__o21ai_4
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18565_ _18565_/A vssd1 vssd1 vccd1 vccd1 _23017_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12989_ _13212_/A _12989_/B vssd1 vssd1 vccd1 vccd1 _12989_/Y sky130_fd_sc_hd__nand2_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15777_ _15752_/X _15753_/Y _15776_/X _15818_/A vssd1 vssd1 vccd1 vccd1 _15777_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17516_ _22665_/Q _16268_/X _17516_/S vssd1 vssd1 vccd1 vccd1 _17517_/A sky130_fd_sc_hd__mux2_1
X_14728_ _22916_/Q _14728_/B vssd1 vssd1 vccd1 vccd1 _14728_/X sky130_fd_sc_hd__and2_1
X_18496_ _22993_/Q _18505_/B vssd1 vssd1 vccd1 vccd1 _18496_/Y sky130_fd_sc_hd__nand2_1
XFILLER_205_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17447_ _17447_/A vssd1 vssd1 vccd1 vccd1 _22634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14659_ _14655_/X _14658_/X _14852_/S vssd1 vssd1 vccd1 vccd1 _14659_/X sky130_fd_sc_hd__mux2_2
XFILLER_159_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17378_ _22609_/Q _14148_/C _17380_/S vssd1 vssd1 vccd1 vccd1 _17379_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19117_ _19117_/A vssd1 vssd1 vccd1 vccd1 _23247_/D sky130_fd_sc_hd__clkbuf_1
X_16329_ _15168_/X _22332_/Q _16333_/S vssd1 vssd1 vccd1 vccd1 _16330_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_334_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19048_ _19048_/A vssd1 vssd1 vccd1 vccd1 _23217_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_303_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_331_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21010_ _21023_/A vssd1 vssd1 vccd1 vccd1 _21010_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput289 _14092_/X vssd1 vssd1 vccd1 vccd1 addr0[4] sky130_fd_sc_hd__buf_2
XFILLER_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_303_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_7 _17296_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22961_ _22961_/CLK _22961_/D vssd1 vssd1 vccd1 vccd1 _22961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21912_ _21885_/A _21884_/A _21883_/Y vssd1 vssd1 vccd1 vccd1 _21913_/B sky130_fd_sc_hd__o21a_1
XFILLER_83_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22892_ _22893_/CLK _22892_/D vssd1 vssd1 vccd1 vccd1 _22892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21843_ _20303_/A _21900_/B _15661_/B _21842_/X vssd1 vssd1 vccd1 vccd1 _21844_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_167_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21774_ _13432_/A _13432_/B _21517_/B _15531_/X vssd1 vssd1 vccd1 vccd1 _21774_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_24_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23513_ _23546_/CLK _23513_/D vssd1 vssd1 vccd1 vccd1 _23513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20725_ _15929_/X _20724_/X _20702_/X vssd1 vssd1 vccd1 vccd1 _20725_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_11_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23444_ _23444_/CLK _23444_/D vssd1 vssd1 vccd1 vccd1 _23444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20656_ _21720_/A _20642_/X _20649_/X vssd1 vssd1 vccd1 vccd1 _20656_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_338_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_353_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23375_ _23407_/CLK _23375_/D vssd1 vssd1 vccd1 vccd1 _23375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20587_ _20895_/A vssd1 vssd1 vccd1 vccd1 _20966_/A sky130_fd_sc_hd__buf_6
XFILLER_319_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_314_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_302_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22326_ _23558_/CLK _22326_/D vssd1 vssd1 vccd1 vccd1 _22326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_353_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_325_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_313_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_341_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_307_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_340_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22257_ _22257_/A _22257_/B vssd1 vssd1 vccd1 vccd1 _22257_/X sky130_fd_sc_hd__or2_1
XFILLER_341_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_322_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12010_ _22275_/Q _23091_/Q _23507_/Q _22436_/Q _12008_/X _12009_/X vssd1 vssd1 vccd1
+ vccd1 _12011_/B sky130_fd_sc_hd__mux4_1
XFILLER_3_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21208_ _14196_/A _14834_/X _21214_/S vssd1 vssd1 vccd1 vccd1 _21209_/B sky130_fd_sc_hd__mux2_8
X_22188_ _22148_/Y _22153_/B _22150_/B vssd1 vssd1 vccd1 vccd1 _22189_/B sky130_fd_sc_hd__o21ai_1
XFILLER_132_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_321_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21139_ _21168_/A vssd1 vssd1 vccd1 vccd1 _21139_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_293_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13961_ _13960_/X _15453_/A _13603_/X _21719_/A vssd1 vssd1 vccd1 vccd1 _13962_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_93_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12912_ _11277_/A _12902_/X _12911_/X _12864_/A vssd1 vssd1 vccd1 vccd1 _20334_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15700_ _23929_/Q vssd1 vssd1 vccd1 vccd1 _21888_/A sky130_fd_sc_hd__buf_2
XFILLER_247_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16680_ _16680_/A _16808_/A vssd1 vssd1 vccd1 vccd1 _16810_/B sky130_fd_sc_hd__nand2_1
X_13892_ _13892_/A _15187_/A vssd1 vssd1 vccd1 vccd1 _13892_/Y sky130_fd_sc_hd__nor2_8
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12843_ _12843_/A vssd1 vssd1 vccd1 vccd1 _12843_/X sky130_fd_sc_hd__buf_6
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15631_ _15631_/A vssd1 vssd1 vccd1 vccd1 _15673_/A sky130_fd_sc_hd__buf_2
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18350_ _18358_/A _18350_/B _18351_/B vssd1 vssd1 vccd1 vccd1 _22943_/D sky130_fd_sc_hd__nor3_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15562_ _14215_/A _21244_/A _15561_/X _11099_/A vssd1 vssd1 vccd1 vccd1 _15562_/X
+ sky130_fd_sc_hd__o22a_1
X_12774_ _12891_/A _13798_/A vssd1 vssd1 vccd1 vccd1 _12774_/Y sky130_fd_sc_hd__nand2_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14513_/A vssd1 vssd1 vccd1 vccd1 _14513_/X sky130_fd_sc_hd__clkbuf_2
X_17301_ _22193_/A _17300_/X _17318_/S vssd1 vssd1 vccd1 vccd1 _17301_/X sky130_fd_sc_hd__mux2_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_48_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23409_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11725_ _11698_/A _11724_/X _11706_/X vssd1 vssd1 vccd1 vccd1 _11725_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18281_ _18317_/A _18286_/C vssd1 vssd1 vccd1 vccd1 _18281_/Y sky130_fd_sc_hd__nor2_1
X_15493_ _15583_/A _15492_/X _12065_/A vssd1 vssd1 vccd1 vccd1 _15493_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_261_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14444_ _14730_/A vssd1 vssd1 vccd1 vccd1 _15346_/A sky130_fd_sc_hd__buf_6
X_17232_ _17232_/A vssd1 vssd1 vccd1 vccd1 _17232_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_348_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11656_ _12842_/A _11643_/X _11655_/X _12797_/A vssd1 vssd1 vccd1 vccd1 _11656_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_302_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17163_ _17163_/A _17163_/B vssd1 vssd1 vccd1 vccd1 _17163_/X sky130_fd_sc_hd__or2_1
XFILLER_317_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14375_ _14665_/S _14369_/X _14381_/B vssd1 vssd1 vccd1 vccd1 _14375_/Y sky130_fd_sc_hd__o21bai_1
X_11587_ _11587_/A _11587_/B vssd1 vssd1 vccd1 vccd1 _11587_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_344_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16114_ _16114_/A _16151_/C vssd1 vssd1 vccd1 vccd1 _16115_/B sky130_fd_sc_hd__xnor2_2
X_13326_ _13629_/A _13330_/B _12809_/Y vssd1 vssd1 vccd1 vccd1 _13327_/B sky130_fd_sc_hd__a21bo_1
XFILLER_127_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17094_ _17268_/A vssd1 vssd1 vccd1 vccd1 _17094_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_346_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16045_ _21077_/A _15663_/X _16043_/Y _16044_/Y vssd1 vssd1 vccd1 vccd1 _16045_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_331_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13257_ _14393_/A _13254_/X _13256_/X vssd1 vssd1 vccd1 vccd1 _13257_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_170_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12208_ _12383_/A _12208_/B vssd1 vssd1 vccd1 vccd1 _12208_/X sky130_fd_sc_hd__or2_1
X_13188_ _13188_/A _13543_/A vssd1 vssd1 vccd1 vccd1 _13574_/A sky130_fd_sc_hd__nor2_4
XFILLER_313_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19804_ _23539_/Q _19210_/A _19804_/S vssd1 vssd1 vccd1 vccd1 _19805_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12139_ _12139_/A _12139_/B vssd1 vssd1 vccd1 vccd1 _12139_/X sky130_fd_sc_hd__or2_1
XFILLER_297_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17996_ _22840_/Q _17990_/X _17986_/X _17995_/X _17983_/X vssd1 vssd1 vccd1 vccd1
+ _17996_/X sky130_fd_sc_hd__a221o_1
XFILLER_300_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19735_ _19213_/X _23508_/Q _19743_/S vssd1 vssd1 vccd1 vccd1 _19736_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16947_ _17022_/B vssd1 vssd1 vccd1 vccd1 _16947_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19666_ _19666_/A vssd1 vssd1 vccd1 vccd1 _23477_/D sky130_fd_sc_hd__clkbuf_1
X_16878_ _16878_/A vssd1 vssd1 vccd1 vccd1 _22540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18617_ _16905_/X _23041_/Q _18619_/S vssd1 vssd1 vccd1 vccd1 _18618_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15829_ _15924_/C _15829_/B vssd1 vssd1 vccd1 vccd1 _15829_/Y sky130_fd_sc_hd__nor2_4
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19597_ _23447_/Q _19223_/A _19599_/S vssd1 vssd1 vccd1 vccd1 _19598_/A sky130_fd_sc_hd__mux2_1
XFILLER_280_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18548_ _18536_/A _18542_/A _18545_/Y _18547_/X vssd1 vssd1 vccd1 vccd1 _23011_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18479_ _18467_/X _18478_/Y _18476_/X vssd1 vssd1 vccd1 vccd1 _22987_/D sky130_fd_sc_hd__a21oi_1
XFILLER_221_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20510_ _23714_/Q _20517_/B _20510_/C vssd1 vssd1 vccd1 vccd1 _20515_/A sky130_fd_sc_hd__and3_1
XFILLER_339_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21490_ _21634_/A vssd1 vssd1 vccd1 vccd1 _22061_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20441_ _20630_/A _20428_/X _20440_/X _20433_/X vssd1 vssd1 vccd1 vccd1 _23695_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_347_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23160_ _23420_/CLK _23160_/D vssd1 vssd1 vccd1 vccd1 _23160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20372_ _20379_/A _21173_/A vssd1 vssd1 vccd1 vccd1 _20372_/Y sky130_fd_sc_hd__nand2_1
XFILLER_323_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22111_ _23839_/Q _22190_/B vssd1 vssd1 vccd1 vccd1 _22111_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23091_ _23507_/CLK _23091_/D vssd1 vssd1 vccd1 vccd1 _23091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22042_ _22161_/A _22042_/B vssd1 vssd1 vccd1 vccd1 _22042_/Y sky130_fd_sc_hd__nand2_1
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22944_ _22947_/CLK _22944_/D vssd1 vssd1 vccd1 vccd1 _22944_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_290_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22875_ _22893_/CLK _22875_/D vssd1 vssd1 vccd1 vccd1 _22875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_357_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21826_ _21826_/A _21829_/A vssd1 vssd1 vccd1 vccd1 _21826_/Y sky130_fd_sc_hd__nand2_1
XFILLER_243_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_325_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_357_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21757_ _21734_/A _21733_/B _21733_/A vssd1 vssd1 vccd1 vccd1 _21758_/B sky130_fd_sc_hd__o21ba_1
XFILLER_12_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11510_ _15929_/A _11500_/X _11509_/X _13765_/A vssd1 vssd1 vccd1 vccd1 _11511_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20708_ _20708_/A _20731_/B vssd1 vssd1 vccd1 vccd1 _20711_/B sky130_fd_sc_hd__and2_2
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12490_ _22455_/Q _22615_/Q _22294_/Q _23430_/Q _12475_/X _12476_/X vssd1 vssd1 vccd1
+ vccd1 _12490_/X sky130_fd_sc_hd__mux4_1
X_21688_ _21725_/B _21688_/B vssd1 vssd1 vccd1 vccd1 _21801_/A sky130_fd_sc_hd__xnor2_2
XFILLER_200_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_339_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11441_ _13091_/A vssd1 vssd1 vccd1 vccd1 _13107_/A sky130_fd_sc_hd__buf_2
XFILLER_221_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23427_ _23491_/CLK _23427_/D vssd1 vssd1 vccd1 vccd1 _23427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20639_ _20639_/A vssd1 vssd1 vccd1 vccd1 _20641_/A sky130_fd_sc_hd__inv_2
XFILLER_326_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14160_ _14394_/A vssd1 vssd1 vccd1 vccd1 _14160_/X sky130_fd_sc_hd__buf_2
X_23358_ _23547_/CLK _23358_/D vssd1 vssd1 vccd1 vccd1 _23358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_299_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11372_ _13287_/A _11372_/B vssd1 vssd1 vccd1 vccd1 _11372_/X sky130_fd_sc_hd__or2_1
XFILLER_354_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_326_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13111_ _23905_/Q _13185_/S _11403_/A _13110_/Y vssd1 vssd1 vccd1 vccd1 _13542_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22309_ _23446_/CLK _22309_/D vssd1 vssd1 vccd1 vccd1 _22309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14091_ _14091_/A vssd1 vssd1 vccd1 vccd1 _14091_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23289_ _23419_/CLK _23289_/D vssd1 vssd1 vccd1 vccd1 _23289_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_166_wb_clk_i _23917_/CLK vssd1 vssd1 vccd1 vccd1 _23874_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_341_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_313_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13042_ _22384_/Q _22416_/Q _22705_/Q _23072_/Q _11432_/A _13037_/X vssd1 vssd1 vccd1
+ vccd1 _13042_/X sky130_fd_sc_hd__mux4_2
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_332_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17850_ _17861_/A vssd1 vssd1 vccd1 vccd1 _17859_/S sky130_fd_sc_hd__buf_2
XFILLER_182_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_293_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16801_ _16804_/A _16801_/B vssd1 vssd1 vccd1 vccd1 _16802_/A sky130_fd_sc_hd__or2_1
XTAP_6997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17781_ _22766_/Q _17614_/X _17787_/S vssd1 vssd1 vccd1 vccd1 _17782_/A sky130_fd_sc_hd__mux2_1
X_14993_ _23722_/Q _23852_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _14993_/X sky130_fd_sc_hd__mux2_2
X_19520_ _19520_/A vssd1 vssd1 vccd1 vccd1 _23412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16732_ _16741_/A _16732_/B vssd1 vssd1 vccd1 vccd1 _16733_/A sky130_fd_sc_hd__or2_1
XFILLER_219_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13944_ _23920_/Q vssd1 vssd1 vccd1 vccd1 _13945_/B sky130_fd_sc_hd__buf_8
XFILLER_262_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19451_ _23382_/Q _18827_/X _19455_/S vssd1 vssd1 vccd1 vccd1 _19452_/A sky130_fd_sc_hd__mux2_1
X_16663_ _16663_/A vssd1 vssd1 vccd1 vccd1 _22478_/D sky130_fd_sc_hd__clkbuf_1
X_13875_ _13875_/A _13875_/B _13875_/C vssd1 vssd1 vccd1 vccd1 _13875_/X sky130_fd_sc_hd__and3_1
XFILLER_62_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18402_ _22962_/Q _18402_/B vssd1 vssd1 vccd1 vccd1 _18409_/C sky130_fd_sc_hd__and2_1
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12826_ _22380_/Q _22412_/Q _22701_/Q _23068_/Q _12825_/X _12672_/A vssd1 vssd1 vccd1
+ vccd1 _12826_/X sky130_fd_sc_hd__mux4_1
XFILLER_250_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15614_ _15367_/A _15608_/X _15613_/X vssd1 vssd1 vccd1 vccd1 _15614_/Y sky130_fd_sc_hd__o21ai_1
X_19382_ _19382_/A vssd1 vssd1 vccd1 vccd1 _23351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_250_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16594_ _16594_/A vssd1 vssd1 vccd1 vccd1 _22447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_349_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18333_ _18358_/A _18333_/B _18334_/B vssd1 vssd1 vccd1 vccd1 _22937_/D sky130_fd_sc_hd__nor3_1
X_12757_ _23223_/Q _23191_/Q _23159_/Q _23127_/Q _12755_/X _12756_/X vssd1 vssd1 vccd1
+ vccd1 _12758_/B sky130_fd_sc_hd__mux4_2
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15545_ _15798_/A _15540_/X _15542_/X _14621_/A _15544_/Y vssd1 vssd1 vccd1 vccd1
+ _15545_/X sky130_fd_sc_hd__o221a_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _22465_/Q _22625_/Q _11708_/S vssd1 vssd1 vccd1 vccd1 _11708_/X sky130_fd_sc_hd__mux2_1
XFILLER_348_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18264_ _18264_/A _18264_/B _18264_/C vssd1 vssd1 vccd1 vccd1 _22916_/D sky130_fd_sc_hd__nor3_1
X_15476_ _15476_/A vssd1 vssd1 vccd1 vccd1 _22274_/D sky130_fd_sc_hd__clkbuf_1
X_12688_ _12836_/A _12686_/X _12687_/X vssd1 vssd1 vccd1 vccd1 _12688_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_202_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17215_ _17283_/A vssd1 vssd1 vccd1 vccd1 _17215_/X sky130_fd_sc_hd__clkbuf_2
X_14427_ _15066_/B _14434_/B vssd1 vssd1 vccd1 vccd1 _15148_/A sky130_fd_sc_hd__nor2_1
XFILLER_336_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11639_ _12007_/A _11639_/B vssd1 vssd1 vccd1 vccd1 _11639_/X sky130_fd_sc_hd__or2_1
XFILLER_175_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18195_ _18195_/A _18195_/B _18195_/C vssd1 vssd1 vccd1 vccd1 _18195_/Y sky130_fd_sc_hd__nand3_1
XFILLER_129_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17146_ _17220_/B vssd1 vssd1 vccd1 vccd1 _17170_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14358_ _14358_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _14358_/Y sky130_fd_sc_hd__nand2_1
XFILLER_344_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_289_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_317_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13309_ _13316_/A _13316_/B _13555_/A vssd1 vssd1 vccd1 vccd1 _13309_/X sky130_fd_sc_hd__a21o_1
X_17077_ _13939_/B _17076_/X _17087_/S vssd1 vssd1 vccd1 vccd1 _17077_/X sky130_fd_sc_hd__mux2_1
XFILLER_305_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14289_ _14287_/Y _13362_/B _14330_/S vssd1 vssd1 vccd1 vccd1 _14373_/A sky130_fd_sc_hd__mux2_1
XFILLER_332_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_289_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16028_ _16028_/A _16028_/B vssd1 vssd1 vccd1 vccd1 _16028_/Y sky130_fd_sc_hd__nand2_1
XFILLER_332_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_300_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater501 _13454_/Y vssd1 vssd1 vccd1 vccd1 output442/A sky130_fd_sc_hd__buf_6
XFILLER_284_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_301_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17979_ _18029_/A vssd1 vssd1 vccd1 vccd1 _17979_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_273_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19718_ _19718_/A vssd1 vssd1 vccd1 vccd1 _23500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20990_ _21051_/A vssd1 vssd1 vccd1 vccd1 _21064_/B sky130_fd_sc_hd__buf_4
XFILLER_226_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_348_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19649_ _19194_/X _23470_/Q _19649_/S vssd1 vssd1 vccd1 vccd1 _19650_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22660_ _23450_/CLK _22660_/D vssd1 vssd1 vccd1 vccd1 _22660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21611_ _13945_/B _21305_/X _21610_/X _21581_/X vssd1 vssd1 vccd1 vccd1 _23920_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_339_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22591_ _22977_/CLK _22591_/D vssd1 vssd1 vccd1 vccd1 _22591_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_205_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21542_ _21542_/A _21546_/B _21542_/C vssd1 vssd1 vccd1 vccd1 _21542_/X sky130_fd_sc_hd__and3_1
XFILLER_355_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21473_ _21472_/A _21472_/C _21472_/B vssd1 vssd1 vccd1 vccd1 _21473_/Y sky130_fd_sc_hd__o21ai_1
X_23212_ _23950_/A _23212_/D vssd1 vssd1 vccd1 vccd1 _23212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_342_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20424_ _23689_/Q _20429_/B vssd1 vssd1 vccd1 vccd1 _20424_/X sky130_fd_sc_hd__or2_1
XFILLER_119_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_335_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23143_ _23367_/CLK _23143_/D vssd1 vssd1 vccd1 vccd1 _23143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_323_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20355_ _20355_/A _20355_/B vssd1 vssd1 vccd1 vccd1 _20355_/Y sky130_fd_sc_hd__nand2_1
XFILLER_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_311_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23074_ _23586_/CLK _23074_/D vssd1 vssd1 vccd1 vccd1 _23074_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20286_ _20272_/X _20660_/A _20284_/X _20285_/X vssd1 vssd1 vccd1 vccd1 _23667_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_6227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_304_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22025_ _22025_/A _22025_/B vssd1 vssd1 vccd1 vccd1 _22025_/Y sky130_fd_sc_hd__nand2_1
XTAP_6249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11990_ _12842_/A _11987_/X _11989_/X _11681_/X vssd1 vssd1 vccd1 vccd1 _11990_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_229_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_291_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22927_ _22929_/CLK _22927_/D vssd1 vssd1 vccd1 vccd1 _22927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13660_ _14211_/A vssd1 vssd1 vccd1 vccd1 _13665_/A sky130_fd_sc_hd__inv_2
X_22858_ _22908_/CLK _22858_/D vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dfxtp_1
XFILLER_231_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_348_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _13340_/A _12611_/B vssd1 vssd1 vccd1 vccd1 _15198_/A sky130_fd_sc_hd__nor2_1
XFILLER_213_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21809_ _21809_/A _21809_/B vssd1 vssd1 vccd1 vccd1 _21810_/B sky130_fd_sc_hd__nor2_1
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _13018_/D _13601_/B _13015_/B vssd1 vssd1 vccd1 vccd1 _13592_/B sky130_fd_sc_hd__o21ba_1
XFILLER_231_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22789_ _22789_/CLK _22789_/D vssd1 vssd1 vccd1 vccd1 _22789_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _15330_/A vssd1 vssd1 vccd1 vccd1 _15330_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_358_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ _11844_/A _12532_/Y _12534_/Y _12541_/X _11240_/A vssd1 vssd1 vccd1 vccd1
+ _12542_/X sky130_fd_sc_hd__o311a_1
XFILLER_197_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_346_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15261_ _23822_/Q vssd1 vssd1 vccd1 vccd1 _21630_/A sky130_fd_sc_hd__buf_2
X_12473_ _22262_/Q _23078_/Q _23494_/Q _22423_/Q _11919_/A _12216_/A vssd1 vssd1 vccd1
+ vccd1 _12474_/B sky130_fd_sc_hd__mux4_2
XFILLER_12_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14212_ _22978_/Q _14137_/A _14980_/A input215/X vssd1 vssd1 vccd1 vccd1 _17655_/A
+ sky130_fd_sc_hd__a22oi_4
X_17000_ _17000_/A vssd1 vssd1 vccd1 vccd1 _17000_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11424_ _11424_/A _11424_/B vssd1 vssd1 vccd1 vccd1 _11424_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_326_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15192_ _15538_/A _15192_/B vssd1 vssd1 vccd1 vccd1 _15192_/Y sky130_fd_sc_hd__nand2_1
XFILLER_327_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_354_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14143_ _14211_/A _16945_/A _14211_/C vssd1 vssd1 vccd1 vccd1 _17648_/A sky130_fd_sc_hd__and3_1
X_11355_ _11288_/X _11326_/X _11340_/X _11354_/X vssd1 vssd1 vccd1 vccd1 _11355_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_314_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_287_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14074_ _14074_/A _14074_/B _14089_/B _14074_/D vssd1 vssd1 vccd1 vccd1 _14074_/X
+ sky130_fd_sc_hd__or4_1
X_18951_ _16819_/X _23174_/Q _18957_/S vssd1 vssd1 vccd1 vccd1 _18952_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_314_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11286_ _12707_/A vssd1 vssd1 vccd1 vccd1 _12745_/A sky130_fd_sc_hd__buf_2
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17902_ _17991_/A _17986_/A vssd1 vssd1 vccd1 vccd1 _17959_/A sky130_fd_sc_hd__and2_2
X_13025_ _14307_/B vssd1 vssd1 vccd1 vccd1 _13026_/B sky130_fd_sc_hd__inv_2
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_295_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18882_ _18882_/A vssd1 vssd1 vccd1 vccd1 _23143_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_343_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_294_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17833_ _22789_/Q _17585_/X _17837_/S vssd1 vssd1 vccd1 vccd1 _17834_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_294_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17764_ _17764_/A vssd1 vssd1 vccd1 vccd1 _22758_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14976_ _21431_/A _14976_/B vssd1 vssd1 vccd1 vccd1 _14977_/B sky130_fd_sc_hd__nor2_1
XFILLER_281_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19503_ _19191_/X _23405_/Q _19505_/S vssd1 vssd1 vccd1 vccd1 _19504_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_63_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23573_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_263_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16715_ _16715_/A vssd1 vssd1 vccd1 vccd1 _22492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_281_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13927_ _13920_/A _13920_/B _12287_/A vssd1 vssd1 vccd1 vccd1 _13928_/B sky130_fd_sc_hd__a21o_1
X_17695_ _17717_/A vssd1 vssd1 vccd1 vccd1 _17704_/S sky130_fd_sc_hd__buf_4
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_401 _13988_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_412 _14033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19434_ _19434_/A vssd1 vssd1 vccd1 vccd1 _23374_/D sky130_fd_sc_hd__clkbuf_1
X_16646_ _16646_/A vssd1 vssd1 vccd1 vccd1 _22470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_423 _14014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13858_ _13858_/A _13875_/B _13875_/C vssd1 vssd1 vccd1 vccd1 _13858_/X sky130_fd_sc_hd__and3_1
XINSDIODE2_434 _23882_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_445 _23945_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_456 _17305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19365_ _19365_/A vssd1 vssd1 vccd1 vccd1 _23343_/D sky130_fd_sc_hd__clkbuf_1
X_12809_ _13534_/A _12809_/B vssd1 vssd1 vccd1 vccd1 _12809_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_467 _22146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16577_ _15710_/X _22440_/Q _16579_/S vssd1 vssd1 vccd1 vccd1 _16578_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_478 _20499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13789_ _13789_/A vssd1 vssd1 vccd1 vccd1 _13829_/B sky130_fd_sc_hd__buf_2
XFILLER_31_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_489 _13956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18316_ _22930_/Q _22931_/Q _22932_/Q _18316_/D vssd1 vssd1 vccd1 vccd1 _18323_/C
+ sky130_fd_sc_hd__and4_2
XFILLER_231_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15528_ _23926_/Q vssd1 vssd1 vccd1 vccd1 _21791_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_337_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19296_ _19204_/X _23313_/Q _19300_/S vssd1 vssd1 vccd1 vccd1 _19297_/A sky130_fd_sc_hd__mux2_1
XFILLER_188_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18247_ _22910_/Q _18253_/B vssd1 vssd1 vccd1 vccd1 _18247_/X sky130_fd_sc_hd__or2_1
X_15459_ _15089_/S _14780_/X _15253_/X vssd1 vssd1 vccd1 vccd1 _15459_/X sky130_fd_sc_hd__a21o_1
XFILLER_318_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_324_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18178_ _18162_/A _18178_/B vssd1 vssd1 vccd1 vccd1 _18178_/X sky130_fd_sc_hd__and2b_1
XFILLER_116_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17129_ _17070_/A _17121_/X _17128_/X _17109_/X vssd1 vssd1 vccd1 vccd1 _17129_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_190_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_305_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20140_ _21294_/A _20140_/B vssd1 vssd1 vccd1 vccd1 _20140_/X sky130_fd_sc_hd__or2_4
XFILLER_143_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_289_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20071_ _23632_/Q _20079_/B _20071_/C vssd1 vssd1 vccd1 vccd1 _20072_/B sky130_fd_sc_hd__and3_2
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_257_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23830_ _23877_/CLK _23830_/D vssd1 vssd1 vccd1 vccd1 _23830_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23761_ _23878_/CLK _23761_/D vssd1 vssd1 vccd1 vccd1 _23761_/Q sky130_fd_sc_hd__dfxtp_4
X_20973_ _22114_/A _20966_/X _20742_/B _20970_/X vssd1 vssd1 vccd1 vccd1 _20973_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_82_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22712_ _22712_/CLK _22712_/D vssd1 vssd1 vccd1 vccd1 _22712_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23692_ _23692_/CLK _23692_/D vssd1 vssd1 vccd1 vccd1 _23692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_281_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22643_ _23585_/CLK _22643_/D vssd1 vssd1 vccd1 vccd1 _22643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_322_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22574_ _23643_/CLK _22574_/D vssd1 vssd1 vccd1 vccd1 _22574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_327_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_327_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21525_ _21546_/B _21542_/C vssd1 vssd1 vccd1 vccd1 _21528_/A sky130_fd_sc_hd__nand2_1
XFILLER_222_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_356_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_327_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21456_ _21456_/A vssd1 vssd1 vccd1 vccd1 _22019_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_309_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_294_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20407_ _20467_/A vssd1 vssd1 vccd1 vccd1 _20428_/A sky130_fd_sc_hd__buf_4
XFILLER_108_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21387_ _21400_/A _21600_/A _21384_/X _21553_/A _21386_/X vssd1 vssd1 vccd1 vccd1
+ _21425_/A sky130_fd_sc_hd__o221a_1
XFILLER_269_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23126_ _23543_/CLK _23126_/D vssd1 vssd1 vccd1 vccd1 _23126_/Q sky130_fd_sc_hd__dfxtp_1
X_11140_ _11774_/A vssd1 vssd1 vccd1 vccd1 _11141_/A sky130_fd_sc_hd__buf_4
XFILLER_351_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20338_ _23674_/Q _20338_/B vssd1 vssd1 vccd1 vccd1 _20338_/X sky130_fd_sc_hd__or2_1
XFILLER_123_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_311_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23057_ _23571_/CLK _23057_/D vssd1 vssd1 vccd1 vccd1 _23057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11071_ _23883_/Q vssd1 vssd1 vccd1 vccd1 _12345_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_6046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20269_ _20174_/X _20265_/X _20267_/Y _20268_/Y _16940_/X vssd1 vssd1 vccd1 vccd1
+ _21025_/A sky130_fd_sc_hd__o32a_4
XFILLER_249_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_295_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput101 dout0[62] vssd1 vssd1 vccd1 vccd1 input101/X sky130_fd_sc_hd__clkbuf_1
XTAP_6068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput112 dout1[14] vssd1 vssd1 vccd1 vccd1 input112/X sky130_fd_sc_hd__clkbuf_1
XTAP_5323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22008_ _22100_/A vssd1 vssd1 vccd1 vccd1 _22161_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput123 dout1[24] vssd1 vssd1 vccd1 vccd1 input123/X sky130_fd_sc_hd__clkbuf_1
XTAP_5334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput134 dout1[34] vssd1 vssd1 vccd1 vccd1 input134/X sky130_fd_sc_hd__buf_2
XTAP_5345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput145 dout1[44] vssd1 vssd1 vccd1 vccd1 input145/X sky130_fd_sc_hd__buf_2
XFILLER_292_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput156 dout1[54] vssd1 vssd1 vccd1 vccd1 input156/X sky130_fd_sc_hd__buf_2
XFILLER_237_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput167 dout1[6] vssd1 vssd1 vccd1 vccd1 input167/X sky130_fd_sc_hd__clkbuf_1
XTAP_5378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14830_ _14218_/X _15332_/A _15331_/A _13829_/B _14829_/Y vssd1 vssd1 vccd1 vccd1
+ _14830_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput178 irq[1] vssd1 vssd1 vccd1 vccd1 _20523_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 jtag_tms vssd1 vssd1 vccd1 vccd1 _18181_/A sky130_fd_sc_hd__buf_12
XFILLER_64_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11973_ _12073_/A vssd1 vssd1 vccd1 vccd1 _11973_/X sky130_fd_sc_hd__buf_4
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14761_ _14761_/A vssd1 vssd1 vccd1 vccd1 _14761_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_291_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16500_ _15710_/X _22407_/Q _16502_/S vssd1 vssd1 vccd1 vccd1 _16501_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _13786_/A _13712_/B vssd1 vssd1 vccd1 vccd1 _13713_/A sky130_fd_sc_hd__and2_4
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14692_ _14632_/Y _14681_/X _14691_/Y vssd1 vssd1 vccd1 vccd1 _14692_/X sky130_fd_sc_hd__o21a_2
X_17480_ _17480_/A vssd1 vssd1 vccd1 vccd1 _22648_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16431_ _16442_/A vssd1 vssd1 vccd1 vccd1 _16440_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_31_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13643_ _13935_/B _13935_/C _13935_/A vssd1 vssd1 vccd1 vccd1 _13942_/B sky130_fd_sc_hd__a21oi_2
XFILLER_108_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19150_ _19150_/A vssd1 vssd1 vccd1 vccd1 _23262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16362_ _15861_/X _22347_/Q _16366_/S vssd1 vssd1 vccd1 vccd1 _16363_/A sky130_fd_sc_hd__mux2_1
X_13574_ _13574_/A _13574_/B vssd1 vssd1 vccd1 vccd1 _13575_/B sky130_fd_sc_hd__xnor2_4
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18101_ _22871_/Q _18096_/X _18100_/X _18090_/X vssd1 vssd1 vccd1 vccd1 _22871_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_347_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12525_ _12532_/A _12525_/B vssd1 vssd1 vccd1 vccd1 _12525_/Y sky130_fd_sc_hd__nor2_1
X_15313_ _15097_/S _15298_/Y _15312_/X _14587_/X vssd1 vssd1 vccd1 vccd1 _15313_/X
+ sky130_fd_sc_hd__a22o_1
X_16293_ _16293_/A vssd1 vssd1 vccd1 vccd1 _22319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_318_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19081_ _19081_/A vssd1 vssd1 vccd1 vccd1 _23232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_181_wb_clk_i _23931_/CLK vssd1 vssd1 vccd1 vccd1 _23938_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_185_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_334_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18032_ _22849_/Q _18016_/X _18031_/X _18029_/X vssd1 vssd1 vccd1 vccd1 _22849_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15244_ _15244_/A _15433_/B vssd1 vssd1 vccd1 vccd1 _15244_/Y sky130_fd_sc_hd__nand2_1
XFILLER_145_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12456_ _12536_/A _12456_/B vssd1 vssd1 vccd1 vccd1 _12456_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_110_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _22830_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_346_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11407_ _12661_/A vssd1 vssd1 vccd1 vccd1 _12891_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15175_ _13833_/A _15119_/B _15111_/X _13737_/A vssd1 vssd1 vccd1 vccd1 _15176_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12387_ _12387_/A _12387_/B vssd1 vssd1 vccd1 vccd1 _12387_/X sky130_fd_sc_hd__or2_1
XFILLER_342_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14126_ _22877_/Q _18198_/B _14122_/X _14125_/Y vssd1 vssd1 vccd1 vccd1 _14126_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11338_ _13287_/A vssd1 vssd1 vccd1 vccd1 _13291_/A sky130_fd_sc_hd__buf_2
XFILLER_153_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19983_ _23608_/Q _19988_/C vssd1 vssd1 vccd1 vccd1 _19986_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_4_9_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_207_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_354_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18934_ _23167_/Q _18856_/X _18940_/S vssd1 vssd1 vccd1 vccd1 _18935_/A sky130_fd_sc_hd__mux2_1
X_14057_ input231/X _14038_/X _14056_/X vssd1 vssd1 vccd1 vccd1 _14057_/X sky130_fd_sc_hd__a21bo_4
XTAP_7270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11269_ _14178_/A _11249_/Y _11269_/S vssd1 vssd1 vccd1 vccd1 _11394_/A sky130_fd_sc_hd__mux2_4
XTAP_7281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13008_ _11515_/A _13007_/X _11537_/A vssd1 vssd1 vccd1 vccd1 _13008_/X sky130_fd_sc_hd__o21a_1
X_18865_ _18865_/A vssd1 vssd1 vccd1 vccd1 _18865_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17816_ _17816_/A vssd1 vssd1 vccd1 vccd1 _22781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_283_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18796_ _23116_/Q _18795_/X _18802_/S vssd1 vssd1 vccd1 vccd1 _18797_/A sky130_fd_sc_hd__mux2_1
XTAP_5890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17747_ _17747_/A vssd1 vssd1 vccd1 vccd1 _22750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_282_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14959_ _14941_/X _14958_/X _14520_/A vssd1 vssd1 vccd1 vccd1 _14959_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_236_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17678_ _22720_/Q _17569_/X _17682_/S vssd1 vssd1 vccd1 vccd1 _17679_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_220 _14924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_231 _15117_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_242 _18804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19417_ _19417_/A vssd1 vssd1 vccd1 vccd1 _23366_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_253 _15510_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16629_ _22463_/Q _16236_/X _16629_/S vssd1 vssd1 vccd1 vccd1 _16630_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_264 _15651_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_275 _21916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_286 _15959_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_356_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19348_ _23336_/Q _18782_/X _19350_/S vssd1 vssd1 vccd1 vccd1 _19349_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_297 _15990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_337_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19279_ _19279_/A vssd1 vssd1 vccd1 vccd1 _23305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_353_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_338_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21310_ _21683_/A vssd1 vssd1 vccd1 vccd1 _21814_/B sky130_fd_sc_hd__buf_2
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22290_ _23522_/CLK _22290_/D vssd1 vssd1 vccd1 vccd1 _22290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_346_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_352_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21241_ _13775_/A _21229_/X _21240_/Y _21236_/X vssd1 vssd1 vccd1 vccd1 _23893_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21172_ _23872_/Q _21168_/X _21171_/X _21163_/X vssd1 vssd1 vccd1 vccd1 _23872_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_264_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20123_ _23647_/Q _23644_/Q _20123_/C _20126_/D vssd1 vssd1 vccd1 vccd1 _20131_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_104_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20054_ _23628_/Q vssd1 vssd1 vccd1 vccd1 _20066_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23813_ _23824_/CLK _23813_/D vssd1 vssd1 vccd1 vccd1 _23813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23744_ _23915_/CLK _23744_/D vssd1 vssd1 vccd1 vccd1 _23744_/Q sky130_fd_sc_hd__dfxtp_1
X_20956_ _23801_/Q _20953_/X _20955_/X _20948_/X vssd1 vssd1 vccd1 vccd1 _23801_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_289_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23675_ _23706_/CLK _23675_/D vssd1 vssd1 vccd1 vccd1 _23675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20887_ _20887_/A vssd1 vssd1 vccd1 vccd1 _23779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22626_ _23568_/CLK _22626_/D vssd1 vssd1 vccd1 vccd1 _22626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22557_ _22977_/CLK _22557_/D vssd1 vssd1 vccd1 vccd1 _22557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_344_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12310_ _12303_/Y _12305_/Y _12307_/Y _12309_/Y _11242_/A vssd1 vssd1 vccd1 vccd1
+ _12311_/C sky130_fd_sc_hd__o221a_1
X_21508_ _21676_/B vssd1 vssd1 vccd1 vccd1 _21515_/B sky130_fd_sc_hd__buf_2
XFILLER_328_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13290_ _22805_/Q _22773_/Q _22674_/Q _22741_/Q _11461_/A _11365_/X vssd1 vssd1 vccd1
+ vccd1 _13291_/B sky130_fd_sc_hd__mux4_1
XFILLER_344_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22488_ _23841_/CLK _22488_/D vssd1 vssd1 vccd1 vccd1 _22488_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_315_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12241_ _12241_/A _12241_/B vssd1 vssd1 vccd1 vccd1 _12241_/Y sky130_fd_sc_hd__nor2_1
X_21439_ _21379_/X _21430_/X _21438_/X _21984_/A vssd1 vssd1 vccd1 vccd1 _21439_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_108_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12172_ _11946_/X _12161_/X _12169_/X _13615_/A _12171_/Y vssd1 vssd1 vccd1 vccd1
+ _13349_/A sky130_fd_sc_hd__o221a_4
XFILLER_107_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11123_ _12660_/A vssd1 vssd1 vccd1 vccd1 _11124_/A sky130_fd_sc_hd__buf_4
X_23109_ _23527_/CLK _23109_/D vssd1 vssd1 vccd1 vccd1 _23109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_311_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16980_ _16980_/A vssd1 vssd1 vccd1 vccd1 _21317_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_111_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_296_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15931_ _15931_/A vssd1 vssd1 vccd1 vccd1 _16084_/A sky130_fd_sc_hd__buf_2
XFILLER_153_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18650_ _23055_/Q _17578_/X _18658_/S vssd1 vssd1 vccd1 vccd1 _18651_/A sky130_fd_sc_hd__mux2_1
X_15862_ _15861_/X _22283_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15863_/A sky130_fd_sc_hd__mux2_1
XTAP_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_329_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17601_ _18827_/A vssd1 vssd1 vccd1 vccd1 _17601_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14813_ _14813_/A vssd1 vssd1 vccd1 vccd1 _22263_/D sky130_fd_sc_hd__clkbuf_1
X_18581_ _18581_/A vssd1 vssd1 vccd1 vccd1 _23024_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _15891_/A _15793_/B vssd1 vssd1 vccd1 vccd1 _15818_/B sky130_fd_sc_hd__nand2_2
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17532_ _22672_/Q _16291_/X _17538_/S vssd1 vssd1 vccd1 vccd1 _17533_/A sky130_fd_sc_hd__mux2_1
XFILLER_280_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ _23655_/Q _14486_/X _14740_/X _14743_/X _15593_/A vssd1 vssd1 vccd1 vccd1
+ _14744_/X sky130_fd_sc_hd__a221o_2
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11956_ _11584_/A _11952_/X _11955_/X vssd1 vssd1 vccd1 vccd1 _11956_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_opt_4_0_wb_clk_i _22899_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_4_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_217_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17463_ _22642_/Q _16297_/X _17465_/S vssd1 vssd1 vccd1 vccd1 _17464_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14675_ _14675_/A _20148_/A vssd1 vssd1 vccd1 vccd1 _14676_/B sky130_fd_sc_hd__nand2_4
X_11887_ _13522_/A _13525_/B vssd1 vssd1 vccd1 vccd1 _13382_/B sky130_fd_sc_hd__or2_1
XFILLER_199_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19202_ _19201_/X _23280_/Q _19211_/S vssd1 vssd1 vccd1 vccd1 _19203_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_338_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16414_ _15422_/X _22369_/Q _16418_/S vssd1 vssd1 vccd1 vccd1 _16415_/A sky130_fd_sc_hd__mux2_1
X_13626_ _21708_/A _13587_/A _15391_/A _13593_/A vssd1 vssd1 vccd1 vccd1 _13956_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_349_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17394_ _17394_/A vssd1 vssd1 vccd1 vccd1 _17394_/Y sky130_fd_sc_hd__inv_2
XFILLER_319_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19133_ _23255_/Q _18830_/X _19135_/S vssd1 vssd1 vccd1 vccd1 _19134_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16345_ _16345_/A vssd1 vssd1 vccd1 vccd1 _22339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_347_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13557_ _13647_/A _16191_/B _16131_/A _13556_/Y _14220_/A vssd1 vssd1 vccd1 vccd1
+ _13686_/B sky130_fd_sc_hd__a311oi_2
XFILLER_346_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_346_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19064_ _19075_/A vssd1 vssd1 vccd1 vccd1 _19073_/S sky130_fd_sc_hd__buf_2
XFILLER_158_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12508_ _11659_/A _12507_/X _11678_/A vssd1 vssd1 vccd1 vccd1 _12508_/X sky130_fd_sc_hd__o21a_1
XFILLER_335_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_334_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_307_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16276_ _22314_/Q _16275_/X _16285_/S vssd1 vssd1 vccd1 vccd1 _16277_/A sky130_fd_sc_hd__mux2_1
X_13488_ _13562_/A vssd1 vssd1 vccd1 vccd1 _13647_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_185_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18015_ _18096_/A vssd1 vssd1 vccd1 vccd1 _18051_/A sky130_fd_sc_hd__buf_2
XFILLER_306_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15227_ _15982_/B vssd1 vssd1 vccd1 vccd1 _16028_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_173_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12439_ _12468_/B _12439_/B _12439_/C vssd1 vssd1 vccd1 vccd1 _13710_/A sky130_fd_sc_hd__nor3_4
Xoutput405 _14026_/X vssd1 vssd1 vccd1 vccd1 din0[9] sky130_fd_sc_hd__buf_2
Xoutput416 _22570_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[17] sky130_fd_sc_hd__buf_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput427 _22580_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[27] sky130_fd_sc_hd__buf_2
XFILLER_315_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput438 _22561_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[8] sky130_fd_sc_hd__buf_2
XFILLER_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15158_ _23918_/Q _15159_/B vssd1 vssd1 vccd1 vccd1 _15274_/C sky130_fd_sc_hd__and2_2
Xoutput449 _22885_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[0] sky130_fd_sc_hd__buf_2
XFILLER_5_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14109_ _22885_/Q vssd1 vssd1 vccd1 vccd1 _14121_/D sky130_fd_sc_hd__clkbuf_2
X_19966_ _23604_/Q _23603_/Q _23602_/Q _23601_/Q vssd1 vssd1 vccd1 vccd1 _19971_/C
+ sky130_fd_sc_hd__and4_1
X_15089_ _15252_/A _15088_/X _15089_/S vssd1 vssd1 vccd1 vccd1 _15090_/B sky130_fd_sc_hd__mux2_2
XFILLER_234_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18917_ _18917_/A vssd1 vssd1 vccd1 vccd1 _23159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19897_ _19897_/A vssd1 vssd1 vccd1 vccd1 _23580_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18848_ _18848_/A vssd1 vssd1 vccd1 vccd1 _23132_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18779_ _18779_/A vssd1 vssd1 vccd1 vccd1 _18779_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_283_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20810_ _20810_/A vssd1 vssd1 vccd1 vccd1 _20810_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21790_ _21790_/A _21790_/B vssd1 vssd1 vccd1 vccd1 _21792_/A sky130_fd_sc_hd__nor2_1
XFILLER_70_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20741_ _16003_/A _20732_/X _20740_/Y vssd1 vssd1 vccd1 vccd1 _20742_/C sky130_fd_sc_hd__a21oi_2
XFILLER_224_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23460_ _23578_/CLK _23460_/D vssd1 vssd1 vccd1 vccd1 _23460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_357_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20672_ _20695_/A _20672_/B _20672_/C vssd1 vssd1 vccd1 vccd1 _20672_/X sky130_fd_sc_hd__or3_1
XFILLER_149_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22411_ _23451_/CLK _22411_/D vssd1 vssd1 vccd1 vccd1 _22411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23391_ _23391_/CLK _23391_/D vssd1 vssd1 vccd1 vccd1 _23391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22342_ _23572_/CLK _22342_/D vssd1 vssd1 vccd1 vccd1 _22342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_326_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_325_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_353_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22273_ _23505_/CLK _22273_/D vssd1 vssd1 vccd1 vccd1 _22273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21224_ _21224_/A vssd1 vssd1 vccd1 vccd1 _23886_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21155_ _23866_/Q _21147_/X _21153_/Y _21154_/X _18192_/X vssd1 vssd1 vccd1 vccd1
+ _23866_/D sky130_fd_sc_hd__o221a_1
XFILLER_144_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_320_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20106_ _20106_/A _20112_/D vssd1 vssd1 vccd1 vccd1 _20107_/C sky130_fd_sc_hd__and2_1
XFILLER_291_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21086_ _20583_/B _21085_/B _21301_/D vssd1 vssd1 vccd1 vccd1 _21086_/X sky130_fd_sc_hd__a21o_1
XFILLER_320_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20037_ _20048_/B _20042_/C _20042_/D _18516_/A vssd1 vssd1 vccd1 vccd1 _20037_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_282_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _12091_/A _11809_/X _11348_/A vssd1 vssd1 vccd1 vccd1 _11810_/X sky130_fd_sc_hd__o21a_1
XFILLER_27_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _22375_/Q _22407_/Q _22696_/Q _23063_/Q _11308_/A _11320_/A vssd1 vssd1 vccd1
+ vccd1 _12790_/X sky130_fd_sc_hd__mux4_2
XFILLER_261_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21988_ _21963_/B _21965_/B _21961_/Y vssd1 vssd1 vccd1 vccd1 _21989_/B sky130_fd_sc_hd__a21o_2
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11741_ _11745_/A vssd1 vssd1 vccd1 vccd1 _11741_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939_ _20969_/A vssd1 vssd1 vccd1 vccd1 _20939_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23727_ _23861_/CLK _23727_/D vssd1 vssd1 vccd1 vccd1 _23727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_270_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11672_ _12029_/A vssd1 vssd1 vccd1 vccd1 _12709_/A sky130_fd_sc_hd__buf_4
X_14460_ _20989_/A _20989_/B _20989_/C vssd1 vssd1 vccd1 vccd1 _20986_/A sky130_fd_sc_hd__or3_4
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23658_ _23818_/CLK _23658_/D vssd1 vssd1 vccd1 vccd1 _23658_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13411_ _14176_/A vssd1 vssd1 vccd1 vccd1 _14675_/A sky130_fd_sc_hd__buf_6
X_22609_ _23646_/CLK _22609_/D vssd1 vssd1 vccd1 vccd1 _22609_/Q sky130_fd_sc_hd__dfxtp_1
X_14391_ _16186_/A vssd1 vssd1 vccd1 vccd1 _14896_/A sky130_fd_sc_hd__clkbuf_4
X_23589_ _23592_/CLK _23589_/D vssd1 vssd1 vccd1 vccd1 _23589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_329_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_328_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_344_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16130_ _16097_/A _14632_/B _14671_/X _15995_/A vssd1 vssd1 vccd1 vccd1 _16130_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_13342_ _13342_/A vssd1 vssd1 vccd1 vccd1 _13625_/A sky130_fd_sc_hd__clkinv_4
XFILLER_154_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_294_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_343_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16061_ _22974_/Q _16177_/S vssd1 vssd1 vccd1 vccd1 _16061_/X sky130_fd_sc_hd__or2_1
X_13273_ _13273_/A _13273_/B vssd1 vssd1 vccd1 vccd1 _13273_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12224_ _22784_/Q _22752_/Q _22653_/Q _22720_/Q _12209_/X _12210_/X vssd1 vssd1 vccd1
+ vccd1 _12225_/B sky130_fd_sc_hd__mux4_1
X_15012_ _15456_/A _14774_/A _14767_/X vssd1 vssd1 vccd1 vccd1 _15012_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_142_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19820_ _23546_/Q _19233_/A _19826_/S vssd1 vssd1 vccd1 vccd1 _19821_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12155_ _12148_/X _12150_/X _12152_/X _12154_/X _11683_/X vssd1 vssd1 vccd1 vccd1
+ _12156_/C sky130_fd_sc_hd__a221o_1
XFILLER_2_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_335_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_257_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11106_ _11106_/A vssd1 vssd1 vccd1 vccd1 _15176_/A sky130_fd_sc_hd__buf_6
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_311_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19751_ _19751_/A vssd1 vssd1 vccd1 vccd1 _23515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16963_ _21294_/B _16984_/B vssd1 vssd1 vccd1 vccd1 _16981_/A sky130_fd_sc_hd__or2_1
X_12086_ _11216_/A _12069_/Y _12076_/X _12085_/X vssd1 vssd1 vccd1 vccd1 _13765_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_311_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18702_ _16819_/X _23078_/Q _18708_/S vssd1 vssd1 vccd1 vccd1 _18703_/A sky130_fd_sc_hd__mux2_1
X_15914_ _14898_/A _15903_/X _15912_/X _15913_/X _15003_/A vssd1 vssd1 vccd1 vccd1
+ _15914_/X sky130_fd_sc_hd__o32a_4
X_19682_ _19242_/X _23485_/Q _19682_/S vssd1 vssd1 vccd1 vccd1 _19683_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16894_ _16894_/A vssd1 vssd1 vccd1 vccd1 _22545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_351_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18633_ _18633_/A vssd1 vssd1 vccd1 vccd1 _23047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_280_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15845_ _15833_/X _15299_/B _15835_/X _15844_/Y _14431_/A vssd1 vssd1 vccd1 vccd1
+ _15845_/X sky130_fd_sc_hd__a221o_1
XFILLER_225_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18564_ _16828_/X _23017_/Q _18564_/S vssd1 vssd1 vccd1 vccd1 _18565_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ _14822_/A _15754_/X _15775_/Y _15673_/A vssd1 vssd1 vccd1 vccd1 _15776_/X
+ sky130_fd_sc_hd__a211o_1
X_12988_ _12988_/A _12988_/B vssd1 vssd1 vccd1 vccd1 _12989_/B sky130_fd_sc_hd__nor2_8
XFILLER_224_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17515_ _17515_/A vssd1 vssd1 vccd1 vccd1 _22664_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14727_ _14897_/A vssd1 vssd1 vccd1 vccd1 _14727_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18495_ _18521_/A vssd1 vssd1 vccd1 vccd1 _18505_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_11939_ _11939_/A _11939_/B vssd1 vssd1 vccd1 vccd1 _13528_/B sky130_fd_sc_hd__nor2_1
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17446_ _22634_/Q _16271_/X _17454_/S vssd1 vssd1 vccd1 vccd1 _17447_/A sky130_fd_sc_hd__mux2_1
X_14658_ _14656_/X _14657_/X _14845_/S vssd1 vssd1 vccd1 vccd1 _14658_/X sky130_fd_sc_hd__mux2_1
XFILLER_296_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13609_ _21846_/A _13603_/X _13608_/Y _13451_/A vssd1 vssd1 vccd1 vccd1 _13966_/A
+ sky130_fd_sc_hd__o22a_2
X_17377_ _17377_/A vssd1 vssd1 vccd1 vccd1 _22608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_308_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14589_ _15903_/B vssd1 vssd1 vccd1 vccd1 _15259_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_220_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19116_ _23247_/Q _18804_/X _19124_/S vssd1 vssd1 vccd1 vccd1 _19117_/A sky130_fd_sc_hd__mux2_1
XFILLER_347_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16328_ _16328_/A vssd1 vssd1 vccd1 vccd1 _22331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19047_ _16854_/X _23217_/Q _19051_/S vssd1 vssd1 vccd1 vccd1 _19048_/A sky130_fd_sc_hd__mux2_1
XFILLER_334_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16259_ _18824_/A vssd1 vssd1 vccd1 vccd1 _16259_/X sky130_fd_sc_hd__buf_2
XFILLER_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_322_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_350_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_303_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_302_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_8 _22193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19949_ _19977_/B _19953_/C vssd1 vssd1 vccd1 vccd1 _19950_/B sky130_fd_sc_hd__and2_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22960_ _22961_/CLK _22960_/D vssd1 vssd1 vccd1 vccd1 _22960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21911_ _21911_/A _21910_/Y vssd1 vssd1 vccd1 vccd1 _21913_/A sky130_fd_sc_hd__or2b_1
XFILLER_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22891_ _23009_/CLK _22891_/D vssd1 vssd1 vccd1 vccd1 _22891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21842_ _21842_/A vssd1 vssd1 vccd1 vccd1 _21842_/X sky130_fd_sc_hd__buf_2
XFILLER_83_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21773_ _21773_/A _21841_/A vssd1 vssd1 vccd1 vccd1 _21773_/X sky130_fd_sc_hd__or2_1
XFILLER_36_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23512_ _23575_/CLK _23512_/D vssd1 vssd1 vccd1 vccd1 _23512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20724_ _20724_/A vssd1 vssd1 vccd1 vccd1 _20724_/X sky130_fd_sc_hd__buf_4
XFILLER_212_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_357_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23443_ _23505_/CLK _23443_/D vssd1 vssd1 vccd1 vccd1 _23443_/Q sky130_fd_sc_hd__dfxtp_1
X_20655_ _20655_/A _20669_/B vssd1 vssd1 vccd1 vccd1 _20658_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23374_ _23534_/CLK _23374_/D vssd1 vssd1 vccd1 vccd1 _23374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20586_ _20774_/A vssd1 vssd1 vccd1 vccd1 _20895_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_325_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_286_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22325_ _23896_/CLK _22325_/D vssd1 vssd1 vccd1 vccd1 _22325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_307_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22256_ _22257_/B _21196_/X _17390_/X vssd1 vssd1 vccd1 vccd1 _23945_/D sky130_fd_sc_hd__o21a_1
XFILLER_118_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21207_ _14196_/B _21202_/X _21206_/Y _21186_/X vssd1 vssd1 vccd1 vccd1 _23881_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_278_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22187_ _22187_/A _22187_/B vssd1 vssd1 vccd1 vccd1 _22189_/A sky130_fd_sc_hd__nand2_1
XFILLER_279_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_321_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21138_ _21097_/A _20890_/B _21158_/A vssd1 vssd1 vccd1 vccd1 _21168_/A sky130_fd_sc_hd__o21ai_4
XFILLER_120_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_321_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21069_ _20754_/A _21008_/A _21068_/X _21061_/X vssd1 vssd1 vccd1 vccd1 _23842_/D
+ sky130_fd_sc_hd__o211a_1
X_13960_ _21081_/A vssd1 vssd1 vccd1 vccd1 _13960_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_280_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12911_ _12707_/X _12904_/X _12906_/X _12910_/X _11378_/A vssd1 vssd1 vccd1 vccd1
+ _12911_/X sky130_fd_sc_hd__a311o_2
XFILLER_274_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13891_ _13890_/B _15112_/A _13890_/Y vssd1 vssd1 vccd1 vccd1 _15187_/A sky130_fd_sc_hd__a21o_4
XFILLER_235_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15630_ _15630_/A vssd1 vssd1 vccd1 vccd1 _17172_/A sky130_fd_sc_hd__buf_6
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _12842_/A vssd1 vssd1 vccd1 vccd1 _12904_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _14801_/A _15546_/Y _15560_/Y _15436_/X vssd1 vssd1 vccd1 vccd1 _15561_/X
+ sky130_fd_sc_hd__o22a_1
X_12773_ _11218_/A _12763_/X _12772_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _13798_/A
+ sky130_fd_sc_hd__a211oi_4
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17300_ _21076_/A _17299_/X _17317_/S vssd1 vssd1 vccd1 vccd1 _17300_/X sky130_fd_sc_hd__mux2_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14753_/A vssd1 vssd1 vccd1 vccd1 _14513_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _18288_/D vssd1 vssd1 vccd1 vccd1 _18286_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_214_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11724_ _23472_/Q _23568_/Q _22532_/Q _22336_/Q _11574_/A _11696_/X vssd1 vssd1 vccd1
+ vccd1 _11724_/X sky130_fd_sc_hd__mux4_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _14792_/A _14676_/B _15492_/S vssd1 vssd1 vccd1 vccd1 _15492_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17231_/A vssd1 vssd1 vccd1 vccd1 _17231_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_302_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11655_ _12105_/A _11655_/B vssd1 vssd1 vccd1 vccd1 _11655_/X sky130_fd_sc_hd__or2_1
X_14443_ _15440_/A vssd1 vssd1 vccd1 vccd1 _14730_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_317_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_88_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23553_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17162_ _21826_/A vssd1 vssd1 vccd1 vccd1 _17163_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11586_ _22471_/Q _22631_/Q _12042_/S vssd1 vssd1 vccd1 vccd1 _11587_/B sky130_fd_sc_hd__mux2_1
X_14374_ _14647_/A vssd1 vssd1 vccd1 vccd1 _14381_/B sky130_fd_sc_hd__buf_2
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16113_ _15676_/X _21278_/A _16112_/X _15365_/X vssd1 vssd1 vccd1 vccd1 _16113_/X
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23047_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13325_ _13608_/A _13350_/A _12812_/B vssd1 vssd1 vccd1 vccd1 _13330_/B sky130_fd_sc_hd__a21o_1
XFILLER_316_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17093_ input79/X input44/X _17132_/S vssd1 vssd1 vccd1 vccd1 _17093_/X sky130_fd_sc_hd__mux2_8
XFILLER_127_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_316_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_344_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16044_ _15480_/X _13562_/B _15663_/X vssd1 vssd1 vccd1 vccd1 _16044_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_142_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_331_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13256_ _21077_/C _13255_/X _11502_/A vssd1 vssd1 vccd1 vccd1 _13256_/X sky130_fd_sc_hd__a21o_1
XFILLER_136_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_331_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_297_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12207_ _22268_/Q _23084_/Q _23500_/Q _22429_/Q _11920_/A _11815_/A vssd1 vssd1 vccd1
+ vccd1 _12208_/B sky130_fd_sc_hd__mux4_2
XFILLER_9_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13187_ _13187_/A _13240_/A vssd1 vssd1 vccd1 vccd1 _13543_/A sky130_fd_sc_hd__nor2_2
XFILLER_97_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_296_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12138_ _22273_/Q _23089_/Q _23505_/Q _22434_/Q _11745_/X _12020_/A vssd1 vssd1 vccd1
+ vccd1 _12139_/B sky130_fd_sc_hd__mux4_1
X_19803_ _19803_/A vssd1 vssd1 vccd1 vccd1 _23538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_340_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17995_ input5/X input280/X _18005_/S vssd1 vssd1 vccd1 vccd1 _17995_/X sky130_fd_sc_hd__mux2_1
XFILLER_312_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19734_ _19756_/A vssd1 vssd1 vccd1 vccd1 _19743_/S sky130_fd_sc_hd__buf_6
X_16946_ _17648_/C _16945_/Y _16949_/A vssd1 vssd1 vccd1 vccd1 _17022_/B sky130_fd_sc_hd__a21oi_1
X_12069_ _11957_/A _12066_/X _12068_/X vssd1 vssd1 vccd1 vccd1 _12069_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19665_ _19217_/X _23477_/Q _19671_/S vssd1 vssd1 vccd1 vccd1 _19666_/A sky130_fd_sc_hd__mux2_1
XFILLER_265_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16877_ _16876_/X _22540_/Q _16877_/S vssd1 vssd1 vccd1 vccd1 _16878_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18616_ _18616_/A vssd1 vssd1 vccd1 vccd1 _23040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ _23933_/Q _15828_/B vssd1 vssd1 vccd1 vccd1 _15829_/B sky130_fd_sc_hd__nor2_1
X_19596_ _19596_/A vssd1 vssd1 vccd1 vccd1 _23446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_252_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18547_ _20324_/A vssd1 vssd1 vccd1 vccd1 _18547_/X sky130_fd_sc_hd__buf_6
XFILLER_252_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15759_ _23801_/Q _14917_/A _15067_/A vssd1 vssd1 vccd1 vccd1 _15759_/X sky130_fd_sc_hd__a21o_1
XFILLER_205_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18478_ _22987_/Q _18478_/B vssd1 vssd1 vccd1 vccd1 _18478_/Y sky130_fd_sc_hd__nand2_1
XFILLER_205_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_339_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17429_ _17429_/A vssd1 vssd1 vccd1 vccd1 _22626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20440_ _23695_/Q _20448_/B vssd1 vssd1 vccd1 vccd1 _20440_/X sky130_fd_sc_hd__or2_1
XFILLER_197_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_308_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23949__508 vssd1 vssd1 vccd1 vccd1 _23949__508/HI localMemory_wb_error_o sky130_fd_sc_hd__conb_1
XFILLER_308_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_307_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20371_ _20226_/X _22119_/A _20370_/X vssd1 vssd1 vccd1 vccd1 _21173_/A sky130_fd_sc_hd__a21oi_4
XFILLER_277_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22110_ _22110_/A _22110_/B vssd1 vssd1 vccd1 vccd1 _22110_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_307_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23090_ _23440_/CLK _23090_/D vssd1 vssd1 vccd1 vccd1 _23090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_304_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_322_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22041_ _22041_/A _22041_/B _22041_/C _22041_/D vssd1 vssd1 vccd1 vccd1 _22042_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_350_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_304_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22943_ _23649_/CLK _22943_/D vssd1 vssd1 vccd1 vccd1 _22943_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_256_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22874_ _22893_/CLK _22874_/D vssd1 vssd1 vccd1 vccd1 _22874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21825_ _21826_/A _21829_/A vssd1 vssd1 vccd1 vccd1 _21827_/A sky130_fd_sc_hd__nor2_1
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21756_ _21756_/A _21756_/B vssd1 vssd1 vccd1 vccd1 _21758_/A sky130_fd_sc_hd__nor2_1
XPHY_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_297_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20707_ _23737_/Q _20697_/X _20705_/X _20706_/X vssd1 vssd1 vccd1 vccd1 _23737_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_4_11_0_wb_clk_i clkbuf_3_5_1_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_11_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21687_ _15379_/Y _22012_/B _21686_/X vssd1 vssd1 vccd1 vccd1 _21688_/B sky130_fd_sc_hd__a21oi_4
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_357_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11440_ _22484_/Q _22644_/Q _13255_/S vssd1 vssd1 vccd1 vccd1 _11440_/X sky130_fd_sc_hd__mux2_1
X_23426_ _23426_/CLK _23426_/D vssd1 vssd1 vccd1 vccd1 _23426_/Q sky130_fd_sc_hd__dfxtp_1
X_20638_ _23727_/Q _20628_/X _20635_/X _20637_/X vssd1 vssd1 vccd1 vccd1 _23727_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23357_ _23549_/CLK _23357_/D vssd1 vssd1 vccd1 vccd1 _23357_/Q sky130_fd_sc_hd__dfxtp_1
X_11371_ _23428_/Q _23044_/Q _23396_/Q _23364_/Q _11364_/A _11365_/A vssd1 vssd1 vccd1
+ vccd1 _11372_/B sky130_fd_sc_hd__mux4_1
X_20569_ _23718_/Q _20542_/X _20568_/X _20559_/X vssd1 vssd1 vccd1 vccd1 _23718_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_299_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22308_ _23444_/CLK _22308_/D vssd1 vssd1 vccd1 vccd1 _22308_/Q sky130_fd_sc_hd__dfxtp_1
X_13110_ _13273_/A _13110_/B vssd1 vssd1 vccd1 vccd1 _13110_/Y sky130_fd_sc_hd__nand2_1
X_14090_ _22592_/Q _14081_/X _13992_/X _14089_/Y vssd1 vssd1 vccd1 vccd1 _14090_/X
+ sky130_fd_sc_hd__a22o_4
X_23288_ _23354_/CLK _23288_/D vssd1 vssd1 vccd1 vccd1 _23288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_341_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ _13041_/A _13041_/B vssd1 vssd1 vccd1 vccd1 _13041_/Y sky130_fd_sc_hd__nor2_1
XFILLER_313_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22239_ _22210_/X _22213_/B _22211_/A vssd1 vssd1 vccd1 vccd1 _22240_/B sky130_fd_sc_hd__a21oi_1
XFILLER_124_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_310_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16800_ _22517_/Q _16729_/A _16730_/A input33/X vssd1 vssd1 vccd1 vccd1 _16801_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_294_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17780_ _17780_/A vssd1 vssd1 vccd1 vccd1 _22765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_135_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _22977_/CLK sky130_fd_sc_hd__clkbuf_16
X_14992_ _23658_/Q _15985_/B vssd1 vssd1 vccd1 vccd1 _14992_/X sky130_fd_sc_hd__or2_1
XFILLER_87_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16731_ _22497_/Q _16729_/X _16730_/X input11/X vssd1 vssd1 vccd1 vccd1 _16732_/B
+ sky130_fd_sc_hd__o22a_1
X_13943_ _13943_/A _13943_/B vssd1 vssd1 vccd1 vccd1 _15256_/A sky130_fd_sc_hd__xnor2_4
XFILLER_281_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19450_ _19450_/A vssd1 vssd1 vccd1 vccd1 _23381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16662_ _22478_/Q _16284_/X _16662_/S vssd1 vssd1 vccd1 vccd1 _16663_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13874_ _13874_/A _13874_/B _13874_/C vssd1 vssd1 vccd1 vccd1 _13874_/X sky130_fd_sc_hd__and3_1
XFILLER_35_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18401_ _18401_/A _18401_/B _18402_/B vssd1 vssd1 vccd1 vccd1 _22961_/D sky130_fd_sc_hd__nor3_1
XFILLER_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15613_ _16004_/A _15612_/Y _15480_/A vssd1 vssd1 vccd1 vccd1 _15613_/X sky130_fd_sc_hd__o21a_1
X_19381_ _23351_/Q _18830_/X _19383_/S vssd1 vssd1 vccd1 vccd1 _19382_/A sky130_fd_sc_hd__mux2_1
X_12825_ _12825_/A vssd1 vssd1 vccd1 vccd1 _12825_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_234_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16593_ _15975_/X _22447_/Q _16601_/S vssd1 vssd1 vccd1 vccd1 _16594_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18332_ _22936_/Q _22937_/Q _18332_/C vssd1 vssd1 vccd1 vccd1 _18334_/B sky130_fd_sc_hd__and3_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15544_ _13531_/A _15196_/X _15543_/X vssd1 vssd1 vccd1 vccd1 _15544_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12756_ _12756_/A vssd1 vssd1 vccd1 vccd1 _12756_/X sky130_fd_sc_hd__buf_6
XFILLER_187_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18263_ _18263_/A _18263_/B _22916_/Q vssd1 vssd1 vccd1 vccd1 _18264_/C sky130_fd_sc_hd__and3_1
X_11707_ _11723_/A _11704_/X _11706_/X vssd1 vssd1 vccd1 vccd1 _11707_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15475_ _15474_/X _22274_/Q _15524_/S vssd1 vssd1 vccd1 vccd1 _15476_/A sky130_fd_sc_hd__mux2_1
X_12687_ _12687_/A vssd1 vssd1 vccd1 vccd1 _12687_/X sky130_fd_sc_hd__buf_2
XFILLER_348_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17214_ _21975_/A _17213_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17214_/X sky130_fd_sc_hd__mux2_1
X_14426_ _14451_/B _14465_/B vssd1 vssd1 vccd1 vccd1 _14434_/B sky130_fd_sc_hd__or2_1
X_18194_ _18188_/A _18188_/B _18178_/X _18195_/A vssd1 vssd1 vccd1 vccd1 _18194_/X
+ sky130_fd_sc_hd__a31o_1
X_11638_ _22278_/Q _23094_/Q _23510_/Q _22439_/Q _11637_/X _12777_/A vssd1 vssd1 vccd1
+ vccd1 _11639_/B sky130_fd_sc_hd__mux4_2
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17145_ _17145_/A _17145_/B vssd1 vssd1 vccd1 vccd1 _17220_/B sky130_fd_sc_hd__and2_1
XFILLER_129_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14357_ _14762_/A _13362_/B _14356_/Y _14351_/S vssd1 vssd1 vccd1 vccd1 _14357_/X
+ sky130_fd_sc_hd__a211o_1
X_11569_ _23222_/Q _23190_/Q _23158_/Q _23126_/Q _12820_/S _12749_/A vssd1 vssd1 vccd1
+ vccd1 _11570_/B sky130_fd_sc_hd__mux4_2
XFILLER_116_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13308_ _13311_/A vssd1 vssd1 vccd1 vccd1 _13555_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_289_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17076_ _14546_/X _17074_/X _17116_/S vssd1 vssd1 vccd1 vccd1 _17076_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14288_ _14288_/A vssd1 vssd1 vccd1 vccd1 _14330_/S sky130_fd_sc_hd__buf_2
XFILLER_332_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_304_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16027_ _14730_/X _16020_/X _16026_/Y _15150_/X vssd1 vssd1 vccd1 vccd1 _16028_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_304_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13239_ _13561_/A _13402_/A _13239_/C vssd1 vssd1 vccd1 vccd1 _13239_/X sky130_fd_sc_hd__and3b_1
XFILLER_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_301_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_300_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater502 _12800_/Y vssd1 vssd1 vccd1 vccd1 _21871_/A sky130_fd_sc_hd__buf_6
X_17978_ _22836_/Q _17972_/X _17896_/X _17977_/X _17966_/X vssd1 vssd1 vccd1 vccd1
+ _17978_/X sky130_fd_sc_hd__a221o_1
XFILLER_242_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16929_ _16929_/A vssd1 vssd1 vccd1 vccd1 _17244_/B sky130_fd_sc_hd__clkbuf_2
X_19717_ _19188_/X _23500_/Q _19721_/S vssd1 vssd1 vccd1 vccd1 _19718_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_348_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19648_ _19648_/A vssd1 vssd1 vccd1 vccd1 _23469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_253_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19579_ _19625_/S vssd1 vssd1 vccd1 vccd1 _19588_/S sky130_fd_sc_hd__buf_4
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21610_ _21377_/X _21589_/X _21595_/Y _21609_/Y vssd1 vssd1 vccd1 vccd1 _21610_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22590_ _22977_/CLK _22590_/D vssd1 vssd1 vccd1 vccd1 _22590_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_178_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21541_ _21542_/C vssd1 vssd1 vccd1 vccd1 _21548_/A sky130_fd_sc_hd__inv_2
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21472_ _21472_/A _21472_/B _21472_/C vssd1 vssd1 vccd1 vccd1 _21472_/X sky130_fd_sc_hd__or3_1
XFILLER_193_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_348_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23211_ _23531_/CLK _23211_/D vssd1 vssd1 vccd1 vccd1 _23211_/Q sky130_fd_sc_hd__dfxtp_1
X_20423_ _20579_/A _20408_/X _20422_/X _20420_/X vssd1 vssd1 vccd1 vccd1 _23688_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_335_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23142_ _23526_/CLK _23142_/D vssd1 vssd1 vccd1 vccd1 _23142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20354_ _15914_/X _20169_/X _20355_/B vssd1 vssd1 vccd1 vccd1 _20354_/X sky130_fd_sc_hd__a21o_1
XFILLER_323_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_351_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23073_ _23073_/CLK _23073_/D vssd1 vssd1 vccd1 vccd1 _23073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_350_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_289_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20285_ _20324_/A vssd1 vssd1 vccd1 vccd1 _20285_/X sky130_fd_sc_hd__clkbuf_2
XTAP_6206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22024_ _22024_/A _22024_/B vssd1 vssd1 vccd1 vccd1 _22025_/B sky130_fd_sc_hd__xnor2_1
XFILLER_304_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_288_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22926_ _22929_/CLK _22926_/D vssd1 vssd1 vccd1 vccd1 _22926_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_216_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_290_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_1_wb_clk_i clkbuf_2_1_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22857_ _22908_/CLK _22857_/D vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dfxtp_1
XFILLER_204_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _13340_/A _12611_/B vssd1 vssd1 vccd1 vccd1 _13942_/A sky130_fd_sc_hd__and2_2
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21808_ _21809_/A _21809_/B vssd1 vssd1 vccd1 vccd1 _21876_/A sky130_fd_sc_hd__and2_1
XFILLER_169_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _12916_/B _13604_/A _13633_/A _13493_/Y vssd1 vssd1 vccd1 vccd1 _13601_/B
+ sky130_fd_sc_hd__o31ai_4
X_22788_ _23578_/CLK _22788_/D vssd1 vssd1 vccd1 vccd1 _22788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12541_ _12523_/A _12536_/Y _12538_/Y _12540_/Y vssd1 vssd1 vccd1 vccd1 _12541_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_358_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21739_ _21739_/A _21739_/B vssd1 vssd1 vccd1 vccd1 _21740_/B sky130_fd_sc_hd__nand2_1
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15260_ _23598_/Q _14450_/X _14455_/X _23630_/Q vssd1 vssd1 vccd1 vccd1 _15260_/X
+ sky130_fd_sc_hd__o22a_2
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12472_ _13505_/A vssd1 vssd1 vccd1 vccd1 _14292_/A sky130_fd_sc_hd__buf_6
XFILLER_138_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_327_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14211_ _14211_/A _14211_/B _14211_/C vssd1 vssd1 vccd1 vccd1 _14980_/A sky130_fd_sc_hd__and3_4
X_23409_ _23409_/CLK _23409_/D vssd1 vssd1 vccd1 vccd1 _23409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11423_ _23331_/Q _23299_/Q _23267_/Q _23555_/Q _11157_/X _11418_/X vssd1 vssd1 vccd1
+ vccd1 _11424_/B sky130_fd_sc_hd__mux4_2
X_15191_ _14243_/Y _15181_/X _15183_/X _15190_/Y vssd1 vssd1 vccd1 vccd1 _21225_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_138_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_326_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14142_ _14148_/A _14148_/B _14148_/C _13662_/B vssd1 vssd1 vccd1 vccd1 _14211_/C
+ sky130_fd_sc_hd__nor4b_4
X_11354_ _13291_/A _11341_/X _11343_/X _15671_/A vssd1 vssd1 vccd1 vccd1 _11354_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_327_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_299_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_314_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11285_ _11285_/A vssd1 vssd1 vccd1 vccd1 _12707_/A sky130_fd_sc_hd__buf_2
X_14073_ _22809_/Q _14027_/X _14072_/X vssd1 vssd1 vccd1 vccd1 _14073_/X sky130_fd_sc_hd__a21o_4
XFILLER_180_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18950_ _18950_/A vssd1 vssd1 vccd1 vccd1 _23173_/D sky130_fd_sc_hd__clkbuf_1
X_17901_ _22813_/Q _17891_/X _17900_/X _17657_/X vssd1 vssd1 vccd1 vccd1 _22813_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_279_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13024_ _13493_/A _13019_/Y _13023_/X vssd1 vssd1 vccd1 vccd1 _13323_/B sky130_fd_sc_hd__a21boi_1
X_18881_ _23143_/Q _18779_/X _18885_/S vssd1 vssd1 vccd1 vccd1 _18882_/A sky130_fd_sc_hd__mux2_1
XTAP_6740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17832_ _17832_/A vssd1 vssd1 vccd1 vccd1 _22788_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17763_ _22758_/Q _17588_/X _17765_/S vssd1 vssd1 vccd1 vccd1 _17764_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14975_ _23915_/Q vssd1 vssd1 vccd1 vccd1 _21431_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19502_ _19502_/A vssd1 vssd1 vccd1 vccd1 _23404_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16714_ _16723_/A _16714_/B vssd1 vssd1 vccd1 vccd1 _16715_/A sky130_fd_sc_hd__or2_1
XFILLER_281_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13926_ _13933_/A _14091_/A vssd1 vssd1 vccd1 vccd1 _13926_/Y sky130_fd_sc_hd__nor2_2
X_17694_ _17694_/A vssd1 vssd1 vccd1 vccd1 _22727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_402 _13989_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19433_ _23374_/Q _18801_/X _19433_/S vssd1 vssd1 vccd1 vccd1 _19434_/A sky130_fd_sc_hd__mux2_1
X_16645_ _22470_/Q _16259_/X _16651_/S vssd1 vssd1 vccd1 vccd1 _16646_/A sky130_fd_sc_hd__mux2_1
XFILLER_290_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_413 _14033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13857_ _13874_/A _13857_/B _13874_/C vssd1 vssd1 vccd1 vccd1 _13857_/X sky130_fd_sc_hd__and3_1
XFILLER_90_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_424 _14127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_435 _23885_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_446 _23946_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19364_ _23343_/Q _18804_/X _19372_/S vssd1 vssd1 vccd1 vccd1 _19365_/A sky130_fd_sc_hd__mux2_1
X_12808_ _23929_/Q _13296_/B _12801_/X vssd1 vssd1 vccd1 vccd1 _12809_/B sky130_fd_sc_hd__o21a_1
XINSDIODE2_457 _22122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16576_ _16576_/A vssd1 vssd1 vccd1 vccd1 _22439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13788_ _13831_/B vssd1 vssd1 vccd1 vccd1 _13789_/A sky130_fd_sc_hd__dlymetal6s2s_1
XINSDIODE2_468 _15176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_479 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18315_ _18315_/A _18315_/B _18315_/C vssd1 vssd1 vccd1 vccd1 _22931_/D sky130_fd_sc_hd__nor3_1
X_15527_ _21771_/A vssd1 vssd1 vccd1 vccd1 _17149_/A sky130_fd_sc_hd__buf_6
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19295_ _19295_/A vssd1 vssd1 vccd1 vccd1 _23312_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_32_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23578_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12739_ _12739_/A vssd1 vssd1 vccd1 vccd1 _13500_/A sky130_fd_sc_hd__buf_4
XFILLER_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_336_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18246_ _22861_/Q _18242_/X _18244_/X _18245_/X vssd1 vssd1 vccd1 vccd1 _22909_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15458_ _15011_/A _14768_/Y _15456_/Y _15457_/Y vssd1 vssd1 vccd1 vccd1 _15458_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14409_ _21550_/A _14550_/B _14433_/S vssd1 vssd1 vccd1 vccd1 _14416_/A sky130_fd_sc_hd__mux2_1
X_18177_ _18118_/X _18126_/S _18176_/Y vssd1 vssd1 vccd1 vccd1 _22890_/D sky130_fd_sc_hd__o21a_1
XFILLER_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ _13625_/A _14792_/A _15388_/Y _12160_/A vssd1 vssd1 vccd1 vccd1 _15389_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_345_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_317_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17128_ _17073_/A _17126_/X _17107_/X _17127_/X vssd1 vssd1 vccd1 vccd1 _17128_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_117_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_289_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_332_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_305_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_289_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_289_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17059_ _22559_/Q _17038_/X _17028_/X _17058_/X vssd1 vssd1 vccd1 vccd1 _22559_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_131_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20070_ _20079_/B _20071_/C _20069_/Y vssd1 vssd1 vccd1 vccd1 _23631_/D sky130_fd_sc_hd__o21a_1
XFILLER_332_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_300_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20972_ _23806_/Q _20969_/X _20971_/X _20964_/X vssd1 vssd1 vccd1 vccd1 _23806_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23760_ _23878_/CLK _23760_/D vssd1 vssd1 vccd1 vccd1 _23760_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_93_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22711_ _23851_/CLK _22711_/D vssd1 vssd1 vccd1 vccd1 _22711_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_281_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23691_ _23696_/CLK _23691_/D vssd1 vssd1 vccd1 vccd1 _23691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22642_ _23880_/CLK _22642_/D vssd1 vssd1 vccd1 vccd1 _22642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_322_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_322_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22573_ _23643_/CLK _22573_/D vssd1 vssd1 vccd1 vccd1 _22573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_328_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21524_ _21521_/Y _21522_/X _16016_/A _21549_/A vssd1 vssd1 vccd1 vccd1 _21542_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_327_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21455_ _21813_/A _21454_/X _21381_/X _23786_/Q vssd1 vssd1 vccd1 vccd1 _21455_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_135_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20406_ _20409_/A _20986_/B vssd1 vssd1 vccd1 vccd1 _20467_/A sky130_fd_sc_hd__or2_1
XFILLER_308_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21386_ _21386_/A _21443_/A vssd1 vssd1 vccd1 vccd1 _21386_/X sky130_fd_sc_hd__or2_1
XFILLER_335_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_323_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23125_ _23543_/CLK _23125_/D vssd1 vssd1 vccd1 vccd1 _23125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20337_ _20302_/X _20335_/X _20336_/Y _21979_/A _20307_/X vssd1 vssd1 vccd1 vccd1
+ _20708_/A sky130_fd_sc_hd__a32o_4
XFILLER_311_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_296_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23056_ _23058_/CLK _23056_/D vssd1 vssd1 vccd1 vccd1 _23056_/Q sky130_fd_sc_hd__dfxtp_1
X_11070_ _14132_/D vssd1 vssd1 vccd1 vccd1 _21335_/A sky130_fd_sc_hd__clkbuf_4
XTAP_6025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20268_ _21708_/B vssd1 vssd1 vccd1 vccd1 _20268_/Y sky130_fd_sc_hd__inv_2
XTAP_6036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput102 dout0[63] vssd1 vssd1 vccd1 vccd1 input102/X sky130_fd_sc_hd__clkbuf_1
X_22007_ _22098_/A vssd1 vssd1 vccd1 vccd1 _22100_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_6069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput113 dout1[15] vssd1 vssd1 vccd1 vccd1 input113/X sky130_fd_sc_hd__clkbuf_1
XTAP_5324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput124 dout1[25] vssd1 vssd1 vccd1 vccd1 input124/X sky130_fd_sc_hd__clkbuf_1
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20199_ _20236_/A _20199_/B vssd1 vssd1 vccd1 vccd1 _20199_/Y sky130_fd_sc_hd__nand2_1
Xinput135 dout1[35] vssd1 vssd1 vccd1 vccd1 input135/X sky130_fd_sc_hd__buf_2
XTAP_5346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput146 dout1[45] vssd1 vssd1 vccd1 vccd1 input146/X sky130_fd_sc_hd__buf_2
XTAP_5357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput157 dout1[55] vssd1 vssd1 vccd1 vccd1 input157/X sky130_fd_sc_hd__buf_2
XFILLER_276_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput168 dout1[7] vssd1 vssd1 vccd1 vccd1 input168/X sky130_fd_sc_hd__clkbuf_2
XTAP_5379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_313_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput179 irq[2] vssd1 vssd1 vccd1 vccd1 _20524_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_292_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _14760_/A vssd1 vssd1 vccd1 vccd1 _14761_/A sky130_fd_sc_hd__clkbuf_4
X_11972_ _11972_/A vssd1 vssd1 vccd1 vccd1 _11972_/X sky130_fd_sc_hd__buf_4
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13711_ _13721_/B _13711_/B vssd1 vssd1 vccd1 vccd1 _13712_/B sky130_fd_sc_hd__nor2_4
X_22909_ _23008_/CLK _22909_/D vssd1 vssd1 vccd1 vccd1 _22909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _14682_/X _14688_/X _14690_/X vssd1 vssd1 vccd1 vccd1 _14691_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23889_ _23907_/CLK _23889_/D vssd1 vssd1 vccd1 vccd1 _23889_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_260_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16430_ _16430_/A vssd1 vssd1 vccd1 vccd1 _22376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13642_ _23922_/Q vssd1 vssd1 vccd1 vccd1 _21673_/A sky130_fd_sc_hd__buf_4
XFILLER_60_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _16361_/A vssd1 vssd1 vccd1 vccd1 _22346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13573_ _13573_/A _13573_/B vssd1 vssd1 vccd1 vccd1 _13574_/B sky130_fd_sc_hd__or2_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18100_ _22870_/Q _18097_/X _18098_/X _23003_/Q _18099_/X vssd1 vssd1 vccd1 vccd1
+ _18100_/X sky130_fd_sc_hd__a221o_1
XFILLER_158_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_297_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15312_ _14898_/X _15299_/X _15309_/X _15311_/X _14937_/X vssd1 vssd1 vccd1 vccd1
+ _15312_/X sky130_fd_sc_hd__o32a_4
XFILLER_40_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_347_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19080_ _16902_/X _23232_/Q _19084_/S vssd1 vssd1 vccd1 vccd1 _19081_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _22261_/Q _23077_/Q _23493_/Q _22422_/Q _11146_/A _11701_/A vssd1 vssd1 vccd1
+ vccd1 _12525_/B sky130_fd_sc_hd__mux4_1
X_16292_ _22319_/Q _16291_/X _16301_/S vssd1 vssd1 vccd1 vccd1 _16293_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_347_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_318_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18031_ hold3/A _18017_/X _18020_/X _22981_/Q _18023_/X vssd1 vssd1 vccd1 vccd1 _18031_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_201_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15243_ _15243_/A _15432_/B vssd1 vssd1 vccd1 vccd1 _15243_/Y sky130_fd_sc_hd__nand2_2
XFILLER_334_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12455_ _22455_/Q _22615_/Q _12457_/S vssd1 vssd1 vccd1 vccd1 _12456_/B sky130_fd_sc_hd__mux2_1
XFILLER_327_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_315_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11406_ _12135_/A vssd1 vssd1 vccd1 vccd1 _12661_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15174_ _15172_/Y _15173_/X _15080_/A vssd1 vssd1 vccd1 vccd1 _15174_/X sky130_fd_sc_hd__a21bo_1
XFILLER_314_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12386_ _22780_/Q _22748_/Q _22649_/Q _22716_/Q _12215_/X _12216_/X vssd1 vssd1 vccd1
+ vccd1 _12387_/B sky130_fd_sc_hd__mux4_1
XFILLER_314_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14125_ _18163_/B _18187_/B vssd1 vssd1 vccd1 vccd1 _14125_/Y sky130_fd_sc_hd__nor2_2
XFILLER_299_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11337_ _13131_/A vssd1 vssd1 vccd1 vccd1 _13287_/A sky130_fd_sc_hd__buf_4
XFILLER_181_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19982_ _23607_/Q _20005_/C _19981_/Y vssd1 vssd1 vccd1 vccd1 _23607_/D sky130_fd_sc_hd__o21a_1
XFILLER_314_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_341_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_287_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_341_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_330_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_354_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18933_ _18933_/A vssd1 vssd1 vccd1 vccd1 _23166_/D sky130_fd_sc_hd__clkbuf_1
X_14056_ _14064_/A _14066_/B _14056_/C vssd1 vssd1 vccd1 vccd1 _14056_/X sky130_fd_sc_hd__or3_1
XFILLER_98_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11268_ _11398_/A _12087_/A vssd1 vssd1 vccd1 vccd1 _11269_/S sky130_fd_sc_hd__nor2_1
XTAP_7271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13007_ _22476_/Q _22636_/Q _22315_/Q _23451_/Q _11532_/A _11533_/A vssd1 vssd1 vccd1
+ vccd1 _13007_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18864_ _18864_/A vssd1 vssd1 vccd1 vccd1 _23137_/D sky130_fd_sc_hd__clkbuf_1
X_11199_ _21077_/C _11199_/B vssd1 vssd1 vccd1 vccd1 _11199_/Y sky130_fd_sc_hd__nand2_1
XTAP_6570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17815_ _22781_/Q _17559_/X _17815_/S vssd1 vssd1 vccd1 vccd1 _17816_/A sky130_fd_sc_hd__mux2_1
X_18795_ _18795_/A vssd1 vssd1 vccd1 vccd1 _18795_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17746_ _22750_/Q _17562_/X _17754_/S vssd1 vssd1 vccd1 vccd1 _17747_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14958_ _15010_/A _14958_/B _14958_/C vssd1 vssd1 vccd1 vccd1 _14958_/X sky130_fd_sc_hd__and3_1
XFILLER_130_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13909_ _23916_/Q vssd1 vssd1 vccd1 vccd1 _15037_/A sky130_fd_sc_hd__buf_2
XFILLER_291_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17677_ _17677_/A vssd1 vssd1 vccd1 vccd1 _22719_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_210 _15595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14889_ _14819_/X _14883_/X _14888_/X vssd1 vssd1 vccd1 vccd1 _14889_/X sky130_fd_sc_hd__a21o_1
XINSDIODE2_221 _14925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_232 _15155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19416_ _23366_/Q _18776_/X _19422_/S vssd1 vssd1 vccd1 vccd1 _19417_/A sky130_fd_sc_hd__mux2_1
X_16628_ _16628_/A vssd1 vssd1 vccd1 vccd1 _22462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_243 _15329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_254 _15560_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_265 _15651_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_276 _21916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_287 _15959_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16559_ _16605_/S vssd1 vssd1 vccd1 vccd1 _16568_/S sky130_fd_sc_hd__buf_4
X_19347_ _19347_/A vssd1 vssd1 vccd1 vccd1 _23335_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_298 _15990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19278_ _19178_/X _23305_/Q _19278_/S vssd1 vssd1 vccd1 vccd1 _19279_/A sky130_fd_sc_hd__mux2_1
XFILLER_337_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18229_ _18242_/A vssd1 vssd1 vccd1 vccd1 _18229_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_324_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21240_ _21240_/A _21240_/B vssd1 vssd1 vccd1 vccd1 _21240_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_333_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21171_ _20731_/A _21158_/X _21142_/A _20509_/C _21161_/X vssd1 vssd1 vccd1 vccd1
+ _21171_/X sky130_fd_sc_hd__a221o_1
XFILLER_171_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20122_ _23647_/Q _20122_/B vssd1 vssd1 vccd1 vccd1 _20124_/B sky130_fd_sc_hd__nor2_1
XFILLER_264_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20053_ _20066_/B _20066_/C _20052_/Y vssd1 vssd1 vccd1 vccd1 _23627_/D sky130_fd_sc_hd__o21a_1
XFILLER_98_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_301_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23812_ _23866_/CLK _23812_/D vssd1 vssd1 vccd1 vccd1 _23812_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23743_ _23915_/CLK _23743_/D vssd1 vssd1 vccd1 vccd1 _23743_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20955_ _21949_/A _20950_/X _20705_/B _20954_/X vssd1 vssd1 vccd1 vccd1 _20955_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_289_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23674_ _23684_/CLK _23674_/D vssd1 vssd1 vccd1 vccd1 _23674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_289_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20886_ _21215_/A _20886_/B vssd1 vssd1 vccd1 vccd1 _20887_/A sky130_fd_sc_hd__and2_1
XFILLER_214_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22625_ _23440_/CLK _22625_/D vssd1 vssd1 vccd1 vccd1 _22625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22556_ _22968_/CLK _22556_/D vssd1 vssd1 vccd1 vccd1 _22556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_356_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_356_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21507_ _13923_/B _21479_/X _21489_/Y _21506_/X _21175_/X vssd1 vssd1 vccd1 vccd1
+ _23917_/D sky130_fd_sc_hd__o221a_1
X_22487_ _23841_/CLK _22487_/D vssd1 vssd1 vccd1 vccd1 _22487_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_108_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_309_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12240_ _23211_/Q _23179_/Q _23147_/Q _23115_/Q _11414_/A _11703_/A vssd1 vssd1 vccd1
+ vccd1 _12241_/B sky130_fd_sc_hd__mux4_1
XFILLER_147_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21438_ _21398_/X _21435_/Y _21437_/Y _21408_/X vssd1 vssd1 vccd1 vccd1 _21438_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_135_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_352_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12171_ _12171_/A _12171_/B vssd1 vssd1 vccd1 vccd1 _12171_/Y sky130_fd_sc_hd__nand2_2
X_21369_ _23815_/Q _23749_/Q vssd1 vssd1 vccd1 vccd1 _21373_/A sky130_fd_sc_hd__nand2_1
XFILLER_150_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_351_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_312_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11122_ _12134_/A vssd1 vssd1 vccd1 vccd1 _12660_/A sky130_fd_sc_hd__buf_6
X_23108_ _23578_/CLK _23108_/D vssd1 vssd1 vccd1 vccd1 _23108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15930_ _15929_/X _15478_/X _16195_/S vssd1 vssd1 vccd1 vccd1 _15930_/Y sky130_fd_sc_hd__a21oi_1
X_23039_ _23423_/CLK _23039_/D vssd1 vssd1 vccd1 vccd1 _23039_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15861_ _19236_/A vssd1 vssd1 vccd1 vccd1 _15861_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _17600_/A vssd1 vssd1 vccd1 vccd1 _22694_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14812_ _14811_/X _22263_/Q _14985_/S vssd1 vssd1 vccd1 vccd1 _14813_/A sky130_fd_sc_hd__mux2_1
X_18580_ _16851_/X _23024_/Q _18586_/S vssd1 vssd1 vccd1 vccd1 _18581_/A sky130_fd_sc_hd__mux2_1
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15792_ _15828_/B _15792_/B vssd1 vssd1 vccd1 vccd1 _15793_/B sky130_fd_sc_hd__or2_1
XFILLER_224_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _17531_/A vssd1 vssd1 vccd1 vccd1 _22671_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14743_ _23751_/Q _15595_/A _15596_/A _14741_/X _14742_/X vssd1 vssd1 vccd1 vccd1
+ _14743_/X sky130_fd_sc_hd__a221o_1
X_11955_ _12671_/A _11954_/X _11961_/A vssd1 vssd1 vccd1 vccd1 _11955_/X sky130_fd_sc_hd__a21o_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17462_ _17462_/A vssd1 vssd1 vccd1 vccd1 _22641_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14674_ _14674_/A vssd1 vssd1 vccd1 vccd1 _14674_/X sky130_fd_sc_hd__clkbuf_4
X_11886_ _13523_/B vssd1 vssd1 vccd1 vccd1 _13525_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_260_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19201_ _19201_/A vssd1 vssd1 vccd1 vccd1 _19201_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16413_ _16413_/A vssd1 vssd1 vccd1 vccd1 _22368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13625_ _13625_/A _13625_/B vssd1 vssd1 vccd1 vccd1 _15391_/A sky130_fd_sc_hd__xnor2_4
X_17393_ _22613_/Q _16927_/B _16927_/A vssd1 vssd1 vccd1 vccd1 _17396_/B sky130_fd_sc_hd__o21ai_1
XFILLER_60_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_349_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19132_ _19132_/A vssd1 vssd1 vccd1 vccd1 _23254_/D sky130_fd_sc_hd__clkbuf_1
X_16344_ _15523_/X _22339_/Q _16344_/S vssd1 vssd1 vccd1 vccd1 _16345_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_319_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13556_ _13562_/A _23942_/Q _23941_/Q vssd1 vssd1 vccd1 vccd1 _13556_/Y sky130_fd_sc_hd__nor3_1
XFILLER_346_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_347_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19063_ _19063_/A vssd1 vssd1 vccd1 vccd1 _23224_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_307_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12507_ _23397_/Q _23013_/Q _23365_/Q _23333_/Q _12501_/X _12502_/X vssd1 vssd1 vccd1
+ vccd1 _12507_/X sky130_fd_sc_hd__mux4_1
X_16275_ _18840_/A vssd1 vssd1 vccd1 vccd1 _16275_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_346_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13487_ _13570_/A vssd1 vssd1 vccd1 vccd1 _13562_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18014_ _18198_/B _18021_/B vssd1 vssd1 vccd1 vccd1 _18096_/A sky130_fd_sc_hd__nor2_4
X_15226_ _15501_/B vssd1 vssd1 vccd1 vccd1 _15982_/B sky130_fd_sc_hd__buf_2
XFILLER_218_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12438_ _12431_/Y _12433_/Y _12435_/Y _12437_/Y _11241_/A vssd1 vssd1 vccd1 vccd1
+ _12439_/C sky130_fd_sc_hd__o221a_1
XFILLER_126_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_315_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput406 _14127_/X vssd1 vssd1 vccd1 vccd1 jtag_tdo sky130_fd_sc_hd__buf_2
XFILLER_315_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput417 _22571_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[18] sky130_fd_sc_hd__buf_2
Xoutput428 _22581_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[28] sky130_fd_sc_hd__buf_2
XFILLER_160_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15157_ _14822_/X _15121_/X _15156_/X _14882_/X vssd1 vssd1 vccd1 vccd1 _15157_/X
+ sky130_fd_sc_hd__a22o_1
Xoutput439 _22562_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[9] sky130_fd_sc_hd__buf_2
X_12369_ _23889_/Q vssd1 vssd1 vccd1 vccd1 _12370_/A sky130_fd_sc_hd__inv_2
XFILLER_114_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_315_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14108_ _22889_/Q _22886_/Q vssd1 vssd1 vccd1 vccd1 _14110_/B sky130_fd_sc_hd__or2_1
XFILLER_287_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19965_ _19976_/B _19960_/B _23604_/Q vssd1 vssd1 vccd1 vccd1 _19970_/B sky130_fd_sc_hd__a21oi_1
X_15088_ _15085_/X _15087_/X _15088_/S vssd1 vssd1 vccd1 vccd1 _15088_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18916_ _23159_/Q _18830_/X _18918_/S vssd1 vssd1 vccd1 vccd1 _18917_/A sky130_fd_sc_hd__mux2_1
X_14039_ _14046_/A _14052_/B _14039_/C vssd1 vssd1 vccd1 vccd1 _14039_/X sky130_fd_sc_hd__or3_1
XTAP_7090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19896_ _16281_/X _23580_/Q _19898_/S vssd1 vssd1 vccd1 vccd1 _19897_/A sky130_fd_sc_hd__mux2_1
XFILLER_268_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18847_ _23132_/Q _18846_/X _18850_/S vssd1 vssd1 vccd1 vccd1 _18848_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18778_ _18778_/A vssd1 vssd1 vccd1 vccd1 _23110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17729_ _17729_/A vssd1 vssd1 vccd1 vccd1 _22743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_282_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20740_ _21078_/A _20724_/X _20733_/X vssd1 vssd1 vccd1 vccd1 _20740_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_251_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20671_ _21790_/A _20648_/X _20670_/Y vssd1 vssd1 vccd1 vccd1 _20672_/C sky130_fd_sc_hd__a21oi_1
XFILLER_211_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22410_ _23068_/CLK _22410_/D vssd1 vssd1 vccd1 vccd1 _22410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23390_ _23547_/CLK _23390_/D vssd1 vssd1 vccd1 vccd1 _23390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_337_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22341_ _23573_/CLK _22341_/D vssd1 vssd1 vccd1 vccd1 _22341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_352_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22272_ _23504_/CLK _22272_/D vssd1 vssd1 vccd1 vccd1 _22272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_353_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21223_ _21258_/A _21223_/B vssd1 vssd1 vccd1 vccd1 _21224_/A sky130_fd_sc_hd__and2_1
XFILLER_88_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_321_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_306_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21154_ _21083_/X _20515_/B _21150_/X vssd1 vssd1 vccd1 vccd1 _21154_/X sky130_fd_sc_hd__a21o_1
XFILLER_105_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20105_ _23642_/Q _23641_/Q vssd1 vssd1 vccd1 vccd1 _20112_/D sky130_fd_sc_hd__and2_1
XFILLER_59_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_320_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21085_ _21085_/A _21085_/B vssd1 vssd1 vccd1 vccd1 _21085_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20036_ _23623_/Q vssd1 vssd1 vccd1 vccd1 _20048_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_291_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_328_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21987_ _21987_/A _22041_/C vssd1 vssd1 vccd1 vccd1 _21989_/A sky130_fd_sc_hd__xnor2_4
XFILLER_57_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11740_ _12144_/A vssd1 vssd1 vccd1 vccd1 _12780_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_199_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23726_ _23755_/CLK _23726_/D vssd1 vssd1 vccd1 vccd1 _23726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20938_ _23795_/Q _20925_/X _20937_/X _20934_/X vssd1 vssd1 vccd1 vccd1 _23795_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11671_ _12842_/A _11670_/X _11631_/A vssd1 vssd1 vccd1 vccd1 _11671_/X sky130_fd_sc_hd__o21a_1
X_23657_ _23818_/CLK _23657_/D vssd1 vssd1 vccd1 vccd1 _23657_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_144_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20869_ _20736_/B _20864_/X _20865_/X _23774_/Q vssd1 vssd1 vccd1 vccd1 _20870_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13410_ _13410_/A _13410_/B _13410_/C _13410_/D vssd1 vssd1 vccd1 vccd1 _13410_/Y
+ sky130_fd_sc_hd__nor4_1
X_22608_ _23646_/CLK _22608_/D vssd1 vssd1 vccd1 vccd1 _22608_/Q sky130_fd_sc_hd__dfxtp_1
X_14390_ _13470_/X _13427_/A _13427_/B _14389_/X vssd1 vssd1 vccd1 vccd1 _14521_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_195_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23588_ _23588_/CLK _23588_/D vssd1 vssd1 vccd1 vccd1 _23588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13341_ _13344_/B _13375_/B vssd1 vssd1 vccd1 vccd1 _13341_/X sky130_fd_sc_hd__or2_1
X_22539_ _23511_/CLK _22539_/D vssd1 vssd1 vccd1 vccd1 _22539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_328_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16060_ _16059_/X _14509_/A _14513_/A _22974_/Q vssd1 vssd1 vccd1 vccd1 _16060_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_185_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13272_ _15929_/A _13262_/X _13271_/X _13765_/A vssd1 vssd1 vccd1 vccd1 _13273_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_183_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15011_ _15011_/A vssd1 vssd1 vccd1 vccd1 _15020_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_12223_ _12387_/A _12222_/X _11819_/A vssd1 vssd1 vccd1 vccd1 _12223_/X sky130_fd_sc_hd__o21a_1
XFILLER_343_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_335_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12154_ _12007_/A _12153_/X _12797_/A vssd1 vssd1 vccd1 vccd1 _12154_/X sky130_fd_sc_hd__o21a_1
XFILLER_151_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_311_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_297_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_296_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11105_ _13421_/A _13470_/A vssd1 vssd1 vccd1 vccd1 _11106_/A sky130_fd_sc_hd__or2_2
X_19750_ _19236_/X _23515_/Q _19754_/S vssd1 vssd1 vccd1 vccd1 _19751_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16962_ _16962_/A _21294_/C vssd1 vssd1 vccd1 vccd1 _16984_/B sky130_fd_sc_hd__or2_1
X_12085_ _12078_/Y _12080_/Y _12082_/Y _12084_/Y _11243_/A vssd1 vssd1 vccd1 vccd1
+ _12085_/X sky130_fd_sc_hd__o221a_1
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_311_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18701_ _18701_/A vssd1 vssd1 vccd1 vccd1 _23077_/D sky130_fd_sc_hd__clkbuf_1
X_15913_ _22938_/Q _15000_/A _15001_/A _22970_/Q vssd1 vssd1 vccd1 vccd1 _15913_/X
+ sky130_fd_sc_hd__o22a_1
X_19681_ _19681_/A vssd1 vssd1 vccd1 vccd1 _23484_/D sky130_fd_sc_hd__clkbuf_1
X_16893_ _16892_/X _22545_/Q _16893_/S vssd1 vssd1 vccd1 vccd1 _16894_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15844_ _15885_/A _15844_/B vssd1 vssd1 vccd1 vccd1 _15844_/Y sky130_fd_sc_hd__nand2_1
X_18632_ _23047_/Q _17553_/X _18636_/S vssd1 vssd1 vccd1 vccd1 _18633_/A sky130_fd_sc_hd__mux2_1
XFILLER_264_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_292_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18563_ _18563_/A vssd1 vssd1 vccd1 vccd1 _23016_/D sky130_fd_sc_hd__clkbuf_1
X_15775_ _15775_/A _15775_/B vssd1 vssd1 vccd1 vccd1 _15775_/Y sky130_fd_sc_hd__nor2_1
X_12987_ _12981_/X _12986_/X _13718_/A vssd1 vssd1 vccd1 vccd1 _12988_/B sky130_fd_sc_hd__o21ai_2
XFILLER_280_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17514_ _22664_/Q _16265_/X _17516_/S vssd1 vssd1 vccd1 vccd1 _17515_/A sky130_fd_sc_hd__mux2_1
X_14726_ _13706_/A _14716_/X _14721_/X _14725_/X vssd1 vssd1 vccd1 vccd1 _21206_/A
+ sky130_fd_sc_hd__a2bb2o_4
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18494_ _18520_/A vssd1 vssd1 vccd1 vccd1 _18494_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11938_ _11939_/A _11939_/B vssd1 vssd1 vccd1 vccd1 _11940_/A sky130_fd_sc_hd__and2_4
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_339_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17445_ _17456_/A vssd1 vssd1 vccd1 vccd1 _17454_/S sky130_fd_sc_hd__buf_2
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14657_ _14330_/X _14297_/X _14664_/S vssd1 vssd1 vccd1 vccd1 _14657_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11869_ _12269_/A vssd1 vssd1 vccd1 vccd1 _11869_/X sky130_fd_sc_hd__buf_4
XFILLER_21_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13608_ _13608_/A _13608_/B vssd1 vssd1 vccd1 vccd1 _13608_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17376_ _22608_/Q _14148_/A _17380_/S vssd1 vssd1 vccd1 vccd1 _17377_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_300_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14588_ _14588_/A vssd1 vssd1 vccd1 vccd1 _15903_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_308_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19115_ _19161_/S vssd1 vssd1 vccd1 vccd1 _19124_/S sky130_fd_sc_hd__buf_4
X_16327_ _15104_/X _22331_/Q _16333_/S vssd1 vssd1 vccd1 vccd1 _16328_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13539_ _12743_/B _13534_/Y _13538_/X _12741_/Y vssd1 vssd1 vccd1 vccd1 _13632_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_347_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19046_ _19046_/A vssd1 vssd1 vccd1 vccd1 _23216_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_307_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16258_ _16258_/A vssd1 vssd1 vccd1 vccd1 _22308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_316_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15209_ _19975_/D _14901_/X _14902_/X _23629_/Q vssd1 vssd1 vccd1 vccd1 _15209_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_126_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16189_ _15676_/A _21283_/A _16188_/Y _20493_/B vssd1 vssd1 vccd1 vccd1 _16189_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_303_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_331_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19948_ _23598_/Q _19944_/B _19947_/Y vssd1 vssd1 vccd1 vccd1 _23598_/D sky130_fd_sc_hd__o21a_1
XFILLER_275_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_9 _22193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19879_ _16255_/X _23572_/Q _19887_/S vssd1 vssd1 vccd1 vccd1 _19880_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21910_ _23832_/Q _23766_/Q vssd1 vssd1 vccd1 vccd1 _21910_/Y sky130_fd_sc_hd__nand2_1
X_22890_ _23009_/CLK _22890_/D vssd1 vssd1 vccd1 vccd1 _22890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21841_ _21841_/A vssd1 vssd1 vccd1 vccd1 _21900_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_167_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21772_ _21790_/A _21845_/A vssd1 vssd1 vccd1 vccd1 _21772_/Y sky130_fd_sc_hd__nor2_1
XPHY_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23511_ _23511_/CLK _23511_/D vssd1 vssd1 vccd1 vccd1 _23511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_358_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20723_ _20723_/A _20731_/B vssd1 vssd1 vccd1 vccd1 _20727_/B sky130_fd_sc_hd__and2_2
XFILLER_24_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_357_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23442_ _23503_/CLK _23442_/D vssd1 vssd1 vccd1 vccd1 _23442_/Q sky130_fd_sc_hd__dfxtp_1
X_20654_ _20654_/A vssd1 vssd1 vccd1 vccd1 _20655_/A sky130_fd_sc_hd__inv_2
XFILLER_286_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20585_ _20585_/A vssd1 vssd1 vccd1 vccd1 _20588_/A sky130_fd_sc_hd__inv_2
XFILLER_104_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23373_ _23407_/CLK _23373_/D vssd1 vssd1 vccd1 vccd1 _23373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_358_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_338_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22324_ _23577_/CLK _22324_/D vssd1 vssd1 vccd1 vccd1 _22324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_286_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_353_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22255_ _22255_/A vssd1 vssd1 vccd1 vccd1 _23944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21206_ _21206_/A _21227_/B vssd1 vssd1 vccd1 vccd1 _21206_/Y sky130_fd_sc_hd__nand2_1
XFILLER_151_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_340_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22186_ _23842_/Q _23776_/Q vssd1 vssd1 vccd1 vccd1 _22187_/B sky130_fd_sc_hd__nand2_1
XFILLER_160_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21137_ _22260_/A _21137_/B vssd1 vssd1 vccd1 vccd1 _23862_/D sky130_fd_sc_hd__nor2_1
XFILLER_235_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21068_ _23842_/Q _21068_/B vssd1 vssd1 vccd1 vccd1 _21068_/X sky130_fd_sc_hd__or2_1
XFILLER_293_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20019_ _23617_/Q _20031_/C _23618_/Q vssd1 vssd1 vccd1 vccd1 _20022_/B sky130_fd_sc_hd__a21oi_1
X_12910_ _12904_/A _12907_/X _12909_/X _12797_/X vssd1 vssd1 vccd1 vccd1 _12910_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_247_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13890_ _13890_/A _13890_/B vssd1 vssd1 vccd1 vccd1 _13890_/Y sky130_fd_sc_hd__nor2_2
XFILLER_101_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12841_ _23934_/Q vssd1 vssd1 vccd1 vccd1 _12841_/Y sky130_fd_sc_hd__inv_2
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15003_/A _15547_/X _15559_/X vssd1 vssd1 vccd1 vccd1 _15560_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_215_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12772_ _12765_/Y _12767_/Y _12769_/Y _12771_/Y _11559_/A vssd1 vssd1 vccd1 vccd1
+ _12772_/X sky130_fd_sc_hd__o221a_2
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14511_ _14933_/A vssd1 vssd1 vccd1 vccd1 _14753_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_187_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11723_/A _11723_/B vssd1 vssd1 vccd1 vccd1 _11723_/Y sky130_fd_sc_hd__nor2_1
XFILLER_214_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23709_ _23714_/CLK _23709_/D vssd1 vssd1 vccd1 vccd1 _23709_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_15_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _14629_/A _15490_/X _15491_/S vssd1 vssd1 vccd1 vccd1 _15491_/X sky130_fd_sc_hd__mux2_1
XFILLER_349_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17230_/A vssd1 vssd1 vccd1 vccd1 _17230_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14442_ _22914_/Q _14868_/B vssd1 vssd1 vccd1 vccd1 _14442_/X sky130_fd_sc_hd__and2_1
XFILLER_159_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _23414_/Q _23030_/Q _23382_/Q _23350_/Q _12029_/A _11676_/A vssd1 vssd1 vccd1
+ vccd1 _11655_/B sky130_fd_sc_hd__mux4_2
XFILLER_302_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17161_ _22811_/Q _17244_/B _17244_/C vssd1 vssd1 vccd1 vccd1 _17169_/A sky130_fd_sc_hd__and3_1
XFILLER_196_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14373_ _14373_/A _15079_/B vssd1 vssd1 vccd1 vccd1 _14647_/A sky130_fd_sc_hd__and2_1
X_11585_ _12119_/S vssd1 vssd1 vccd1 vccd1 _12042_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_7_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16112_ _14690_/X _16094_/Y _16098_/X _17298_/A _15964_/A vssd1 vssd1 vccd1 vccd1
+ _16112_/X sky130_fd_sc_hd__o32a_1
XFILLER_344_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13324_ _13601_/A _13324_/B vssd1 vssd1 vccd1 vccd1 _13400_/A sky130_fd_sc_hd__xnor2_4
XFILLER_317_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17092_ _17276_/A vssd1 vssd1 vccd1 vccd1 _17132_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_183_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16043_ _15318_/A _16038_/X _16042_/Y vssd1 vssd1 vccd1 vccd1 _16043_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_127_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13255_ _22482_/Q _22642_/Q _13255_/S vssd1 vssd1 vccd1 vccd1 _13255_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_332_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12206_ _12206_/A vssd1 vssd1 vccd1 vccd1 _12596_/B sky130_fd_sc_hd__buf_2
XFILLER_313_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_57_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23572_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13186_ _13187_/A _13240_/A vssd1 vssd1 vccd1 vccd1 _13188_/A sky130_fd_sc_hd__and2_2
XFILLER_124_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19802_ _23538_/Q _19207_/A _19804_/S vssd1 vssd1 vccd1 vccd1 _19803_/A sky130_fd_sc_hd__mux2_1
X_12137_ _23923_/Q vssd1 vssd1 vccd1 vccd1 _12137_/Y sky130_fd_sc_hd__inv_2
XFILLER_296_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17994_ _22840_/Q _17981_/X _17993_/X _17979_/X vssd1 vssd1 vccd1 vccd1 _22840_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_229_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_300_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19733_ _19733_/A vssd1 vssd1 vccd1 vccd1 _23507_/D sky130_fd_sc_hd__clkbuf_1
X_16945_ _16945_/A _16945_/B vssd1 vssd1 vccd1 vccd1 _16945_/Y sky130_fd_sc_hd__nand2_1
X_12068_ _12082_/A _12067_/X _11230_/A vssd1 vssd1 vccd1 vccd1 _12068_/X sky130_fd_sc_hd__o21a_1
XFILLER_237_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19664_ _19664_/A vssd1 vssd1 vccd1 vccd1 _23476_/D sky130_fd_sc_hd__clkbuf_1
X_16876_ _19226_/A vssd1 vssd1 vccd1 vccd1 _16876_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_265_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18615_ _16902_/X _23040_/Q _18619_/S vssd1 vssd1 vccd1 vccd1 _18616_/A sky130_fd_sc_hd__mux2_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _23933_/Q _15828_/B vssd1 vssd1 vccd1 vccd1 _15924_/C sky130_fd_sc_hd__and2_2
XFILLER_92_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19595_ _23446_/Q _19220_/A _19599_/S vssd1 vssd1 vccd1 vccd1 _19596_/A sky130_fd_sc_hd__mux2_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18546_ _21220_/A vssd1 vssd1 vccd1 vccd1 _20324_/A sky130_fd_sc_hd__clkbuf_2
X_15758_ _23737_/Q _23867_/Q _16138_/S vssd1 vssd1 vccd1 vccd1 _15758_/X sky130_fd_sc_hd__mux2_1
XFILLER_240_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14709_ _22980_/Q _14137_/A _14980_/A input237/X vssd1 vssd1 vccd1 vccd1 _21350_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_178_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18477_ _18467_/X _18475_/Y _18476_/X vssd1 vssd1 vccd1 vccd1 _22986_/D sky130_fd_sc_hd__a21oi_1
X_15689_ _23799_/Q _15219_/X _14606_/X vssd1 vssd1 vccd1 vccd1 _15689_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_339_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17428_ _22626_/Q _16246_/X _17432_/S vssd1 vssd1 vccd1 vccd1 _17429_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_348_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17359_ _17359_/A vssd1 vssd1 vccd1 vccd1 _22600_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_348_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20370_ _20227_/X _20368_/X _20369_/Y _20196_/X vssd1 vssd1 vccd1 vccd1 _20370_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_308_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_307_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_3_1_wb_clk_i clkbuf_3_3_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19029_ _16828_/X _23209_/Q _19029_/S vssd1 vssd1 vccd1 vccd1 _19030_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22040_ _22040_/A _22040_/B vssd1 vssd1 vccd1 vccd1 _22040_/Y sky130_fd_sc_hd__nand2_1
XFILLER_288_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22942_ _22947_/CLK _22942_/D vssd1 vssd1 vccd1 vccd1 _22942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22873_ _23592_/CLK _22873_/D vssd1 vssd1 vccd1 vccd1 _22873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21824_ _21793_/A _21793_/B _21792_/A vssd1 vssd1 vccd1 vccd1 _21828_/A sky130_fd_sc_hd__a21oi_2
XFILLER_225_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21755_ _23827_/Q _23761_/Q vssd1 vssd1 vccd1 vccd1 _21756_/B sky130_fd_sc_hd__nor2_1
XFILLER_24_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_357_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_297_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20706_ _20763_/A vssd1 vssd1 vccd1 vccd1 _20706_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21686_ _20264_/A _21841_/A _21619_/B _15377_/X vssd1 vssd1 vccd1 vccd1 _21686_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_196_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23425_ _23453_/CLK _23425_/D vssd1 vssd1 vccd1 vccd1 _23425_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20637_ _20763_/A vssd1 vssd1 vccd1 vccd1 _20637_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_326_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23356_ _23420_/CLK _23356_/D vssd1 vssd1 vccd1 vccd1 _23356_/Q sky130_fd_sc_hd__dfxtp_1
X_11370_ _23332_/Q _23300_/Q _23268_/Q _23556_/Q _11468_/A _11365_/X vssd1 vssd1 vccd1
+ vccd1 _11370_/X sky130_fd_sc_hd__mux4_1
X_20568_ _20591_/A _20779_/B _20568_/C vssd1 vssd1 vccd1 vccd1 _20568_/X sky130_fd_sc_hd__or3_1
XFILLER_326_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22307_ _23571_/CLK _22307_/D vssd1 vssd1 vccd1 vccd1 _22307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_353_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_291_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_341_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23287_ _23543_/CLK _23287_/D vssd1 vssd1 vccd1 vccd1 _23287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_314_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_298_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20499_ _21077_/D _20499_/B _21517_/B vssd1 vssd1 vccd1 vccd1 _20500_/B sky130_fd_sc_hd__and3_1
XFILLER_316_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13040_ _23232_/Q _23200_/Q _23168_/Q _23136_/Q _13032_/S _11435_/A vssd1 vssd1 vccd1
+ vccd1 _13041_/B sky130_fd_sc_hd__mux4_1
XFILLER_4_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22238_ _16194_/X _22235_/Y _22236_/X _21767_/X vssd1 vssd1 vccd1 vccd1 _22238_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22169_ _22168_/Y _22142_/C _22142_/B vssd1 vssd1 vccd1 vccd1 _22170_/B sky130_fd_sc_hd__a21oi_2
XFILLER_133_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14991_ _19934_/B _14901_/X _14902_/X _23626_/Q vssd1 vssd1 vccd1 vccd1 _14991_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_278_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_294_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16730_ _16730_/A vssd1 vssd1 vccd1 vccd1 _16730_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13942_ _13942_/A _13942_/B vssd1 vssd1 vccd1 vccd1 _13943_/B sky130_fd_sc_hd__or2_2
XFILLER_293_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_332_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16661_ _16661_/A vssd1 vssd1 vccd1 vccd1 _22477_/D sky130_fd_sc_hd__clkbuf_1
X_13873_ _13873_/A vssd1 vssd1 vccd1 vccd1 _13873_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_175_wb_clk_i _23931_/CLK vssd1 vssd1 vccd1 vccd1 _23942_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18400_ _22960_/Q _22961_/Q _18400_/C vssd1 vssd1 vccd1 vccd1 _18402_/B sky130_fd_sc_hd__and3_1
XFILLER_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15612_ _15701_/C _15612_/B vssd1 vssd1 vccd1 vccd1 _15612_/Y sky130_fd_sc_hd__nor2_2
XFILLER_290_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12824_ _12926_/A _12824_/B vssd1 vssd1 vccd1 vccd1 _12824_/Y sky130_fd_sc_hd__nor2_1
XFILLER_262_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19380_ _19380_/A vssd1 vssd1 vccd1 vccd1 _23350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_290_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16592_ _16592_/A vssd1 vssd1 vccd1 vccd1 _16601_/S sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_104_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23391_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18331_ _15833_/X _18332_/C _22937_/Q vssd1 vssd1 vccd1 vccd1 _18333_/B sky130_fd_sc_hd__a21oi_1
X_15543_ _12005_/Y _14259_/A _14674_/A _13615_/A vssd1 vssd1 vccd1 vccd1 _15543_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12755_ _12755_/A vssd1 vssd1 vccd1 vccd1 _12755_/X sky130_fd_sc_hd__buf_4
XFILLER_188_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ _18263_/A _18263_/B _22916_/Q vssd1 vssd1 vccd1 vccd1 _18264_/B sky130_fd_sc_hd__a21oi_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _11706_/A vssd1 vssd1 vccd1 vccd1 _11706_/X sky130_fd_sc_hd__clkbuf_4
X_15474_ _19207_/A vssd1 vssd1 vccd1 vccd1 _15474_/X sky130_fd_sc_hd__clkbuf_2
X_12686_ _22376_/Q _22408_/Q _22697_/Q _23064_/Q _12977_/S _12685_/X vssd1 vssd1 vccd1
+ vccd1 _12686_/X sky130_fd_sc_hd__mux4_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17213_ _14393_/X _17009_/S _17212_/X vssd1 vssd1 vccd1 vccd1 _17213_/X sky130_fd_sc_hd__o21a_1
X_14425_ _21448_/B _15929_/A _14421_/S _14424_/X vssd1 vssd1 vccd1 vccd1 _14465_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_30_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_348_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18193_ _18118_/X _18163_/A _18186_/X _18191_/X _18192_/X vssd1 vssd1 vccd1 vccd1
+ _22892_/D sky130_fd_sc_hd__o221a_1
X_11637_ _11637_/A vssd1 vssd1 vccd1 vccd1 _11637_/X sky130_fd_sc_hd__buf_4
XFILLER_202_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_357_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17144_ _17144_/A vssd1 vssd1 vccd1 vccd1 _17172_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_345_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14356_ _14358_/A _14356_/B vssd1 vssd1 vccd1 vccd1 _14356_/Y sky130_fd_sc_hd__nor2_1
XFILLER_317_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11568_ _11568_/A vssd1 vssd1 vccd1 vccd1 _12749_/A sky130_fd_sc_hd__buf_6
XFILLER_155_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13307_ _13307_/A _16128_/S vssd1 vssd1 vccd1 vccd1 _13311_/A sky130_fd_sc_hd__nor2_1
XFILLER_116_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_345_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17075_ _17222_/B vssd1 vssd1 vccd1 vccd1 _17116_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_171_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14287_ _14356_/B vssd1 vssd1 vccd1 vccd1 _14287_/Y sky130_fd_sc_hd__clkinv_2
X_11499_ _11502_/A _11498_/X _11236_/A vssd1 vssd1 vccd1 vccd1 _11499_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_226_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16026_ _23712_/Q _15210_/X _16025_/X vssd1 vssd1 vccd1 vccd1 _16026_/Y sky130_fd_sc_hd__o21ai_4
X_13238_ _13574_/A _13579_/A vssd1 vssd1 vccd1 vccd1 _13239_/C sky130_fd_sc_hd__nor2_1
XFILLER_108_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_313_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_300_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13169_ _13218_/A _13169_/B vssd1 vssd1 vccd1 vccd1 _13169_/X sky130_fd_sc_hd__or2_1
XFILLER_111_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17977_ input1/X input267/X _17987_/S vssd1 vssd1 vccd1 vccd1 _17977_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater503 _13455_/Y vssd1 vssd1 vccd1 vccd1 output441/A sky130_fd_sc_hd__buf_6
XFILLER_300_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_300_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19716_ _19716_/A vssd1 vssd1 vccd1 vccd1 _23499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_348_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16928_ _17237_/A vssd1 vssd1 vccd1 vccd1 _17109_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_238_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19647_ _19191_/X _23469_/Q _19649_/S vssd1 vssd1 vccd1 vccd1 _19648_/A sky130_fd_sc_hd__mux2_1
XFILLER_226_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16859_ _16859_/A vssd1 vssd1 vccd1 vccd1 _22534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19578_ _19578_/A vssd1 vssd1 vccd1 vccd1 _23438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18529_ _18520_/X _18528_/Y _18264_/A vssd1 vssd1 vccd1 vccd1 _23006_/D sky130_fd_sc_hd__a21oi_1
XFILLER_178_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21540_ _21516_/X _21538_/X _21539_/Y vssd1 vssd1 vccd1 vccd1 _23918_/D sky130_fd_sc_hd__a21oi_1
XFILLER_328_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_327_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21471_ _21403_/A _21401_/A _21403_/B _21432_/Y _21400_/Y vssd1 vssd1 vccd1 vccd1
+ _21472_/C sky130_fd_sc_hd__o311a_1
XFILLER_21_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23210_ _23466_/CLK _23210_/D vssd1 vssd1 vccd1 vccd1 _23210_/Q sky130_fd_sc_hd__dfxtp_1
X_20422_ _23688_/Q _20429_/B vssd1 vssd1 vccd1 vccd1 _20422_/X sky130_fd_sc_hd__or2_1
XFILLER_119_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_323_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23141_ _23527_/CLK _23141_/D vssd1 vssd1 vccd1 vccd1 _23141_/Q sky130_fd_sc_hd__dfxtp_1
X_20353_ _20353_/A _20400_/B vssd1 vssd1 vccd1 vccd1 _20355_/B sky130_fd_sc_hd__nor2_1
XFILLER_335_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_350_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23072_ _23391_/CLK _23072_/D vssd1 vssd1 vccd1 vccd1 _23072_/Q sky130_fd_sc_hd__dfxtp_1
X_20284_ _23667_/Q _20338_/B vssd1 vssd1 vccd1 vccd1 _20284_/X sky130_fd_sc_hd__or2_1
XFILLER_136_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_304_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_351_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22023_ _22023_/A _22023_/B vssd1 vssd1 vccd1 vccd1 _22024_/B sky130_fd_sc_hd__nor2_1
XTAP_6229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_289_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_303_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23370_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_275_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22925_ _22929_/CLK _22925_/D vssd1 vssd1 vccd1 vccd1 _22925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22856_ _22908_/CLK _22856_/D vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21807_ _17163_/A _21867_/A _21806_/X _21556_/X vssd1 vssd1 vccd1 vccd1 _21809_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22787_ _23567_/CLK _22787_/D vssd1 vssd1 vccd1 vccd1 _22787_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _23901_/Q _12539_/X _11843_/A vssd1 vssd1 vccd1 vccd1 _12540_/Y sky130_fd_sc_hd__o21ai_1
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21738_ _21738_/A _21741_/A vssd1 vssd1 vccd1 vccd1 _21739_/B sky130_fd_sc_hd__or2_1
XFILLER_40_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12471_ _12468_/X _12469_/Y _12470_/Y vssd1 vssd1 vccd1 vccd1 _13505_/A sky130_fd_sc_hd__a21oi_2
XFILLER_358_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21669_ _21669_/A _21669_/B vssd1 vssd1 vccd1 vccd1 _21669_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_327_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14210_ _15618_/A vssd1 vssd1 vccd1 vccd1 _14210_/X sky130_fd_sc_hd__clkbuf_4
X_23408_ _23951_/A _23408_/D vssd1 vssd1 vccd1 vccd1 _23408_/Q sky130_fd_sc_hd__dfxtp_1
X_11422_ _13259_/A _11421_/X _11236_/X vssd1 vssd1 vccd1 vccd1 _11422_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_327_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15190_ _13739_/A _15186_/Y _15189_/Y _13875_/C vssd1 vssd1 vccd1 vccd1 _15190_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_126_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_314_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14141_ _23012_/Q _18536_/A _18537_/B vssd1 vssd1 vccd1 vccd1 _16945_/A sky130_fd_sc_hd__or3_4
XFILLER_126_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_327_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11353_ _11353_/A vssd1 vssd1 vccd1 vccd1 _15671_/A sky130_fd_sc_hd__buf_8
X_23339_ _23531_/CLK _23339_/D vssd1 vssd1 vccd1 vccd1 _23339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_327_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_342_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14072_ _14072_/A _14072_/B _14072_/C vssd1 vssd1 vccd1 vccd1 _14072_/X sky130_fd_sc_hd__and3_1
XFILLER_314_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11284_ _11284_/A vssd1 vssd1 vccd1 vccd1 _11285_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17900_ _18009_/B _17894_/X _17896_/X _14119_/C _17899_/X vssd1 vssd1 vccd1 vccd1
+ _17900_/X sky130_fd_sc_hd__a221o_1
X_13023_ _13492_/B _13388_/B vssd1 vssd1 vccd1 vccd1 _13023_/X sky130_fd_sc_hd__or2_1
XFILLER_341_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18880_ _18880_/A vssd1 vssd1 vccd1 vccd1 _23142_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17831_ _22788_/Q _17582_/X _17837_/S vssd1 vssd1 vccd1 vccd1 _17832_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17762_ _17762_/A vssd1 vssd1 vccd1 vccd1 _22757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14974_ _23915_/Q _14976_/B vssd1 vssd1 vccd1 vccd1 _15049_/C sky130_fd_sc_hd__and2_1
X_19501_ _19188_/X _23404_/Q _19505_/S vssd1 vssd1 vccd1 vccd1 _19502_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16713_ _22492_/Q _16711_/X _16712_/X input37/X vssd1 vssd1 vccd1 vccd1 _16714_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_75_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13925_ _13918_/X _15078_/A _13923_/Y _13924_/X vssd1 vssd1 vccd1 vccd1 _14091_/A
+ sky130_fd_sc_hd__a211o_4
X_17693_ _22727_/Q _17591_/X _17693_/S vssd1 vssd1 vccd1 vccd1 _17694_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19432_ _19432_/A vssd1 vssd1 vccd1 vccd1 _23373_/D sky130_fd_sc_hd__clkbuf_1
X_16644_ _16644_/A vssd1 vssd1 vccd1 vccd1 _22469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_263_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_403 _13990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13856_ _13856_/A vssd1 vssd1 vccd1 vccd1 _13856_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_290_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_414 _14037_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_425 _13432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_436 _23885_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12807_ _12807_/A vssd1 vssd1 vccd1 vccd1 _12807_/Y sky130_fd_sc_hd__inv_2
X_19363_ _19409_/S vssd1 vssd1 vccd1 vccd1 _19372_/S sky130_fd_sc_hd__buf_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_447 _14073_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16575_ _15668_/X _22439_/Q _16579_/S vssd1 vssd1 vccd1 vccd1 _16576_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13787_ _13787_/A vssd1 vssd1 vccd1 vccd1 _13787_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_458 _21681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_469 _12801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18314_ _18314_/A _22931_/Q _18314_/C vssd1 vssd1 vccd1 vccd1 _18315_/C sky130_fd_sc_hd__and3_1
XFILLER_188_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_349_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12738_ _13184_/A _12738_/B _12738_/C vssd1 vssd1 vccd1 vccd1 _21900_/A sky130_fd_sc_hd__nand3_4
X_15526_ _22993_/Q _15620_/A _15621_/A input221/X vssd1 vssd1 vccd1 vccd1 _21791_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_176_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ _19201_/X _23312_/Q _19300_/S vssd1 vssd1 vccd1 vccd1 _19295_/A sky130_fd_sc_hd__mux2_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_337_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18245_ _18245_/A vssd1 vssd1 vccd1 vccd1 _18245_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15457_ _15088_/S _15014_/X _15491_/S vssd1 vssd1 vccd1 vccd1 _15457_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_336_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12669_ _22796_/Q _22764_/Q _22665_/Q _22732_/Q _12750_/S _12041_/X vssd1 vssd1 vccd1
+ vccd1 _12670_/B sky130_fd_sc_hd__mux4_2
X_14408_ _22904_/Q _14153_/X _14164_/A _22597_/Q vssd1 vssd1 vccd1 vccd1 _14550_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_352_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_72_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23354_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18176_ _18170_/X _18173_/X _18175_/X vssd1 vssd1 vccd1 vccd1 _18176_/Y sky130_fd_sc_hd__a21oi_1
X_15388_ _13497_/A _14251_/A _14760_/A vssd1 vssd1 vccd1 vccd1 _15388_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17127_ _17283_/A vssd1 vssd1 vccd1 vccd1 _17127_/X sky130_fd_sc_hd__clkbuf_2
X_14339_ _12602_/A _14276_/B _15171_/A vssd1 vssd1 vccd1 vccd1 _14339_/X sky130_fd_sc_hd__mux2_1
XFILLER_317_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_289_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17058_ _17000_/X _17051_/X _17056_/X _17057_/X vssd1 vssd1 vccd1 vccd1 _17058_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16009_ _21078_/A _15617_/X _15618_/X vssd1 vssd1 vccd1 vccd1 _16009_/Y sky130_fd_sc_hd__o21ai_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_297_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20971_ _22116_/A _20966_/X _20736_/B _20970_/X vssd1 vssd1 vccd1 vccd1 _20971_/X
+ sky130_fd_sc_hd__a211o_1
X_22710_ _23846_/CLK _22710_/D vssd1 vssd1 vccd1 vccd1 _22710_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23690_ _23696_/CLK _23690_/D vssd1 vssd1 vccd1 vccd1 _23690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22641_ _23422_/CLK _22641_/D vssd1 vssd1 vccd1 vccd1 _22641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_322_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22572_ _23646_/CLK _22572_/D vssd1 vssd1 vccd1 vccd1 _22572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_322_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_328_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21523_ _16016_/A _21549_/A _21521_/Y _21522_/X vssd1 vssd1 vccd1 vccd1 _21546_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_355_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_327_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21454_ _21454_/A _21454_/B vssd1 vssd1 vccd1 vccd1 _21454_/X sky130_fd_sc_hd__xor2_1
XFILLER_308_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_309_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20405_ _20213_/A _20765_/A _20404_/X _20392_/X vssd1 vssd1 vccd1 vccd1 _23684_/D
+ sky130_fd_sc_hd__o211a_1
X_21385_ _11084_/A _21518_/A _21482_/A vssd1 vssd1 vccd1 vccd1 _21553_/A sky130_fd_sc_hd__a21o_1
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23124_ _23543_/CLK _23124_/D vssd1 vssd1 vccd1 vccd1 _23124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_335_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20336_ _20355_/A _20336_/B vssd1 vssd1 vccd1 vccd1 _20336_/Y sky130_fd_sc_hd__nand2_1
XFILLER_350_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23055_ _23567_/CLK _23055_/D vssd1 vssd1 vccd1 vccd1 _23055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20267_ _20376_/A _20267_/B vssd1 vssd1 vccd1 vccd1 _20267_/Y sky130_fd_sc_hd__nor2_1
XTAP_6037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_288_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22006_ _21999_/A _21984_/X _22005_/Y _21896_/X vssd1 vssd1 vccd1 vccd1 _23933_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput103 dout0[6] vssd1 vssd1 vccd1 vccd1 input103/X sky130_fd_sc_hd__buf_2
Xinput114 dout1[16] vssd1 vssd1 vccd1 vccd1 input114/X sky130_fd_sc_hd__clkbuf_1
XTAP_5325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20198_ _14939_/B _20154_/X _20199_/B vssd1 vssd1 vccd1 vccd1 _20198_/X sky130_fd_sc_hd__a21o_1
Xinput125 dout1[26] vssd1 vssd1 vccd1 vccd1 input125/X sky130_fd_sc_hd__clkbuf_1
XFILLER_277_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput136 dout1[36] vssd1 vssd1 vccd1 vccd1 input136/X sky130_fd_sc_hd__buf_2
XTAP_5347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput147 dout1[46] vssd1 vssd1 vccd1 vccd1 input147/X sky130_fd_sc_hd__buf_2
XFILLER_292_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput158 dout1[56] vssd1 vssd1 vccd1 vccd1 input158/X sky130_fd_sc_hd__buf_2
XTAP_5369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput169 dout1[8] vssd1 vssd1 vccd1 vccd1 input169/X sky130_fd_sc_hd__clkbuf_1
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ _11141_/A _11970_/X _11598_/X vssd1 vssd1 vccd1 vccd1 _11971_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_245_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13710_ _13710_/A _13718_/D vssd1 vssd1 vccd1 vccd1 _13711_/B sky130_fd_sc_hd__nand2_4
X_22908_ _22908_/CLK _22908_/D vssd1 vssd1 vccd1 vccd1 _22908_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _14690_/A vssd1 vssd1 vccd1 vccd1 _14690_/X sky130_fd_sc_hd__clkbuf_4
X_23888_ _23888_/CLK _23888_/D vssd1 vssd1 vccd1 vccd1 _23888_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_260_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13641_ _13647_/A vssd1 vssd1 vccd1 vccd1 _21293_/A sky130_fd_sc_hd__clkbuf_4
X_22839_ _23632_/CLK _22839_/D vssd1 vssd1 vccd1 vccd1 _22839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _15823_/X _22346_/Q _16366_/S vssd1 vssd1 vccd1 vccd1 _16361_/A sky130_fd_sc_hd__mux2_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _23936_/Q vssd1 vssd1 vccd1 vccd1 _22087_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_213_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_347_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_319_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15311_ _18296_/A _14932_/X _14934_/X _22956_/Q vssd1 vssd1 vccd1 vccd1 _15311_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_200_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _12523_/A _12523_/B vssd1 vssd1 vccd1 vccd1 _12523_/Y sky130_fd_sc_hd__nor2_1
X_16291_ _18856_/A vssd1 vssd1 vccd1 vccd1 _16291_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_169_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18030_ hold3/A _18016_/X _18028_/X _18029_/X vssd1 vssd1 vccd1 vccd1 _22848_/D sky130_fd_sc_hd__o211a_1
X_15242_ _15242_/A vssd1 vssd1 vccd1 vccd1 _22269_/D sky130_fd_sc_hd__clkbuf_1
X_12454_ _11843_/A _12446_/Y _12448_/Y _12451_/Y _12453_/Y vssd1 vssd1 vccd1 vccd1
+ _12454_/X sky130_fd_sc_hd__o32a_1
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11405_ _11910_/A vssd1 vssd1 vccd1 vccd1 _12135_/A sky130_fd_sc_hd__buf_2
X_15173_ _13736_/B _15119_/B _15111_/X _13879_/B _14725_/A vssd1 vssd1 vccd1 vccd1
+ _15173_/X sky130_fd_sc_hd__o221a_1
X_12385_ _11330_/A _12384_/X _11819_/A vssd1 vssd1 vccd1 vccd1 _12385_/X sky130_fd_sc_hd__o21a_1
XFILLER_315_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14124_ _22893_/Q _18188_/B vssd1 vssd1 vccd1 vccd1 _18187_/B sky130_fd_sc_hd__or2_1
XFILLER_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11336_ _13229_/A vssd1 vssd1 vccd1 vccd1 _13131_/A sky130_fd_sc_hd__clkbuf_4
X_19981_ _19981_/A _19988_/C vssd1 vssd1 vccd1 vccd1 _19981_/Y sky130_fd_sc_hd__nor2_1
XFILLER_299_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_315_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18932_ _23166_/Q _18852_/X _18940_/S vssd1 vssd1 vccd1 vccd1 _18933_/A sky130_fd_sc_hd__mux2_1
XFILLER_286_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14055_ _14069_/B vssd1 vssd1 vccd1 vccd1 _14066_/B sky130_fd_sc_hd__clkbuf_1
XTAP_7250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11267_ _11267_/A vssd1 vssd1 vccd1 vccd1 _12087_/A sky130_fd_sc_hd__buf_2
XFILLER_4_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13006_ _13006_/A _13006_/B vssd1 vssd1 vccd1 vccd1 _13006_/X sky130_fd_sc_hd__or2_1
XTAP_7283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18863_ _23137_/Q _18862_/X _18866_/S vssd1 vssd1 vccd1 vccd1 _18864_/A sky130_fd_sc_hd__mux2_1
XTAP_6560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11198_ _22485_/Q _22645_/Q _13254_/S vssd1 vssd1 vccd1 vccd1 _11199_/B sky130_fd_sc_hd__mux2_1
XTAP_6571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_190_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23525_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17814_ _17814_/A vssd1 vssd1 vccd1 vccd1 _22780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18794_ _18794_/A vssd1 vssd1 vccd1 vccd1 _23115_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17745_ _17802_/S vssd1 vssd1 vccd1 vccd1 _17754_/S sky130_fd_sc_hd__buf_6
XFILLER_236_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14957_ _14384_/X _16034_/B _14956_/X _14839_/X vssd1 vssd1 vccd1 vccd1 _14958_/C
+ sky130_fd_sc_hd__o22a_2
XFILLER_303_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13908_ _13933_/A _14087_/A vssd1 vssd1 vccd1 vccd1 _13908_/Y sky130_fd_sc_hd__nor2_2
XFILLER_235_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_200 _13951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17676_ _22719_/Q _17566_/X _17682_/S vssd1 vssd1 vccd1 vccd1 _17677_/A sky130_fd_sc_hd__mux2_1
XFILLER_251_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14888_ _15367_/A _21384_/B _15479_/A vssd1 vssd1 vccd1 vccd1 _14888_/X sky130_fd_sc_hd__a21o_1
XINSDIODE2_211 _14494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19415_ _19415_/A vssd1 vssd1 vccd1 vccd1 _23365_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_222 _14939_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16627_ _22462_/Q _16233_/X _16629_/S vssd1 vssd1 vccd1 vccd1 _16628_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_233 _15155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_244 _15329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13839_ _15113_/A _13874_/C vssd1 vssd1 vccd1 vccd1 _13863_/B sky130_fd_sc_hd__nand2_2
XFILLER_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_255 _15602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_266 _15651_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19346_ _23335_/Q _18779_/X _19350_/S vssd1 vssd1 vccd1 vccd1 _19347_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_277 _15767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_288 _15959_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16558_ _16558_/A vssd1 vssd1 vccd1 vccd1 _22431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_338_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_299 _15990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15509_ _23827_/Q _14907_/A _15505_/X _15508_/X _14923_/A vssd1 vssd1 vccd1 vccd1
+ _15509_/X sky130_fd_sc_hd__a221o_1
X_19277_ _19277_/A vssd1 vssd1 vccd1 vccd1 _23304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16489_ _15474_/X _22402_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _16490_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_337_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18228_ _22855_/Q _18216_/X _18227_/X _18219_/X vssd1 vssd1 vccd1 vccd1 _22903_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_325_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_346_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18159_ _18159_/A _18159_/B vssd1 vssd1 vccd1 vccd1 _18160_/A sky130_fd_sc_hd__and2_1
XFILLER_175_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_333_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_352_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21170_ _23871_/Q _21168_/X _21169_/X _21163_/X vssd1 vssd1 vccd1 vccd1 _23871_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_321_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20121_ _20121_/A vssd1 vssd1 vccd1 vccd1 _20137_/A sky130_fd_sc_hd__buf_6
XFILLER_171_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20052_ _20066_/B _20066_/C _18268_/A vssd1 vssd1 vccd1 vccd1 _20052_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_258_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_286_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23811_ _23866_/CLK _23811_/D vssd1 vssd1 vccd1 vccd1 _23811_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_274_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23742_ _23915_/CLK _23742_/D vssd1 vssd1 vccd1 vccd1 _23742_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20954_ _20970_/A vssd1 vssd1 vccd1 vccd1 _20954_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23673_ _23706_/CLK _23673_/D vssd1 vssd1 vccd1 vccd1 _23673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20885_ _20762_/B _20810_/A _20811_/A _23779_/Q vssd1 vssd1 vccd1 vccd1 _20886_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_289_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22624_ _23047_/CLK _22624_/D vssd1 vssd1 vccd1 vccd1 _22624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22555_ _22968_/CLK _22555_/D vssd1 vssd1 vccd1 vccd1 _22555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21506_ _21491_/X _21498_/X _21505_/X vssd1 vssd1 vccd1 vccd1 _21506_/X sky130_fd_sc_hd__a21o_1
XFILLER_356_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22486_ _22520_/CLK _22486_/D vssd1 vssd1 vccd1 vccd1 _22486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_315_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21437_ _21437_/A _22197_/B vssd1 vssd1 vccd1 vccd1 _21437_/Y sky130_fd_sc_hd__nor2_1
XFILLER_257_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_324_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_324_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12170_ _12170_/A vssd1 vssd1 vccd1 vccd1 _12171_/B sky130_fd_sc_hd__inv_2
XFILLER_107_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21368_ _22025_/A vssd1 vssd1 vccd1 vccd1 _21418_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11121_ _12260_/A vssd1 vssd1 vccd1 vccd1 _12134_/A sky130_fd_sc_hd__buf_8
X_23107_ _23459_/CLK _23107_/D vssd1 vssd1 vccd1 vccd1 _23107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_218_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20319_ _15738_/A _20215_/X _20318_/X vssd1 vssd1 vccd1 vccd1 _20319_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_296_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21299_ _21465_/A vssd1 vssd1 vccd1 vccd1 _21479_/A sky130_fd_sc_hd__buf_4
XFILLER_104_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23038_ _23550_/CLK _23038_/D vssd1 vssd1 vccd1 vccd1 _23038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_277_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_276_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15860_ _18843_/A vssd1 vssd1 vccd1 vccd1 _19236_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_277_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14811_ _19172_/A vssd1 vssd1 vccd1 vccd1 _14811_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _21950_/A _15790_/C _23932_/Q vssd1 vssd1 vccd1 vccd1 _15792_/B sky130_fd_sc_hd__a21oi_1
XFILLER_291_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _22671_/Q _16287_/X _17538_/S vssd1 vssd1 vccd1 vccd1 _17531_/A sky130_fd_sc_hd__mux2_1
XFILLER_292_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11954_ _22308_/Q _23444_/Q _12043_/S vssd1 vssd1 vccd1 vccd1 _11954_/X sky130_fd_sc_hd__mux2_1
XFILLER_245_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14742_ _14916_/A vssd1 vssd1 vccd1 vccd1 _14742_/X sky130_fd_sc_hd__buf_4
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17461_ _22641_/Q _16294_/X _17465_/S vssd1 vssd1 vccd1 vccd1 _17462_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14673_ _20205_/A _15176_/A vssd1 vssd1 vccd1 vccd1 _14674_/A sky130_fd_sc_hd__nor2_4
X_11885_ _11828_/B _21596_/A _11884_/Y vssd1 vssd1 vccd1 vccd1 _13523_/B sky130_fd_sc_hd__a21bo_1
XFILLER_225_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19200_ _19200_/A vssd1 vssd1 vccd1 vccd1 _23279_/D sky130_fd_sc_hd__clkbuf_1
X_16412_ _15372_/X _22368_/Q _16418_/S vssd1 vssd1 vccd1 vccd1 _16413_/A sky130_fd_sc_hd__mux2_1
X_13624_ _23923_/Q vssd1 vssd1 vccd1 vccd1 _21708_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_260_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17392_ _21185_/A vssd1 vssd1 vccd1 vccd1 _21681_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_347_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19131_ _23254_/Q _18827_/X _19135_/S vssd1 vssd1 vccd1 vccd1 _19132_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16343_ _16343_/A vssd1 vssd1 vccd1 vccd1 _22338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13555_ _13555_/A _13555_/B vssd1 vssd1 vccd1 vccd1 _16131_/A sky130_fd_sc_hd__xnor2_4
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_319_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_346_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12506_ _12506_/A _12506_/B vssd1 vssd1 vccd1 vccd1 _12506_/X sky130_fd_sc_hd__or2_1
X_19062_ _16876_/X _23224_/Q _19062_/S vssd1 vssd1 vccd1 vccd1 _19063_/A sky130_fd_sc_hd__mux2_1
X_16274_ _16274_/A vssd1 vssd1 vccd1 vccd1 _22313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_347_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ _14206_/A _13655_/A vssd1 vssd1 vccd1 vccd1 _14220_/A sky130_fd_sc_hd__and2_4
XFILLER_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18013_ _18009_/C _17894_/X _18009_/X _18011_/X _18012_/X vssd1 vssd1 vccd1 vccd1
+ _22845_/D sky130_fd_sc_hd__o2111a_1
X_15225_ _14592_/X _15209_/X _15224_/X _14748_/X vssd1 vssd1 vccd1 vccd1 _15225_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_9_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12437_ _12421_/A _12436_/X _11229_/A vssd1 vssd1 vccd1 vccd1 _12437_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_138_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput407 _22585_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_ack_o sky130_fd_sc_hd__buf_2
XFILLER_315_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15156_ _14520_/A _15124_/X _15139_/Y _15155_/X _14587_/X vssd1 vssd1 vccd1 vccd1
+ _15156_/X sky130_fd_sc_hd__a32o_1
XFILLER_314_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput418 _22572_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[19] sky130_fd_sc_hd__buf_2
XFILLER_299_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12368_ _13763_/A _12368_/B _13714_/B vssd1 vssd1 vccd1 vccd1 _12368_/X sky130_fd_sc_hd__and3_1
Xoutput429 _22582_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[29] sky130_fd_sc_hd__buf_2
XFILLER_330_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_299_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14107_ _18166_/B vssd1 vssd1 vccd1 vccd1 _14107_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_287_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11319_ _12777_/A vssd1 vssd1 vccd1 vccd1 _11320_/A sky130_fd_sc_hd__buf_4
X_19964_ _19976_/B _19960_/B _19963_/Y vssd1 vssd1 vccd1 vccd1 _23603_/D sky130_fd_sc_hd__o21a_1
X_15087_ _15086_/Y _14781_/X _15133_/A vssd1 vssd1 vccd1 vccd1 _15087_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12299_ _22782_/Q _22750_/Q _22651_/Q _22718_/Q _12242_/S _11611_/A vssd1 vssd1 vccd1
+ vccd1 _12299_/X sky130_fd_sc_hd__mux4_2
XFILLER_80_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18915_ _18915_/A vssd1 vssd1 vccd1 vccd1 _23158_/D sky130_fd_sc_hd__clkbuf_1
X_14038_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14038_/X sky130_fd_sc_hd__buf_2
XTAP_7080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19895_ _19895_/A vssd1 vssd1 vccd1 vccd1 _23579_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_312_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18846_ _18846_/A vssd1 vssd1 vccd1 vccd1 _18846_/X sky130_fd_sc_hd__clkbuf_2
XTAP_6390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18777_ _23110_/Q _18776_/X _18786_/S vssd1 vssd1 vccd1 vccd1 _18778_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15989_ _23839_/Q _15593_/X _15985_/X _15988_/X _14923_/X vssd1 vssd1 vccd1 vccd1
+ _15989_/X sky130_fd_sc_hd__a221o_1
XFILLER_103_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17728_ _22743_/Q _17642_/X _17730_/S vssd1 vssd1 vccd1 vccd1 _17729_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17659_ _19771_/A vssd1 vssd1 vccd1 vccd1 _19555_/B sky130_fd_sc_hd__buf_8
XFILLER_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20670_ _17149_/A _20642_/X _20649_/X vssd1 vssd1 vccd1 vccd1 _20670_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_338_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19329_ _19252_/X _23328_/Q _19333_/S vssd1 vssd1 vccd1 vccd1 _19330_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_338_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_337_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22340_ _23572_/CLK _22340_/D vssd1 vssd1 vccd1 vccd1 _22340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22271_ _23503_/CLK _22271_/D vssd1 vssd1 vccd1 vccd1 _22271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21222_ _14548_/X _15121_/X _21257_/S vssd1 vssd1 vccd1 vccd1 _21223_/B sky130_fd_sc_hd__mux2_1
XFILLER_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_333_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21153_ _21153_/A _21177_/B vssd1 vssd1 vccd1 vccd1 _21153_/Y sky130_fd_sc_hd__nor2_1
XFILLER_321_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20104_ _23641_/Q _20106_/A _23642_/Q vssd1 vssd1 vccd1 vccd1 _20107_/B sky130_fd_sc_hd__a21oi_1
XFILLER_59_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21084_ _21084_/A _21084_/B vssd1 vssd1 vccd1 vccd1 _21085_/B sky130_fd_sc_hd__nor2_1
XFILLER_293_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20035_ _20041_/A _20035_/B _20048_/C vssd1 vssd1 vccd1 vccd1 _23622_/D sky130_fd_sc_hd__nor3_1
XFILLER_258_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_301_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21986_ _21999_/A _21845_/A _21985_/X _21847_/A vssd1 vssd1 vccd1 vccd1 _22041_/C
+ sky130_fd_sc_hd__o22a_2
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_328_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23725_ _23755_/CLK _23725_/D vssd1 vssd1 vccd1 vccd1 _23725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20937_ _17133_/X _20936_/X _20665_/B _20926_/X vssd1 vssd1 vccd1 vccd1 _20937_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _22374_/Q _22406_/Q _22695_/Q _23062_/Q _12716_/A _11669_/X vssd1 vssd1 vccd1
+ vccd1 _11670_/X sky130_fd_sc_hd__mux4_1
X_23656_ _23818_/CLK _23656_/D vssd1 vssd1 vccd1 vccd1 _23656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20868_ _20868_/A vssd1 vssd1 vccd1 vccd1 _23773_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22607_ _23646_/CLK _22607_/D vssd1 vssd1 vccd1 vccd1 _22607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23587_ _23893_/CLK _23587_/D vssd1 vssd1 vccd1 vccd1 _23587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_356_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20799_ _20608_/B _20791_/X _20792_/X _23755_/Q vssd1 vssd1 vccd1 vccd1 _20800_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13340_ _13340_/A _13340_/B vssd1 vssd1 vccd1 vccd1 _13375_/B sky130_fd_sc_hd__nor2_1
X_22538_ _23572_/CLK _22538_/D vssd1 vssd1 vccd1 vccd1 _22538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_316_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13271_ _13264_/Y _13266_/Y _13268_/Y _13270_/Y _11247_/X vssd1 vssd1 vccd1 vccd1
+ _13271_/X sky130_fd_sc_hd__o221a_1
XFILLER_154_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_343_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_294_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22469_ _22632_/CLK _22469_/D vssd1 vssd1 vccd1 vccd1 _22469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_129_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23602_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_185_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15010_ _15010_/A _15010_/B vssd1 vssd1 vccd1 vccd1 _15010_/Y sky130_fd_sc_hd__nor2_1
X_12222_ _23212_/Q _23180_/Q _23148_/Q _23116_/Q _12215_/X _12216_/X vssd1 vssd1 vccd1
+ vccd1 _12222_/X sky130_fd_sc_hd__mux4_2
XFILLER_151_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12153_ _22466_/Q _22626_/Q _22305_/Q _23441_/Q _11741_/X _12025_/A vssd1 vssd1 vccd1
+ vccd1 _12153_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_335_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11104_ _23891_/Q vssd1 vssd1 vccd1 vccd1 _13470_/A sky130_fd_sc_hd__buf_2
XFILLER_297_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16961_ _11069_/D _16957_/X _17317_/S vssd1 vssd1 vccd1 vccd1 _16961_/X sky130_fd_sc_hd__mux2_1
X_12084_ _11582_/A _12083_/X _11230_/A vssd1 vssd1 vccd1 vccd1 _12084_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_311_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18700_ _16813_/X _23077_/Q _18708_/S vssd1 vssd1 vccd1 vccd1 _18701_/A sky130_fd_sc_hd__mux2_1
X_15912_ _22970_/Q _15911_/X _15982_/B vssd1 vssd1 vccd1 vccd1 _15912_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19680_ _19239_/X _23484_/Q _19682_/S vssd1 vssd1 vccd1 vccd1 _19681_/A sky130_fd_sc_hd__mux2_1
X_16892_ _19242_/A vssd1 vssd1 vccd1 vccd1 _16892_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_249_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18631_ _18631_/A vssd1 vssd1 vccd1 vccd1 _23046_/D sky130_fd_sc_hd__clkbuf_1
X_15843_ _14516_/A _15836_/X _15842_/Y _15652_/X vssd1 vssd1 vccd1 vccd1 _15844_/B
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18562_ _16825_/X _23016_/Q _18564_/S vssd1 vssd1 vccd1 vccd1 _18563_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12986_ _11233_/A _12983_/X _12985_/X _11559_/X vssd1 vssd1 vccd1 vccd1 _12986_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15774_ _14586_/A _15767_/X _15773_/X _14690_/A vssd1 vssd1 vccd1 vccd1 _15775_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ _17513_/A vssd1 vssd1 vccd1 vccd1 _22663_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_280_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14725_ _14725_/A _15287_/A vssd1 vssd1 vccd1 vccd1 _14725_/X sky130_fd_sc_hd__or2_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18493_ _18480_/X _18492_/Y _18490_/X vssd1 vssd1 vccd1 vccd1 _22992_/D sky130_fd_sc_hd__a21oi_1
XFILLER_261_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11937_ _13518_/A _13340_/A _13340_/B vssd1 vssd1 vccd1 vccd1 _11937_/X sky130_fd_sc_hd__or3_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17444_ _17444_/A vssd1 vssd1 vccd1 vccd1 _22633_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14656_ _14327_/X _14329_/X _14660_/S vssd1 vssd1 vccd1 vccd1 _14656_/X sky130_fd_sc_hd__mux2_1
X_11868_ _11348_/A _11861_/Y _11863_/Y _11865_/Y _11867_/Y vssd1 vssd1 vccd1 vccd1
+ _11868_/X sky130_fd_sc_hd__o32a_1
XFILLER_300_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13607_ _15582_/A _13612_/A vssd1 vssd1 vccd1 vccd1 _13608_/B sky130_fd_sc_hd__nor2_2
XFILLER_300_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17375_ _17375_/A vssd1 vssd1 vccd1 vccd1 _22607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14587_ _15815_/A vssd1 vssd1 vccd1 vccd1 _14587_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11799_ _11799_/A vssd1 vssd1 vccd1 vccd1 _11799_/X sky130_fd_sc_hd__buf_4
XFILLER_159_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19114_ _19114_/A vssd1 vssd1 vccd1 vccd1 _23246_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16326_ _16326_/A vssd1 vssd1 vccd1 vccd1 _22330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_319_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13538_ _15678_/A _13538_/B vssd1 vssd1 vccd1 vccd1 _13538_/X sky130_fd_sc_hd__or2_1
XFILLER_185_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19045_ _16851_/X _23216_/Q _19051_/S vssd1 vssd1 vccd1 vccd1 _19046_/A sky130_fd_sc_hd__mux2_1
X_16257_ _22308_/Q _16255_/X _16269_/S vssd1 vssd1 vccd1 vccd1 _16258_/A sky130_fd_sc_hd__mux2_1
X_13469_ _14216_/A _14216_/B vssd1 vssd1 vccd1 vccd1 _13879_/B sky130_fd_sc_hd__nand2_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15208_ _23597_/Q vssd1 vssd1 vccd1 vccd1 _19975_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_309_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_350_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16188_ _16188_/A _16188_/B vssd1 vssd1 vccd1 vccd1 _16188_/Y sky130_fd_sc_hd__nand2_1
XFILLER_316_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_315_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15139_ _15139_/A _15139_/B vssd1 vssd1 vccd1 vccd1 _15139_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_287_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_331_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19947_ _19950_/A _19953_/C vssd1 vssd1 vccd1 vccd1 _19947_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_330_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19878_ _19900_/A vssd1 vssd1 vccd1 vccd1 _19887_/S sky130_fd_sc_hd__buf_6
XFILLER_110_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18829_ _18829_/A vssd1 vssd1 vccd1 vccd1 _23126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21840_ _21840_/A vssd1 vssd1 vccd1 vccd1 _21847_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_270_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21771_ _21771_/A _21865_/A vssd1 vssd1 vccd1 vccd1 _21771_/X sky130_fd_sc_hd__or2_1
XFILLER_36_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23510_ _23510_/CLK _23510_/D vssd1 vssd1 vccd1 vccd1 _23510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20722_ _23740_/Q _20697_/X _20721_/X _20706_/X vssd1 vssd1 vccd1 vccd1 _23740_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_357_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23441_ _23441_/CLK _23441_/D vssd1 vssd1 vccd1 vccd1 _23441_/Q sky130_fd_sc_hd__dfxtp_1
X_20653_ _23729_/Q _20628_/X _20652_/X _20637_/X vssd1 vssd1 vccd1 vccd1 _23729_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_338_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23372_ _23950_/A _23372_/D vssd1 vssd1 vccd1 vccd1 _23372_/Q sky130_fd_sc_hd__dfxtp_1
X_20584_ _23720_/Q _20542_/X _20583_/X _20559_/X vssd1 vssd1 vccd1 vccd1 _23720_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_353_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_358_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22323_ _23893_/CLK _22323_/D vssd1 vssd1 vccd1 vccd1 _22323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_307_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22254_ _22254_/A _22254_/B vssd1 vssd1 vccd1 vccd1 _22255_/A sky130_fd_sc_hd__and2_1
XFILLER_164_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21205_ _11069_/C _21202_/X _21204_/Y _21186_/X vssd1 vssd1 vccd1 vccd1 _23880_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_254_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22185_ _23842_/Q _23776_/Q vssd1 vssd1 vccd1 vccd1 _22187_/A sky130_fd_sc_hd__or2_1
XFILLER_155_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21136_ _23862_/Q _21135_/X _21124_/A _21033_/A vssd1 vssd1 vccd1 vccd1 _21137_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21067_ _20749_/A _21047_/X _21066_/X _21061_/X vssd1 vssd1 vccd1 vccd1 _23841_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20018_ _23617_/Q _20026_/C _20017_/Y vssd1 vssd1 vccd1 vccd1 _23617_/D sky130_fd_sc_hd__o21a_1
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_261_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12840_ _12816_/X _12667_/X _11402_/A _12839_/Y vssd1 vssd1 vccd1 vccd1 _13029_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_46_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12871_/A _12770_/X _11232_/A vssd1 vssd1 vccd1 vccd1 _12771_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21969_ _23834_/Q _23768_/Q vssd1 vssd1 vccd1 vccd1 _21971_/A sky130_fd_sc_hd__and2_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11722_ _22272_/Q _23088_/Q _23504_/Q _22433_/Q _12120_/S _11163_/A vssd1 vssd1 vccd1
+ vccd1 _11723_/B sky130_fd_sc_hd__mux4_1
X_14510_ _14510_/A _14510_/B vssd1 vssd1 vccd1 vccd1 _14933_/A sky130_fd_sc_hd__or2_2
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15085_/X _15083_/X _15490_/S vssd1 vssd1 vccd1 vccd1 _15490_/X sky130_fd_sc_hd__mux2_1
X_23708_ _23714_/CLK _23708_/D vssd1 vssd1 vccd1 vccd1 _23708_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23639_ _23652_/CLK _23639_/D vssd1 vssd1 vccd1 vccd1 _23639_/Q sky130_fd_sc_hd__dfxtp_1
X_11653_ _11653_/A vssd1 vssd1 vccd1 vccd1 _11676_/A sky130_fd_sc_hd__buf_2
X_14441_ _14728_/B vssd1 vssd1 vccd1 vccd1 _14868_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17160_ _17158_/X _17159_/Y _17163_/B vssd1 vssd1 vccd1 vccd1 _17160_/Y sky130_fd_sc_hd__o21ai_1
X_14372_ _14370_/X _14371_/Y _14175_/Y vssd1 vssd1 vccd1 vccd1 _15079_/B sky130_fd_sc_hd__o21a_4
X_11584_ _11584_/A vssd1 vssd1 vccd1 vccd1 _11587_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_344_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_316_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16111_ _14755_/X _16099_/X _16110_/X vssd1 vssd1 vccd1 vccd1 _17298_/A sky130_fd_sc_hd__o21ai_4
X_13323_ _13323_/A _13323_/B vssd1 vssd1 vccd1 vccd1 _13324_/B sky130_fd_sc_hd__nand2_2
X_17091_ _17091_/A vssd1 vssd1 vccd1 vccd1 _17091_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_344_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13254_ _22321_/Q _23457_/Q _13254_/S vssd1 vssd1 vccd1 vccd1 _13254_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16042_ _16004_/A _16041_/Y _14807_/A vssd1 vssd1 vccd1 vccd1 _16042_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_344_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_297_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12205_ _11911_/B _13727_/A _12204_/Y vssd1 vssd1 vccd1 vccd1 _12235_/A sky130_fd_sc_hd__a21oi_4
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_324_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13185_ _13165_/Y _20362_/A _13185_/S vssd1 vssd1 vccd1 vccd1 _13240_/A sky130_fd_sc_hd__mux2_2
XFILLER_313_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_296_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19801_ _19801_/A vssd1 vssd1 vccd1 vccd1 _23537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12136_ _13470_/A _12157_/S _11400_/A _12135_/Y vssd1 vssd1 vccd1 vccd1 _12159_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_123_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17993_ _22839_/Q _17990_/X _17986_/X _17992_/X _17983_/X vssd1 vssd1 vccd1 vccd1
+ _17993_/X sky130_fd_sc_hd__a221o_1
XFILLER_215_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19732_ _19210_/X _23507_/Q _19732_/S vssd1 vssd1 vccd1 vccd1 _19733_/A sky130_fd_sc_hd__mux2_1
X_16944_ _16944_/A _16966_/A _14147_/B vssd1 vssd1 vccd1 vccd1 _16945_/B sky130_fd_sc_hd__or3b_1
X_12067_ _22370_/Q _22402_/Q _22691_/Q _23058_/Q _11700_/X _11839_/A vssd1 vssd1 vccd1
+ vccd1 _12067_/X sky130_fd_sc_hd__mux4_1
XFILLER_284_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_97_wb_clk_i _22899_/CLK vssd1 vssd1 vccd1 vccd1 _23522_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19663_ _19213_/X _23476_/Q _19671_/S vssd1 vssd1 vccd1 vccd1 _19664_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16875_ _16875_/A vssd1 vssd1 vccd1 vccd1 _22539_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_26_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23491_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18614_ _18614_/A vssd1 vssd1 vccd1 vccd1 _23039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_265_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15826_ _15826_/A vssd1 vssd1 vccd1 vccd1 _21077_/B sky130_fd_sc_hd__buf_6
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19594_ _19594_/A vssd1 vssd1 vccd1 vccd1 _23445_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18545_ _22877_/Q _18203_/C _18542_/A _16945_/A vssd1 vssd1 vccd1 vccd1 _18545_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_206_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15757_ _23673_/Q _16137_/B vssd1 vssd1 vccd1 vccd1 _15757_/X sky130_fd_sc_hd__or2_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _23483_/Q _23579_/Q _22543_/Q _22347_/Q _12819_/S _11166_/A vssd1 vssd1 vccd1
+ vccd1 _12969_/X sky130_fd_sc_hd__mux4_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14708_ _14708_/A vssd1 vssd1 vccd1 vccd1 _22262_/D sky130_fd_sc_hd__clkbuf_1
X_18476_ _18476_/A vssd1 vssd1 vccd1 vccd1 _18476_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_221_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15688_ _23735_/Q _23865_/Q _16022_/S vssd1 vssd1 vccd1 vccd1 _15688_/X sky130_fd_sc_hd__mux2_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17427_ _17427_/A vssd1 vssd1 vccd1 vccd1 _22625_/D sky130_fd_sc_hd__clkbuf_1
X_14639_ _14639_/A vssd1 vssd1 vccd1 vccd1 _14853_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_202_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17358_ _22600_/Q input194/X _17358_/S vssd1 vssd1 vccd1 vccd1 _17359_/A sky130_fd_sc_hd__mux2_1
XFILLER_308_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16309_ _17471_/A _17471_/B _18770_/B vssd1 vssd1 vccd1 vccd1 _19843_/A sky130_fd_sc_hd__or3_1
XFILLER_146_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17289_ _17289_/A vssd1 vssd1 vccd1 vccd1 _17289_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_335_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_307_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19028_ _19028_/A vssd1 vssd1 vccd1 vccd1 _23208_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_350_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_288_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22941_ _23649_/CLK _22941_/D vssd1 vssd1 vccd1 vccd1 _22941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22872_ _23592_/CLK _22872_/D vssd1 vssd1 vccd1 vccd1 _22872_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_283_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21823_ _23829_/Q _22214_/S _21822_/Y _21634_/A vssd1 vssd1 vccd1 vccd1 _21831_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21754_ _23827_/Q _23761_/Q vssd1 vssd1 vccd1 vccd1 _21756_/A sky130_fd_sc_hd__and2_1
XPHY_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20705_ _20727_/A _20705_/B _20705_/C vssd1 vssd1 vccd1 vccd1 _20705_/X sky130_fd_sc_hd__or3_1
XFILLER_358_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21685_ _15080_/A _21556_/X _21849_/A vssd1 vssd1 vccd1 vccd1 _21725_/B sky130_fd_sc_hd__o21a_1
XFILLER_196_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23424_ _23424_/CLK _23424_/D vssd1 vssd1 vccd1 vccd1 _23424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_357_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_339_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_338_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20636_ _20963_/A vssd1 vssd1 vccd1 vccd1 _20763_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_196_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23355_ _23549_/CLK _23355_/D vssd1 vssd1 vccd1 vccd1 _23355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_338_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20567_ _21317_/A _20563_/X _20566_/X vssd1 vssd1 vccd1 vccd1 _20568_/C sky130_fd_sc_hd__o21a_1
XFILLER_20_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22306_ _23570_/CLK _22306_/D vssd1 vssd1 vccd1 vccd1 _22306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_326_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_326_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23286_ _23414_/CLK _23286_/D vssd1 vssd1 vccd1 vccd1 _23286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_307_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20498_ _21615_/A vssd1 vssd1 vccd1 vccd1 _21517_/B sky130_fd_sc_hd__buf_2
XFILLER_106_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22237_ _22235_/Y _22236_/X _16194_/X vssd1 vssd1 vccd1 vccd1 _22237_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22168_ _22168_/A vssd1 vssd1 vccd1 vccd1 _22168_/Y sky130_fd_sc_hd__inv_2
XTAP_6934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_294_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21119_ _21121_/A _21119_/B vssd1 vssd1 vccd1 vccd1 _23855_/D sky130_fd_sc_hd__nor2_1
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_293_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14990_ _23594_/Q vssd1 vssd1 vccd1 vccd1 _19934_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_22099_ _22099_/A vssd1 vssd1 vccd1 vccd1 _22101_/A sky130_fd_sc_hd__inv_2
XFILLER_59_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13941_ _16679_/B _14095_/A vssd1 vssd1 vccd1 vccd1 _13941_/Y sky130_fd_sc_hd__nor2_1
XFILLER_235_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16660_ _22477_/Q _16281_/X _16662_/S vssd1 vssd1 vccd1 vccd1 _16661_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13872_ _13967_/B _13872_/B vssd1 vssd1 vccd1 vccd1 _13873_/A sky130_fd_sc_hd__and2_1
XFILLER_262_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15611_ _21826_/A _15611_/B vssd1 vssd1 vccd1 vccd1 _15612_/B sky130_fd_sc_hd__nor2_1
X_12823_ _23228_/Q _23196_/Q _23164_/Q _23132_/Q _12680_/X _12637_/X vssd1 vssd1 vccd1
+ vccd1 _12824_/B sky130_fd_sc_hd__mux4_2
X_16591_ _16591_/A vssd1 vssd1 vccd1 vccd1 _22446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_262_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18330_ _15833_/X _18332_/C _18329_/Y vssd1 vssd1 vccd1 vccd1 _22936_/D sky130_fd_sc_hd__o21a_1
XFILLER_243_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15542_ _14671_/S _15541_/Y _15253_/X vssd1 vssd1 vccd1 vccd1 _15542_/X sky130_fd_sc_hd__a21o_1
X_12754_ _12754_/A vssd1 vssd1 vccd1 vccd1 _12871_/A sky130_fd_sc_hd__buf_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18261_ _20121_/A vssd1 vssd1 vccd1 vccd1 _18264_/A sky130_fd_sc_hd__buf_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11705_/A vssd1 vssd1 vccd1 vccd1 _11706_/A sky130_fd_sc_hd__buf_4
X_12685_ _12685_/A vssd1 vssd1 vccd1 vccd1 _12685_/X sky130_fd_sc_hd__buf_6
X_15473_ _18814_/A vssd1 vssd1 vccd1 vccd1 _19207_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_144_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _22929_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_230_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17212_ _16989_/X _15815_/B _17170_/B _23482_/Q _17202_/Y vssd1 vssd1 vccd1 vccd1
+ _17212_/X sky130_fd_sc_hd__a221o_1
X_11636_ _12091_/A vssd1 vssd1 vccd1 vccd1 _12007_/A sky130_fd_sc_hd__clkbuf_4
X_14424_ _22712_/Q _16942_/A _14551_/B vssd1 vssd1 vccd1 vccd1 _14424_/X sky130_fd_sc_hd__or3_1
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18192_ _21681_/A vssd1 vssd1 vccd1 vccd1 _18192_/X sky130_fd_sc_hd__buf_12
XFILLER_129_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_329_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_317_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17143_ input84/X input49/X _17200_/S vssd1 vssd1 vccd1 vccd1 _17143_/X sky130_fd_sc_hd__mux2_8
X_11567_ _11949_/A vssd1 vssd1 vccd1 vccd1 _11568_/A sky130_fd_sc_hd__buf_4
X_14355_ _14358_/A vssd1 vssd1 vccd1 vccd1 _14762_/A sky130_fd_sc_hd__buf_2
XFILLER_128_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_345_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13306_ _13306_/A _13306_/B vssd1 vssd1 vccd1 vccd1 _16128_/S sky130_fd_sc_hd__nor2_1
XFILLER_305_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17074_ _23469_/Q _17061_/X _17062_/X _17042_/X _15230_/X vssd1 vssd1 vccd1 vccd1
+ _17074_/X sky130_fd_sc_hd__a32o_1
XFILLER_157_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14286_ _14672_/B _11489_/B _14317_/S vssd1 vssd1 vccd1 vccd1 _14286_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11498_ _22386_/Q _22418_/Q _22707_/Q _23074_/Q _11432_/X _11435_/X vssd1 vssd1 vccd1
+ vccd1 _11498_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_344_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13237_ _13237_/A _13573_/A vssd1 vssd1 vccd1 vccd1 _13579_/A sky130_fd_sc_hd__nor2_2
X_16025_ _23840_/Q _15211_/X _16021_/X _16024_/X _15222_/X vssd1 vssd1 vccd1 vccd1
+ _16025_/X sky130_fd_sc_hd__a221o_1
XFILLER_237_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_297_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13168_ _23486_/Q _23582_/Q _22546_/Q _22350_/Q _11532_/X _11544_/A vssd1 vssd1 vccd1
+ vccd1 _13169_/B sky130_fd_sc_hd__mux4_2
XFILLER_301_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12119_ _22466_/Q _22626_/Q _12119_/S vssd1 vssd1 vccd1 vccd1 _12119_/X sky130_fd_sc_hd__mux2_1
X_17976_ _22836_/Q _17965_/X _17975_/X _17963_/X vssd1 vssd1 vccd1 vccd1 _22836_/D
+ sky130_fd_sc_hd__o211a_1
X_13099_ _11235_/A _13087_/Y _13093_/Y _13095_/Y _13098_/Y vssd1 vssd1 vccd1 vccd1
+ _13099_/X sky130_fd_sc_hd__o32a_1
XFILLER_284_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater504 _12634_/Y vssd1 vssd1 vccd1 vccd1 _20296_/A sky130_fd_sc_hd__buf_6
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19715_ _19185_/X _23499_/Q _19721_/S vssd1 vssd1 vccd1 vccd1 _19716_/A sky130_fd_sc_hd__mux2_1
X_16927_ _16927_/A _16927_/B vssd1 vssd1 vccd1 vccd1 _17237_/A sky130_fd_sc_hd__nor2_4
XFILLER_300_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_348_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19646_ _19646_/A vssd1 vssd1 vccd1 vccd1 _23468_/D sky130_fd_sc_hd__clkbuf_1
X_16858_ _16857_/X _22534_/Q _16861_/S vssd1 vssd1 vccd1 vccd1 _16859_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_309_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15809_ _23834_/Q _15211_/A _15805_/X _15808_/X _15222_/A vssd1 vssd1 vccd1 vccd1
+ _15809_/X sky130_fd_sc_hd__a221o_1
X_19577_ _23438_/Q _19194_/A _19577_/S vssd1 vssd1 vccd1 vccd1 _19578_/A sky130_fd_sc_hd__mux2_1
XFILLER_280_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16789_ _16795_/A _16789_/B vssd1 vssd1 vccd1 vccd1 _16790_/A sky130_fd_sc_hd__or2_1
XFILLER_111_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18528_ _23006_/Q _18530_/B vssd1 vssd1 vccd1 vccd1 _18528_/Y sky130_fd_sc_hd__nand2_1
XFILLER_234_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_339_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18459_ _18451_/X _18458_/Y _22260_/A vssd1 vssd1 vccd1 vccd1 _22979_/D sky130_fd_sc_hd__a21oi_1
XFILLER_178_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21470_ _21468_/Y _21470_/B vssd1 vssd1 vccd1 vccd1 _21472_/B sky130_fd_sc_hd__and2b_1
XFILLER_355_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20421_ _20570_/A _20408_/X _20419_/X _20420_/X vssd1 vssd1 vccd1 vccd1 _23687_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_335_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23140_ _23578_/CLK _23140_/D vssd1 vssd1 vccd1 vccd1 _23140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_308_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20352_ _23676_/Q _20177_/A _20351_/Y _20324_/X vssd1 vssd1 vccd1 vccd1 _23676_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_308_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23071_ _23583_/CLK _23071_/D vssd1 vssd1 vccd1 vccd1 _23071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_350_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20283_ _20344_/A vssd1 vssd1 vccd1 vccd1 _20338_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_290_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_289_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22022_ _23836_/Q _23770_/Q vssd1 vssd1 vccd1 vccd1 _22023_/B sky130_fd_sc_hd__nor2_1
XTAP_6219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_331_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_291_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22924_ _22929_/CLK _22924_/D vssd1 vssd1 vccd1 vccd1 _22924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22855_ _22908_/CLK _22855_/D vssd1 vssd1 vccd1 vccd1 _22855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21806_ _20296_/A _21870_/A _15612_/Y _22046_/A vssd1 vssd1 vccd1 vccd1 _21806_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22786_ _23054_/CLK _22786_/D vssd1 vssd1 vccd1 vccd1 _22786_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21737_ _21737_/A _21741_/A vssd1 vssd1 vccd1 vccd1 _21739_/A sky130_fd_sc_hd__nand2_1
XFILLER_358_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12470_ _11949_/A _11404_/B _12520_/S vssd1 vssd1 vccd1 vccd1 _12470_/Y sky130_fd_sc_hd__o21ai_1
X_21668_ _21627_/Y _21632_/B _21629_/B vssd1 vssd1 vccd1 vccd1 _21669_/B sky130_fd_sc_hd__o21ai_4
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11421_ _23491_/Q _23587_/Q _22551_/Q _22355_/Q _13254_/S _11418_/X vssd1 vssd1 vccd1
+ vccd1 _11421_/X sky130_fd_sc_hd__mux4_1
XFILLER_345_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20619_ _13939_/B _20563_/X _20618_/X vssd1 vssd1 vccd1 vccd1 _20620_/C sky130_fd_sc_hd__o21a_1
X_23407_ _23407_/CLK _23407_/D vssd1 vssd1 vccd1 vccd1 _23407_/Q sky130_fd_sc_hd__dfxtp_1
X_21599_ _21596_/X _21597_/X _21598_/X vssd1 vssd1 vccd1 vccd1 _21599_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_327_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14140_ _23010_/Q vssd1 vssd1 vccd1 vccd1 _18537_/B sky130_fd_sc_hd__inv_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11352_ _11352_/A vssd1 vssd1 vccd1 vccd1 _11353_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23338_ _23370_/CLK _23338_/D vssd1 vssd1 vccd1 vccd1 _23338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14071_ _14071_/A vssd1 vssd1 vccd1 vccd1 _14072_/A sky130_fd_sc_hd__buf_2
X_11283_ _11630_/A vssd1 vssd1 vccd1 vccd1 _11284_/A sky130_fd_sc_hd__clkbuf_4
X_23269_ _23397_/CLK _23269_/D vssd1 vssd1 vccd1 vccd1 _23269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ _13022_/A _13022_/B vssd1 vssd1 vccd1 vccd1 _13388_/B sky130_fd_sc_hd__nand2_1
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17830_ _17830_/A vssd1 vssd1 vccd1 vccd1 _22787_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17761_ _22757_/Q _17585_/X _17765_/S vssd1 vssd1 vccd1 vccd1 _17762_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14973_ _16004_/A vssd1 vssd1 vccd1 vccd1 _15161_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_294_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19500_ _19500_/A vssd1 vssd1 vccd1 vccd1 _23403_/D sky130_fd_sc_hd__clkbuf_1
X_16712_ _16730_/A vssd1 vssd1 vccd1 vccd1 _16712_/X sky130_fd_sc_hd__clkbuf_2
X_13924_ _14220_/A vssd1 vssd1 vccd1 vccd1 _13924_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_208_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17692_ _17692_/A vssd1 vssd1 vccd1 vccd1 _22726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19431_ _23373_/Q _18798_/X _19433_/S vssd1 vssd1 vccd1 vccd1 _19432_/A sky130_fd_sc_hd__mux2_1
X_16643_ _22469_/Q _16255_/X _16651_/S vssd1 vssd1 vccd1 vccd1 _16644_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13855_ _13855_/A _13855_/B vssd1 vssd1 vccd1 vccd1 _13856_/A sky130_fd_sc_hd__and2_1
XINSDIODE2_404 _13880_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_415 _14044_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_426 _11068_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12806_ _13599_/A _13532_/D vssd1 vssd1 vccd1 vccd1 _12806_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_437 _23911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19362_ _19362_/A vssd1 vssd1 vccd1 vccd1 _23342_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_448 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16574_ _16574_/A vssd1 vssd1 vccd1 vccd1 _22438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13786_ _13786_/A _13786_/B vssd1 vssd1 vccd1 vccd1 _13787_/A sky130_fd_sc_hd__and2_1
XINSDIODE2_459 _21220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18313_ _18314_/A _18314_/C _22931_/Q vssd1 vssd1 vccd1 vccd1 _18315_/B sky130_fd_sc_hd__a21oi_1
XFILLER_188_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15525_ _15525_/A vssd1 vssd1 vccd1 vccd1 _22275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12725_/X _12730_/X _12732_/X _12736_/X _11276_/A vssd1 vssd1 vccd1 vccd1
+ _12738_/C sky130_fd_sc_hd__a221o_1
X_19293_ _19293_/A vssd1 vssd1 vccd1 vccd1 _23311_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18244_ _22909_/Q _18253_/B vssd1 vssd1 vccd1 vccd1 _18244_/X sky130_fd_sc_hd__or2_1
XFILLER_230_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_337_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15456_ _15456_/A _15456_/B vssd1 vssd1 vccd1 vccd1 _15456_/Y sky130_fd_sc_hd__nor2_1
X_12668_ _12698_/A vssd1 vssd1 vccd1 vccd1 _12818_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14407_ _23907_/Q vssd1 vssd1 vccd1 vccd1 _21550_/A sky130_fd_sc_hd__buf_8
XFILLER_128_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11619_ _12117_/A _11619_/B vssd1 vssd1 vccd1 vccd1 _11619_/X sky130_fd_sc_hd__or2_1
X_18175_ _18423_/A vssd1 vssd1 vccd1 vccd1 _18175_/X sky130_fd_sc_hd__buf_4
X_15387_ _14859_/Y _15386_/Y _15387_/S vssd1 vssd1 vccd1 vccd1 _15387_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12599_ _14368_/A _12602_/A vssd1 vssd1 vccd1 vccd1 _12600_/B sky130_fd_sc_hd__and2_1
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17126_ _21737_/A _17125_/X _17137_/S vssd1 vssd1 vccd1 vccd1 _17126_/X sky130_fd_sc_hd__mux2_1
XFILLER_345_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14338_ _14343_/S vssd1 vssd1 vccd1 vccd1 _15171_/A sky130_fd_sc_hd__buf_2
XFILLER_171_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_333_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17057_ _17109_/A vssd1 vssd1 vccd1 vccd1 _17057_/X sky130_fd_sc_hd__clkbuf_2
X_14269_ _14281_/A vssd1 vssd1 vccd1 vccd1 _14329_/S sky130_fd_sc_hd__buf_2
XFILLER_320_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16008_ _21526_/A vssd1 vssd1 vccd1 vccd1 _21078_/A sky130_fd_sc_hd__buf_6
XFILLER_83_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_41_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23058_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ _17959_/A vssd1 vssd1 vccd1 vccd1 _17959_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_300_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20970_ _20970_/A vssd1 vssd1 vccd1 vccd1 _20970_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19629_ _19697_/S vssd1 vssd1 vccd1 vccd1 _19638_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_241_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22640_ _23583_/CLK _22640_/D vssd1 vssd1 vccd1 vccd1 _22640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_280_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22571_ _23646_/CLK _22571_/D vssd1 vssd1 vccd1 vccd1 _22571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_356_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21522_ _21522_/A _21619_/B vssd1 vssd1 vccd1 vccd1 _21522_/X sky130_fd_sc_hd__and2_1
XFILLER_355_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21453_ _21543_/B _21428_/B _21452_/X vssd1 vssd1 vccd1 vccd1 _21454_/B sky130_fd_sc_hd__a21oi_1
XFILLER_175_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20404_ _23684_/Q _20404_/B vssd1 vssd1 vccd1 vccd1 _20404_/X sky130_fd_sc_hd__or2_1
XFILLER_324_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21384_ _21520_/A _21384_/B vssd1 vssd1 vccd1 vccd1 _21384_/X sky130_fd_sc_hd__or2_1
XFILLER_107_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23123_ _23507_/CLK _23123_/D vssd1 vssd1 vccd1 vccd1 _23123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20335_ _15815_/B _20169_/X _20336_/B vssd1 vssd1 vccd1 vccd1 _20335_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_311_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23054_ _23054_/CLK _23054_/D vssd1 vssd1 vccd1 vccd1 _23054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20266_ _20275_/A vssd1 vssd1 vccd1 vccd1 _20376_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_134_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_350_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22005_ _21307_/X _21990_/X _21997_/Y _22004_/X _21410_/X vssd1 vssd1 vccd1 vccd1
+ _22005_/Y sky130_fd_sc_hd__o2111ai_2
XFILLER_115_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput104 dout0[7] vssd1 vssd1 vccd1 vccd1 input104/X sky130_fd_sc_hd__buf_2
XFILLER_298_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20197_ _11483_/X _21422_/A _20197_/S vssd1 vssd1 vccd1 vccd1 _20199_/B sky130_fd_sc_hd__mux2_1
Xinput115 dout1[17] vssd1 vssd1 vccd1 vccd1 input115/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput126 dout1[27] vssd1 vssd1 vccd1 vccd1 input126/X sky130_fd_sc_hd__clkbuf_1
XTAP_5337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput137 dout1[37] vssd1 vssd1 vccd1 vccd1 input137/X sky130_fd_sc_hd__buf_2
XFILLER_277_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput148 dout1[47] vssd1 vssd1 vccd1 vccd1 input148/X sky130_fd_sc_hd__buf_2
XTAP_5359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput159 dout1[57] vssd1 vssd1 vccd1 vccd1 input159/X sky130_fd_sc_hd__buf_2
XFILLER_276_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_292_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _23412_/Q _23028_/Q _23380_/Q _23348_/Q _12755_/A _11568_/A vssd1 vssd1 vccd1
+ vccd1 _11970_/X sky130_fd_sc_hd__mux4_2
XFILLER_229_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22907_ _22929_/CLK _22907_/D vssd1 vssd1 vccd1 vccd1 _22907_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23887_ _23888_/CLK _23887_/D vssd1 vssd1 vccd1 vccd1 _23887_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13640_ _13640_/A vssd1 vssd1 vccd1 vccd1 _17385_/B sky130_fd_sc_hd__buf_12
X_22838_ _23632_/CLK _22838_/D vssd1 vssd1 vccd1 vccd1 _22838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_260_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_346_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _13581_/A _17267_/A _13490_/A _13570_/Y vssd1 vssd1 vccd1 vccd1 _13983_/A
+ sky130_fd_sc_hd__o211a_2
X_22769_ _23451_/CLK _22769_/D vssd1 vssd1 vccd1 vccd1 _22769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15310_ _22924_/Q vssd1 vssd1 vccd1 vccd1 _18296_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _23461_/Q _23557_/Q _22521_/Q _22325_/Q _12535_/S _11609_/A vssd1 vssd1 vccd1
+ vccd1 _12523_/B sky130_fd_sc_hd__mux4_1
XFILLER_358_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16290_ _16290_/A vssd1 vssd1 vccd1 vccd1 _22318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_346_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15241_ _15240_/X _22269_/Q _15284_/S vssd1 vssd1 vccd1 vccd1 _15242_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12453_ _12465_/A _12452_/X _11843_/A vssd1 vssd1 vccd1 vccd1 _12453_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_138_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_327_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11404_ _11404_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _11910_/A sky130_fd_sc_hd__and2_1
X_15172_ _14241_/A _15109_/B _15425_/A vssd1 vssd1 vccd1 vccd1 _15172_/Y sky130_fd_sc_hd__a21oi_1
X_12384_ _23208_/Q _23176_/Q _23144_/Q _23112_/Q _11646_/A _11651_/A vssd1 vssd1 vccd1
+ vccd1 _12384_/X sky130_fd_sc_hd__mux4_1
XFILLER_338_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_299_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_338_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_342_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14123_ _22891_/Q _22890_/Q vssd1 vssd1 vccd1 vccd1 _18163_/B sky130_fd_sc_hd__or2_2
X_11335_ _13006_/A vssd1 vssd1 vccd1 vccd1 _13229_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19980_ _23607_/Q _23606_/Q _19980_/C vssd1 vssd1 vccd1 vccd1 _19988_/C sky130_fd_sc_hd__and3_1
XFILLER_193_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_330_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18931_ _18931_/A vssd1 vssd1 vccd1 vccd1 _18940_/S sky130_fd_sc_hd__buf_6
XFILLER_125_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_314_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14054_ _14049_/X _13827_/B _14041_/X input230/X vssd1 vssd1 vccd1 vccd1 _14054_/X
+ sky130_fd_sc_hd__a22o_4
X_11266_ _11404_/A _12371_/B vssd1 vssd1 vccd1 vccd1 _11267_/A sky130_fd_sc_hd__nand2_1
XFILLER_137_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13005_ _22799_/Q _22767_/Q _22668_/Q _22735_/Q _12733_/X _12734_/X vssd1 vssd1 vccd1
+ vccd1 _13006_/B sky130_fd_sc_hd__mux4_1
XTAP_7284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18862_ _18862_/A vssd1 vssd1 vccd1 vccd1 _18862_/X sky130_fd_sc_hd__clkbuf_2
XTAP_6550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11197_ _11493_/S vssd1 vssd1 vccd1 vccd1 _13254_/S sky130_fd_sc_hd__clkbuf_4
XTAP_7295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_295_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17813_ _22780_/Q _17556_/X _17815_/S vssd1 vssd1 vccd1 vccd1 _17814_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18793_ _23115_/Q _18792_/X _18802_/S vssd1 vssd1 vccd1 vccd1 _18794_/A sky130_fd_sc_hd__mux2_1
XFILLER_295_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17744_ _17744_/A vssd1 vssd1 vccd1 vccd1 _22749_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14956_ _14951_/Y _14955_/X _15341_/S vssd1 vssd1 vccd1 vccd1 _14956_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13907_ _17033_/A _13906_/Y _13931_/A vssd1 vssd1 vccd1 vccd1 _14087_/A sky130_fd_sc_hd__mux2_8
X_17675_ _17675_/A vssd1 vssd1 vccd1 vccd1 _22718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14887_ _16191_/A vssd1 vssd1 vccd1 vccd1 _15479_/A sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_201 _16808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_212 _14520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19414_ _23365_/Q _18769_/X _19422_/S vssd1 vssd1 vccd1 vccd1 _19415_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_223 _14960_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16626_ _16626_/A vssd1 vssd1 vccd1 vccd1 _22461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_290_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13838_ _13861_/A _14056_/C vssd1 vssd1 vccd1 vccd1 _13838_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_234 _15995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_245 _17103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_256 _15606_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19345_ _19345_/A vssd1 vssd1 vccd1 vccd1 _23334_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_267 _15656_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16557_ _15283_/X _22431_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _16558_/A sky130_fd_sc_hd__mux2_1
X_13769_ _14019_/C _13739_/X _13768_/Y _13746_/X vssd1 vssd1 vccd1 vccd1 _13770_/B
+ sky130_fd_sc_hd__o2bb2a_4
XINSDIODE2_278 _15767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_289 _15959_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15508_ _23763_/Q _14911_/A _14913_/A _15506_/X _15507_/X vssd1 vssd1 vccd1 vccd1
+ _15508_/X sky130_fd_sc_hd__a221o_1
X_19276_ _19175_/X _23304_/Q _19278_/S vssd1 vssd1 vccd1 vccd1 _19277_/A sky130_fd_sc_hd__mux2_1
XFILLER_338_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16488_ _16488_/A vssd1 vssd1 vccd1 vccd1 _22401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_349_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18227_ _22903_/Q _18227_/B vssd1 vssd1 vccd1 vccd1 _18227_/X sky130_fd_sc_hd__or2_1
XFILLER_31_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_337_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15439_ _22959_/Q _15501_/B vssd1 vssd1 vccd1 vccd1 _15439_/X sky130_fd_sc_hd__or2_1
XFILLER_164_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_306_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18158_ _14119_/A _22882_/Q _18158_/S vssd1 vssd1 vccd1 vccd1 _18159_/B sky130_fd_sc_hd__mux2_1
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_317_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17109_ _17109_/A vssd1 vssd1 vccd1 vccd1 _17109_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_264_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18089_ _22867_/Q _18082_/X _18083_/X _23000_/Q _18084_/X vssd1 vssd1 vccd1 vccd1
+ _18089_/X sky130_fd_sc_hd__a221o_1
XFILLER_333_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_321_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20120_ _20120_/A _20120_/B _20122_/B vssd1 vssd1 vccd1 vccd1 _23646_/D sky130_fd_sc_hd__nor3_1
XFILLER_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20051_ _20051_/A _20056_/D vssd1 vssd1 vccd1 vccd1 _20066_/C sky130_fd_sc_hd__and2_1
XFILLER_320_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23810_ _23810_/CLK _23810_/D vssd1 vssd1 vccd1 vccd1 _23810_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20953_ _20969_/A vssd1 vssd1 vccd1 vccd1 _20953_/X sky130_fd_sc_hd__clkbuf_2
X_23741_ _23874_/CLK _23741_/D vssd1 vssd1 vccd1 vccd1 _23741_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20884_ _20884_/A vssd1 vssd1 vccd1 vccd1 _23778_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23672_ _23704_/CLK _23672_/D vssd1 vssd1 vccd1 vccd1 _23672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22623_ _23566_/CLK _22623_/D vssd1 vssd1 vccd1 vccd1 _22623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_289_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22554_ _23693_/CLK _22554_/D vssd1 vssd1 vccd1 vccd1 _22554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21505_ _13471_/A _21504_/X _21465_/A vssd1 vssd1 vccd1 vccd1 _21505_/X sky130_fd_sc_hd__a21bo_1
XFILLER_195_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22485_ _23588_/CLK _22485_/D vssd1 vssd1 vccd1 vccd1 _22485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_309_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21436_ _21575_/A vssd1 vssd1 vccd1 vccd1 _22197_/B sky130_fd_sc_hd__buf_2
XFILLER_147_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21367_ _21816_/A vssd1 vssd1 vccd1 vccd1 _22025_/A sky130_fd_sc_hd__buf_2
XFILLER_351_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_352_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11120_ _12468_/B vssd1 vssd1 vccd1 vccd1 _12260_/A sky130_fd_sc_hd__buf_8
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23106_ _23554_/CLK _23106_/D vssd1 vssd1 vccd1 vccd1 _23106_/Q sky130_fd_sc_hd__dfxtp_1
X_20318_ _21900_/A _20368_/B vssd1 vssd1 vccd1 vccd1 _20318_/X sky130_fd_sc_hd__or2_1
XFILLER_123_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_311_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21298_ _21328_/A vssd1 vssd1 vccd1 vccd1 _21465_/A sky130_fd_sc_hd__buf_2
XFILLER_311_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23037_ _23547_/CLK _23037_/D vssd1 vssd1 vccd1 vccd1 _23037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_324_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20249_ _15312_/X _20169_/A _20250_/B vssd1 vssd1 vccd1 vccd1 _20249_/X sky130_fd_sc_hd__a21o_1
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _18779_/A vssd1 vssd1 vccd1 vccd1 _19172_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _23932_/Q _21950_/A _15790_/C vssd1 vssd1 vccd1 vccd1 _15828_/B sky130_fd_sc_hd__and3_1
XFILLER_264_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_291_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ _23719_/Q _23849_/Q _16171_/S vssd1 vssd1 vccd1 vccd1 _14741_/X sky130_fd_sc_hd__mux2_2
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ _11953_/A vssd1 vssd1 vccd1 vccd1 _12671_/A sky130_fd_sc_hd__buf_6
XFILLER_251_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23939_ _23942_/CLK _23939_/D vssd1 vssd1 vccd1 vccd1 _23939_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ _17460_/A vssd1 vssd1 vccd1 vccd1 _22640_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _14840_/S _14672_/B vssd1 vssd1 vccd1 vccd1 _14676_/A sky130_fd_sc_hd__nand2_1
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11884_ _21601_/A _11884_/B vssd1 vssd1 vccd1 vccd1 _11884_/Y sky130_fd_sc_hd__nand2_2
XFILLER_45_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16411_ _16411_/A vssd1 vssd1 vccd1 vccd1 _22367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13623_ _13623_/A _13623_/B vssd1 vssd1 vccd1 vccd1 _15453_/A sky130_fd_sc_hd__xnor2_4
X_17391_ _13669_/A _17012_/X _17387_/X _17390_/X vssd1 vssd1 vccd1 vccd1 _22612_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_260_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19130_ _19130_/A vssd1 vssd1 vccd1 vccd1 _23253_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_347_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16342_ _15474_/X _22338_/Q _16344_/S vssd1 vssd1 vccd1 vccd1 _16343_/A sky130_fd_sc_hd__mux2_1
XFILLER_349_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13554_ _13554_/A _13554_/B vssd1 vssd1 vccd1 vccd1 _16191_/B sky130_fd_sc_hd__xnor2_4
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19061_ _19061_/A vssd1 vssd1 vccd1 vccd1 _23223_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12505_ _23301_/Q _23269_/Q _23237_/Q _23525_/Q _12501_/X _12502_/X vssd1 vssd1 vccd1
+ vccd1 _12506_/B sky130_fd_sc_hd__mux4_1
X_16273_ _22313_/Q _16271_/X _16285_/S vssd1 vssd1 vccd1 vccd1 _16274_/A sky130_fd_sc_hd__mux2_1
X_13485_ _13779_/A _19969_/D vssd1 vssd1 vccd1 vccd1 _13655_/A sky130_fd_sc_hd__nand2_2
XFILLER_201_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18012_ _20790_/A vssd1 vssd1 vccd1 vccd1 _18012_/X sky130_fd_sc_hd__buf_12
XFILLER_201_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15224_ _23693_/Q _15210_/X _15223_/X vssd1 vssd1 vccd1 vccd1 _15224_/X sky130_fd_sc_hd__o21a_2
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_346_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12436_ _23463_/Q _23559_/Q _22523_/Q _22327_/Q _12244_/A _12292_/A vssd1 vssd1 vccd1
+ vccd1 _12436_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15155_ _14431_/X _15140_/X _15152_/X _15154_/X _14518_/X vssd1 vssd1 vccd1 vccd1
+ _15155_/X sky130_fd_sc_hd__o32a_4
Xoutput408 _22553_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[0] sky130_fd_sc_hd__buf_2
XFILLER_154_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput419 _22554_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[1] sky130_fd_sc_hd__buf_2
X_12367_ _11214_/A _12353_/X _12357_/Y _12366_/X vssd1 vssd1 vccd1 vccd1 _13714_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_181_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_314_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14106_ _18188_/A _18188_/B _22891_/Q vssd1 vssd1 vccd1 vccd1 _18166_/B sky130_fd_sc_hd__and3_2
XFILLER_99_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11318_ _11457_/B vssd1 vssd1 vccd1 vccd1 _12777_/A sky130_fd_sc_hd__clkbuf_4
X_19963_ _19976_/B _19960_/B _19962_/X vssd1 vssd1 vccd1 vccd1 _19963_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_180_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15086_ _15086_/A vssd1 vssd1 vccd1 vccd1 _15086_/Y sky130_fd_sc_hd__clkinv_2
X_12298_ _11837_/A _12295_/X _12297_/X vssd1 vssd1 vccd1 vccd1 _12298_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18914_ _23158_/Q _18827_/X _18918_/S vssd1 vssd1 vccd1 vccd1 _18915_/A sky130_fd_sc_hd__mux2_1
XFILLER_268_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11249_ _13765_/A _11249_/B _11249_/C vssd1 vssd1 vccd1 vccd1 _11249_/Y sky130_fd_sc_hd__nor3_4
X_14037_ input220/X _14027_/X _14036_/X vssd1 vssd1 vccd1 vccd1 _14037_/X sky130_fd_sc_hd__a21o_4
XTAP_7070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19894_ _16278_/X _23579_/Q _19898_/S vssd1 vssd1 vccd1 vccd1 _19895_/A sky130_fd_sc_hd__mux2_1
XTAP_7092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_295_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18845_ _18845_/A vssd1 vssd1 vccd1 vccd1 _23131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18776_ _18776_/A vssd1 vssd1 vccd1 vccd1 _18776_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15988_ _23775_/Q _15595_/X _15596_/X _15986_/X _15987_/X vssd1 vssd1 vccd1 vccd1
+ _15988_/X sky130_fd_sc_hd__a221o_2
XFILLER_243_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17727_ _17727_/A vssd1 vssd1 vccd1 vccd1 _22742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14939_ _15097_/S _14939_/B vssd1 vssd1 vccd1 vccd1 _14939_/X sky130_fd_sc_hd__or2_1
XFILLER_264_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17658_ _16940_/X _17653_/B _17655_/Y _17657_/X vssd1 vssd1 vccd1 vccd1 _22712_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_36_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16609_ _16677_/S vssd1 vssd1 vccd1 vccd1 _16618_/S sky130_fd_sc_hd__buf_4
XFILLER_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17589_ _22691_/Q _17588_/X _17592_/S vssd1 vssd1 vccd1 vccd1 _17590_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19328_ _19328_/A vssd1 vssd1 vccd1 vccd1 _23327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_338_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19259_ _19258_/X _23298_/Q _19259_/S vssd1 vssd1 vccd1 vccd1 _19260_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_337_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22270_ _23502_/CLK _22270_/D vssd1 vssd1 vccd1 vccd1 _22270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21221_ _21260_/S vssd1 vssd1 vccd1 vccd1 _21257_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_306_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_352_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_305_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_333_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21152_ _23865_/Q _21147_/X _21149_/Y _21151_/X _18192_/X vssd1 vssd1 vccd1 vccd1
+ _23865_/D sky130_fd_sc_hd__o221a_1
XFILLER_117_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20103_ _23641_/Q _20106_/A _20102_/Y vssd1 vssd1 vccd1 vccd1 _23641_/D sky130_fd_sc_hd__a21oi_1
XFILLER_259_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21083_ _21083_/A vssd1 vssd1 vccd1 vccd1 _21083_/X sky130_fd_sc_hd__buf_4
XFILLER_113_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20034_ _23620_/Q _20034_/B _20034_/C _20042_/D vssd1 vssd1 vccd1 vccd1 _20048_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_274_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21985_ _20340_/A _21870_/A _15829_/Y _21842_/A vssd1 vssd1 vccd1 vccd1 _21985_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_26_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23724_ _23755_/CLK _23724_/D vssd1 vssd1 vccd1 vccd1 _23724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ _20936_/A vssd1 vssd1 vccd1 vccd1 _20936_/X sky130_fd_sc_hd__buf_4
XFILLER_310_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_8_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_8_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_27_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23655_ _23818_/CLK _23655_/D vssd1 vssd1 vccd1 vccd1 _23655_/Q sky130_fd_sc_hd__dfxtp_1
X_20867_ _20879_/A _20867_/B vssd1 vssd1 vccd1 vccd1 _20868_/A sky130_fd_sc_hd__and2_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22606_ _23646_/CLK _22606_/D vssd1 vssd1 vccd1 vccd1 _22606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23586_ _23586_/CLK _23586_/D vssd1 vssd1 vccd1 vccd1 _23586_/Q sky130_fd_sc_hd__dfxtp_1
X_20798_ _20798_/A vssd1 vssd1 vccd1 vccd1 _23754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22537_ _23349_/CLK _22537_/D vssd1 vssd1 vccd1 vccd1 _22537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_319_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_356_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_344_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_316_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13270_ _13253_/A _13269_/X _11236_/X vssd1 vssd1 vccd1 vccd1 _13270_/Y sky130_fd_sc_hd__o21ai_1
X_22468_ _23571_/CLK _22468_/D vssd1 vssd1 vccd1 vccd1 _22468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12221_ _12383_/A _12221_/B vssd1 vssd1 vccd1 vccd1 _12221_/X sky130_fd_sc_hd__or2_1
X_21419_ _23817_/Q _21418_/A _21418_/Y _21377_/X vssd1 vssd1 vccd1 vccd1 _21419_/X
+ sky130_fd_sc_hd__o211a_2
X_22399_ _23567_/CLK _22399_/D vssd1 vssd1 vccd1 vccd1 _22399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_335_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12152_ _12780_/A _12152_/B vssd1 vssd1 vccd1 vccd1 _12152_/X sky130_fd_sc_hd__or2_1
XFILLER_151_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_169_wb_clk_i _23917_/CLK vssd1 vssd1 vccd1 vccd1 _23876_/CLK sky130_fd_sc_hd__clkbuf_16
X_11103_ _23893_/Q vssd1 vssd1 vccd1 vccd1 _14176_/A sky130_fd_sc_hd__buf_2
XFILLER_151_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_300_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16960_ _17248_/A vssd1 vssd1 vccd1 vccd1 _17317_/S sky130_fd_sc_hd__clkbuf_2
X_12083_ _23474_/Q _23570_/Q _22534_/Q _22338_/Q _11894_/S _11566_/A vssd1 vssd1 vccd1
+ vccd1 _12083_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15911_ _14730_/A _15904_/X _15910_/X _14748_/A vssd1 vssd1 vccd1 vccd1 _15911_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_277_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16891_ _16891_/A vssd1 vssd1 vccd1 vccd1 _22544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18630_ _23046_/Q _17550_/X _18636_/S vssd1 vssd1 vccd1 vccd1 _18631_/A sky130_fd_sc_hd__mux2_1
XFILLER_292_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15842_ _23707_/Q _14905_/X _15841_/X vssd1 vssd1 vccd1 vccd1 _15842_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_264_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_351_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ _18561_/A vssd1 vssd1 vccd1 vccd1 _23015_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _15801_/A _15341_/X _15769_/Y _15772_/X vssd1 vssd1 vccd1 vccd1 _15773_/X
+ sky130_fd_sc_hd__o211a_2
X_12985_ _12985_/A _12985_/B vssd1 vssd1 vccd1 vccd1 _12985_/X sky130_fd_sc_hd__or2_1
XFILLER_264_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ _22663_/Q _16262_/X _17516_/S vssd1 vssd1 vccd1 vccd1 _17513_/A sky130_fd_sc_hd__mux2_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _14724_/A _14724_/B vssd1 vssd1 vccd1 vccd1 _15287_/A sky130_fd_sc_hd__nand2_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18492_ _22992_/Q _18492_/B vssd1 vssd1 vccd1 vccd1 _18492_/Y sky130_fd_sc_hd__nand2_1
XFILLER_261_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ _12913_/S _20234_/A _11935_/X vssd1 vssd1 vccd1 vccd1 _13340_/B sky130_fd_sc_hd__a21bo_4
XFILLER_73_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17443_ _22633_/Q _16268_/X _17443_/S vssd1 vssd1 vccd1 vccd1 _17444_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14655_ _14653_/Y _14654_/X _14845_/S vssd1 vssd1 vccd1 vccd1 _14655_/X sky130_fd_sc_hd__mux2_2
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _12097_/A _11866_/X _11680_/A vssd1 vssd1 vccd1 vccd1 _11867_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_220_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13606_ _12893_/Y _13603_/X _13605_/Y _13451_/A vssd1 vssd1 vccd1 vccd1 _13974_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_319_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17374_ _22607_/Q _14148_/B _17380_/S vssd1 vssd1 vccd1 vccd1 _17375_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14586_ _14586_/A vssd1 vssd1 vccd1 vccd1 _15815_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11798_ _12324_/A vssd1 vssd1 vccd1 vccd1 _11799_/A sky130_fd_sc_hd__buf_6
XFILLER_9_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19113_ _23246_/Q _18801_/X _19113_/S vssd1 vssd1 vccd1 vccd1 _19114_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16325_ _15044_/X _22330_/Q _16333_/S vssd1 vssd1 vccd1 vccd1 _16326_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13537_ _13535_/Y _15582_/A _13536_/Y vssd1 vssd1 vccd1 vccd1 _13538_/B sky130_fd_sc_hd__o21a_1
XFILLER_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_319_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19044_ _19044_/A vssd1 vssd1 vccd1 vccd1 _23215_/D sky130_fd_sc_hd__clkbuf_1
X_16256_ _16288_/A vssd1 vssd1 vccd1 vccd1 _16269_/S sky130_fd_sc_hd__buf_4
X_13468_ _13367_/C _13593_/A _13587_/A _23911_/Q vssd1 vssd1 vccd1 vccd1 _14216_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15207_ _22954_/Q vssd1 vssd1 vccd1 vccd1 _15207_/X sky130_fd_sc_hd__buf_2
X_12419_ _12570_/A _12419_/B vssd1 vssd1 vccd1 vccd1 _12419_/Y sky130_fd_sc_hd__nor2_1
X_16187_ _14586_/A _16179_/X _16186_/X vssd1 vssd1 vccd1 vccd1 _16188_/B sky130_fd_sc_hd__a21o_1
X_13399_ _13399_/A _13399_/B vssd1 vssd1 vccd1 vccd1 _13399_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_331_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15138_ _14632_/A _15915_/B _15137_/X _14839_/X vssd1 vssd1 vccd1 vccd1 _15139_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_315_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_288_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_331_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_303_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19946_ _23598_/Q _19975_/D _19971_/B vssd1 vssd1 vccd1 vccd1 _19953_/C sky130_fd_sc_hd__and3_1
X_15069_ _23723_/Q _23853_/Q _16171_/S vssd1 vssd1 vccd1 vccd1 _15069_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19877_ _19877_/A vssd1 vssd1 vccd1 vccd1 _23571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_295_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18828_ _23126_/Q _18827_/X _18834_/S vssd1 vssd1 vccd1 vccd1 _18829_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18759_ _16902_/X _23104_/Q _18763_/S vssd1 vssd1 vccd1 vccd1 _18760_/A sky130_fd_sc_hd__mux2_1
XFILLER_270_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21770_ _17133_/X _21612_/X _21769_/Y _21581_/X vssd1 vssd1 vccd1 vccd1 _23925_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20721_ _20727_/A _20721_/B _20721_/C vssd1 vssd1 vccd1 vccd1 _20721_/X sky130_fd_sc_hd__or3_1
XFILLER_251_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23440_ _23440_/CLK _23440_/D vssd1 vssd1 vccd1 vccd1 _23440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20652_ _20665_/A _20652_/B _20652_/C vssd1 vssd1 vccd1 vccd1 _20652_/X sky130_fd_sc_hd__or3_1
XFILLER_17_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23371_ _23531_/CLK _23371_/D vssd1 vssd1 vccd1 vccd1 _23371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20583_ _20591_/A _20583_/B _20583_/C vssd1 vssd1 vccd1 vccd1 _20583_/X sky130_fd_sc_hd__or3_1
XFILLER_104_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22322_ _23586_/CLK _22322_/D vssd1 vssd1 vccd1 vccd1 _22322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22253_ _23944_/Q _20536_/B _22253_/S vssd1 vssd1 vccd1 vccd1 _22254_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_opt_3_0_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21204_ _21204_/A _21227_/B vssd1 vssd1 vccd1 vccd1 _21204_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22184_ _23810_/Q _21746_/X _22183_/X _21395_/X vssd1 vssd1 vccd1 vccd1 _22184_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_333_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21135_ _21161_/A vssd1 vssd1 vccd1 vccd1 _21135_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21066_ _23841_/Q _21068_/B vssd1 vssd1 vccd1 vccd1 _21066_/X sky130_fd_sc_hd__or2_1
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20017_ _23617_/Q _20026_/C _19962_/X vssd1 vssd1 vccd1 vccd1 _20017_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_171_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _23479_/Q _23575_/Q _22539_/Q _22343_/Q _12920_/A _12746_/X vssd1 vssd1 vccd1
+ vccd1 _12770_/X sky130_fd_sc_hd__mux4_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21968_ _21944_/X _21947_/B _21945_/A vssd1 vssd1 vccd1 vccd1 _21972_/A sky130_fd_sc_hd__a21oi_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _11698_/A _11720_/X _11713_/X vssd1 vssd1 vccd1 vccd1 _11721_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23707_ _23714_/CLK _23707_/D vssd1 vssd1 vccd1 vccd1 _23707_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20919_ _13939_/B _20908_/X _20620_/B _20912_/X vssd1 vssd1 vccd1 vccd1 _20919_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21899_ _21899_/A _22044_/A vssd1 vssd1 vccd1 vccd1 _21899_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _16168_/B vssd1 vssd1 vccd1 vccd1 _14728_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_187_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23638_ _23652_/CLK _23638_/D vssd1 vssd1 vccd1 vccd1 _23638_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11652_/A vssd1 vssd1 vccd1 vccd1 _11653_/A sky130_fd_sc_hd__buf_8
XFILLER_302_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_357_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14371_ _14371_/A _14371_/B _20214_/A vssd1 vssd1 vccd1 vccd1 _14371_/Y sky130_fd_sc_hd__nor3_4
X_11583_ _11957_/A vssd1 vssd1 vccd1 vccd1 _12698_/A sky130_fd_sc_hd__clkbuf_4
X_23569_ _23571_/CLK _23569_/D vssd1 vssd1 vccd1 vccd1 _23569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16110_ _22943_/Q _14988_/B _16100_/X _16109_/Y _14898_/A vssd1 vssd1 vccd1 vccd1
+ _16110_/X sky130_fd_sc_hd__a221o_1
XFILLER_210_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_344_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13322_ _13605_/A _13329_/A _13322_/C vssd1 vssd1 vccd1 vccd1 _13323_/A sky130_fd_sc_hd__nand3_2
X_17090_ _22562_/Q _17038_/X _17083_/X _17089_/X vssd1 vssd1 vccd1 vccd1 _22562_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_182_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_344_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16041_ _16077_/B _16041_/B vssd1 vssd1 vccd1 vccd1 _16041_/Y sky130_fd_sc_hd__nor2_2
XFILLER_109_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13253_ _13253_/A _13253_/B vssd1 vssd1 vccd1 vccd1 _13253_/Y sky130_fd_sc_hd__nor2_1
XFILLER_313_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12204_ _23906_/Q _11911_/B _12415_/S vssd1 vssd1 vccd1 vccd1 _12204_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_312_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13184_ _13184_/A _13184_/B _13184_/C vssd1 vssd1 vccd1 vccd1 _20362_/A sky130_fd_sc_hd__nand3_4
XFILLER_151_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_297_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19800_ _23537_/Q _19204_/A _19804_/S vssd1 vssd1 vccd1 vccd1 _19801_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12135_ _12135_/A _13858_/A vssd1 vssd1 vccd1 vccd1 _12135_/Y sky130_fd_sc_hd__nand2_1
X_17992_ input4/X input270/X _18005_/S vssd1 vssd1 vccd1 vccd1 _17992_/X sky130_fd_sc_hd__mux2_1
XFILLER_313_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_296_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_313_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16943_ _16935_/B _22249_/C _16943_/C _17145_/A vssd1 vssd1 vccd1 vccd1 _17648_/C
+ sky130_fd_sc_hd__and4b_1
X_19731_ _19731_/A vssd1 vssd1 vccd1 vccd1 _23506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_278_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12066_ _23218_/Q _23186_/Q _23154_/Q _23122_/Q _11972_/A _11949_/A vssd1 vssd1 vccd1
+ vccd1 _12066_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16874_ _16873_/X _22539_/Q _16877_/S vssd1 vssd1 vccd1 vccd1 _16875_/A sky130_fd_sc_hd__mux2_1
X_19662_ _19684_/A vssd1 vssd1 vccd1 vccd1 _19671_/S sky130_fd_sc_hd__buf_6
XFILLER_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18613_ _16899_/X _23039_/Q _18619_/S vssd1 vssd1 vccd1 vccd1 _18614_/A sky130_fd_sc_hd__mux2_1
X_15825_ _15825_/A vssd1 vssd1 vccd1 vccd1 _22282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19593_ _23445_/Q _19217_/A _19599_/S vssd1 vssd1 vccd1 vccd1 _19594_/A sky130_fd_sc_hd__mux2_1
XFILLER_253_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _23609_/Q _14901_/A _14902_/A _23641_/Q vssd1 vssd1 vccd1 vccd1 _15756_/X
+ sky130_fd_sc_hd__o22a_4
X_18544_ _20134_/A _18544_/B vssd1 vssd1 vccd1 vccd1 _23010_/D sky130_fd_sc_hd__nor2_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12968_ _12968_/A _12968_/B vssd1 vssd1 vccd1 vccd1 _12968_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_66_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23544_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ _14706_/X _22262_/Q _14985_/S vssd1 vssd1 vccd1 vccd1 _14708_/A sky130_fd_sc_hd__mux2_1
X_18475_ _22986_/Q _18478_/B vssd1 vssd1 vccd1 vccd1 _18475_/Y sky130_fd_sc_hd__nand2_1
X_11919_ _11919_/A vssd1 vssd1 vccd1 vccd1 _11920_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15687_ _23671_/Q _16021_/B vssd1 vssd1 vccd1 vccd1 _15687_/X sky130_fd_sc_hd__or2_1
X_12899_ _22475_/Q _22635_/Q _22314_/Q _23450_/Q _12733_/A _12844_/A vssd1 vssd1 vccd1
+ vccd1 _12900_/B sky130_fd_sc_hd__mux4_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _22625_/Q _16243_/X _17432_/S vssd1 vssd1 vccd1 vccd1 _17427_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14638_ _14309_/X _14268_/X _14646_/S vssd1 vssd1 vccd1 vccd1 _14638_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17357_ _17357_/A vssd1 vssd1 vccd1 vccd1 _22599_/D sky130_fd_sc_hd__clkbuf_1
X_14569_ _14569_/A vssd1 vssd1 vccd1 vccd1 _15676_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_202_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16308_ _16308_/A vssd1 vssd1 vccd1 vccd1 _22324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17288_ _22165_/A vssd1 vssd1 vccd1 vccd1 _22166_/A sky130_fd_sc_hd__buf_8
XFILLER_174_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19027_ _16825_/X _23208_/Q _19029_/S vssd1 vssd1 vccd1 vccd1 _19028_/A sky130_fd_sc_hd__mux2_1
X_16239_ _18804_/A vssd1 vssd1 vccd1 vccd1 _16239_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_288_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_318_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19929_ _19934_/C _19929_/B vssd1 vssd1 vccd1 vccd1 _23593_/D sky130_fd_sc_hd__nor2_1
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22940_ _23649_/CLK _22940_/D vssd1 vssd1 vccd1 vccd1 _22940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_290_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22871_ _23592_/CLK _22871_/D vssd1 vssd1 vccd1 vccd1 _22871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21822_ _22242_/B _21822_/B vssd1 vssd1 vccd1 vccd1 _21822_/Y sky130_fd_sc_hd__nand2_1
XFILLER_325_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21753_ _23795_/Q _21746_/X _21752_/Y _21660_/X vssd1 vssd1 vccd1 vccd1 _21753_/X
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20704_ _15753_/A _20701_/X _20703_/Y vssd1 vssd1 vccd1 vccd1 _20705_/C sky130_fd_sc_hd__a21oi_2
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21684_ _21925_/A _21842_/A _21840_/A vssd1 vssd1 vccd1 vccd1 _21849_/A sky130_fd_sc_hd__a21o_2
XFILLER_357_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23423_ _23423_/CLK _23423_/D vssd1 vssd1 vccd1 vccd1 _23423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20635_ _20665_/A _20635_/B _20635_/C vssd1 vssd1 vccd1 vccd1 _20635_/X sky130_fd_sc_hd__or3_1
XFILLER_133_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_338_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_326_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23354_ _23354_/CLK _23354_/D vssd1 vssd1 vccd1 vccd1 _23354_/Q sky130_fd_sc_hd__dfxtp_1
X_20566_ _11069_/C _20564_/X _20732_/A vssd1 vssd1 vccd1 vccd1 _20566_/X sky130_fd_sc_hd__a21o_1
XFILLER_353_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22305_ _23568_/CLK _22305_/D vssd1 vssd1 vccd1 vccd1 _22305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23285_ _23541_/CLK _23285_/D vssd1 vssd1 vccd1 vccd1 _23285_/Q sky130_fd_sc_hd__dfxtp_1
X_20497_ _21482_/A vssd1 vssd1 vccd1 vccd1 _21615_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22236_ _17315_/X _22218_/A _22223_/A _21676_/B vssd1 vssd1 vccd1 vccd1 _22236_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22167_ _22167_/A _22166_/Y vssd1 vssd1 vccd1 vccd1 _22170_/A sky130_fd_sc_hd__or2b_1
XTAP_6924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21118_ _23855_/Q _21110_/X _21111_/X _20616_/A vssd1 vssd1 vccd1 vccd1 _21119_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_6957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_294_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22098_ _22098_/A _22100_/B vssd1 vssd1 vccd1 vccd1 _22099_/A sky130_fd_sc_hd__nand2_1
XFILLER_121_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_332_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21049_ _21163_/A vssd1 vssd1 vccd1 vccd1 _21049_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13940_ _13918_/X _13936_/X _13939_/Y _13924_/X vssd1 vssd1 vccd1 vccd1 _14095_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_208_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13871_ _13871_/A _13871_/B vssd1 vssd1 vccd1 vccd1 _13872_/B sky130_fd_sc_hd__nor2_4
XFILLER_47_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15610_ _21826_/A _15611_/B vssd1 vssd1 vccd1 vccd1 _15701_/C sky130_fd_sc_hd__and2_2
XFILLER_62_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12822_ _13195_/A _12819_/X _12821_/X vssd1 vssd1 vccd1 vccd1 _12822_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16590_ _15936_/X _22446_/Q _16590_/S vssd1 vssd1 vccd1 vccd1 _16591_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15541_ _15541_/A vssd1 vssd1 vccd1 vccd1 _15541_/Y sky130_fd_sc_hd__inv_2
X_12753_ _12749_/X _12750_/X _12752_/X vssd1 vssd1 vccd1 vccd1 _12753_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _20067_/A vssd1 vssd1 vccd1 vccd1 _20121_/A sky130_fd_sc_hd__clkbuf_4
X_11704_ _22368_/Q _22400_/Q _22689_/Q _23056_/Q _11700_/X _11839_/A vssd1 vssd1 vccd1
+ vccd1 _11704_/X sky130_fd_sc_hd__mux4_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15472_ _15470_/X _21741_/A _15708_/S vssd1 vssd1 vccd1 vccd1 _18814_/A sky130_fd_sc_hd__mux2_8
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12684_ _12978_/S vssd1 vssd1 vccd1 vccd1 _12977_/S sky130_fd_sc_hd__buf_6
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _23932_/Q vssd1 vssd1 vccd1 vccd1 _21975_/A sky130_fd_sc_hd__clkbuf_16
X_14423_ _22901_/Q _14394_/A _14164_/A _22594_/Q vssd1 vssd1 vccd1 vccd1 _14551_/B
+ sky130_fd_sc_hd__a22o_1
X_18191_ _18191_/A _18191_/B _18191_/C _18191_/D vssd1 vssd1 vccd1 vccd1 _18191_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_230_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11635_ _12401_/A vssd1 vssd1 vccd1 vccd1 _12091_/A sky130_fd_sc_hd__buf_4
XFILLER_357_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17142_ _17276_/A vssd1 vssd1 vccd1 vccd1 _17200_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_357_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14354_ _14354_/A _14840_/S vssd1 vssd1 vccd1 vccd1 _14354_/X sky130_fd_sc_hd__or2b_1
XFILLER_317_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11566_ _11566_/A vssd1 vssd1 vccd1 vccd1 _11949_/A sky130_fd_sc_hd__buf_6
XFILLER_156_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_184_wb_clk_i clkbuf_opt_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23926_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13305_ _13306_/A _13306_/B vssd1 vssd1 vccd1 vccd1 _13307_/A sky130_fd_sc_hd__and2_1
XFILLER_345_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_305_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17073_ _17073_/A vssd1 vssd1 vccd1 vccd1 _17073_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_344_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14285_ _14282_/X _14283_/X _14646_/S vssd1 vssd1 vccd1 vccd1 _14285_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11497_ _11497_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _11497_/Y sky130_fd_sc_hd__nor2_1
XFILLER_183_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_113_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23327_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16024_ _23776_/Q _15215_/X _15216_/X _16022_/X _16023_/X vssd1 vssd1 vccd1 vccd1
+ _16024_/X sky130_fd_sc_hd__a221o_4
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13236_ _13242_/A _13241_/A vssd1 vssd1 vccd1 vccd1 _13573_/A sky130_fd_sc_hd__nor2_1
XFILLER_109_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_298_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13167_ _13216_/A _13167_/B vssd1 vssd1 vccd1 vccd1 _13167_/X sky130_fd_sc_hd__or2_1
XFILLER_97_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ _22789_/Q _22757_/Q _22658_/Q _22725_/Q _11151_/A _11953_/A vssd1 vssd1 vccd1
+ vccd1 _12118_/X sky130_fd_sc_hd__mux4_2
XFILLER_257_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17975_ _22835_/Q _17972_/X _17959_/A input266/X _17966_/X vssd1 vssd1 vccd1 vccd1
+ _17975_/X sky130_fd_sc_hd__a221o_1
X_13098_ _13107_/A _13097_/X _11235_/A vssd1 vssd1 vccd1 vccd1 _13098_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_306_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater505 _12037_/Y vssd1 vssd1 vccd1 vccd1 _20279_/A sky130_fd_sc_hd__buf_6
XFILLER_78_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19714_ _19714_/A vssd1 vssd1 vccd1 vccd1 _23498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_284_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12049_ _12056_/A _12048_/X _12687_/A vssd1 vssd1 vccd1 vccd1 _12049_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_242_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16926_ input68/X input43/X _17219_/S vssd1 vssd1 vccd1 vccd1 _16926_/X sky130_fd_sc_hd__mux2_8
XFILLER_272_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_348_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19645_ _19188_/X _23468_/Q _19649_/S vssd1 vssd1 vccd1 vccd1 _19646_/A sky130_fd_sc_hd__mux2_1
XFILLER_348_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16857_ _19207_/A vssd1 vssd1 vccd1 vccd1 _16857_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15808_ _23770_/Q _15215_/A _15216_/A _15806_/X _15807_/X vssd1 vssd1 vccd1 vccd1
+ _15808_/X sky130_fd_sc_hd__a221o_2
X_16788_ _22513_/Q _16783_/X _16784_/X input28/X vssd1 vssd1 vccd1 vccd1 _16789_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_65_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19576_ _19576_/A vssd1 vssd1 vccd1 vccd1 _23437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18527_ _18520_/X _18526_/Y _18516_/X vssd1 vssd1 vccd1 vccd1 _23005_/D sky130_fd_sc_hd__a21oi_1
X_15739_ _16186_/A _15723_/Y _15738_/Y _14586_/A vssd1 vssd1 vccd1 vccd1 _15739_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_244_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18458_ _22979_/Q _18465_/B vssd1 vssd1 vccd1 vccd1 _18458_/Y sky130_fd_sc_hd__nand2_1
XFILLER_339_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17409_ _17409_/A vssd1 vssd1 vccd1 vccd1 _22617_/D sky130_fd_sc_hd__clkbuf_1
X_18389_ _15351_/A _18392_/C _18380_/X vssd1 vssd1 vccd1 vccd1 _18389_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_53_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_336_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20420_ _20445_/A vssd1 vssd1 vccd1 vccd1 _20420_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_354_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20351_ _20379_/A _21165_/A vssd1 vssd1 vccd1 vccd1 _20351_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23070_ _23070_/CLK _23070_/D vssd1 vssd1 vccd1 vccd1 _23070_/Q sky130_fd_sc_hd__dfxtp_1
X_20282_ _20192_/X _21766_/A _20280_/Y _20281_/X vssd1 vssd1 vccd1 vccd1 _20660_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_134_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_350_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22021_ _23836_/Q _23770_/Q vssd1 vssd1 vccd1 vccd1 _22023_/A sky130_fd_sc_hd__and2_1
XTAP_6209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_289_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_350_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_331_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_288_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22923_ _22923_/CLK _22923_/D vssd1 vssd1 vccd1 vccd1 _22923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22854_ _22908_/CLK _22854_/D vssd1 vssd1 vccd1 vccd1 _22854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21805_ _15616_/A _21556_/X _21721_/X vssd1 vssd1 vccd1 vccd1 _21809_/A sky130_fd_sc_hd__o21a_1
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22785_ _23367_/CLK _22785_/D vssd1 vssd1 vccd1 vccd1 _22785_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21736_ _21709_/B _21711_/B _21709_/A vssd1 vssd1 vccd1 vccd1 _21740_/A sky130_fd_sc_hd__a21bo_1
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21667_ _21667_/A _21667_/B vssd1 vssd1 vccd1 vccd1 _21669_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11420_ _11424_/A _11420_/B vssd1 vssd1 vccd1 vccd1 _11420_/Y sky130_fd_sc_hd__nor2_1
X_23406_ _23534_/CLK _23406_/D vssd1 vssd1 vccd1 vccd1 _23406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20618_ _14546_/X _20617_/X _20598_/X vssd1 vssd1 vccd1 vccd1 _20618_/X sky130_fd_sc_hd__a21o_1
XFILLER_354_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21598_ _21840_/A vssd1 vssd1 vccd1 vccd1 _21598_/X sky130_fd_sc_hd__buf_2
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_327_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_327_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11351_ _11537_/A vssd1 vssd1 vccd1 vccd1 _11352_/A sky130_fd_sc_hd__buf_2
X_23337_ _23369_/CLK _23337_/D vssd1 vssd1 vccd1 vccd1 _23337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20549_ _20549_/A vssd1 vssd1 vccd1 vccd1 _20724_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_341_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14070_ input239/X _14058_/X _14069_/X vssd1 vssd1 vccd1 vccd1 _14070_/X sky130_fd_sc_hd__a21bo_4
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_298_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23268_ _23578_/CLK _23268_/D vssd1 vssd1 vccd1 vccd1 _23268_/Q sky130_fd_sc_hd__dfxtp_1
X_11282_ _11282_/A vssd1 vssd1 vccd1 vccd1 _11630_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_141_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13021_ _23931_/Q _13020_/Y _13296_/B vssd1 vssd1 vccd1 vccd1 _13022_/B sky130_fd_sc_hd__mux2_1
XFILLER_152_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22219_ _22219_/A _22219_/B vssd1 vssd1 vccd1 vccd1 _22219_/X sky130_fd_sc_hd__or2_1
XFILLER_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23199_ _23582_/CLK _23199_/D vssd1 vssd1 vccd1 vccd1 _23199_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_343_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17760_ _17760_/A vssd1 vssd1 vccd1 vccd1 _22756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14972_ _16079_/A vssd1 vssd1 vccd1 vccd1 _16004_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16711_ _16729_/A vssd1 vssd1 vccd1 vccd1 _16711_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13923_ _13931_/A _13923_/B vssd1 vssd1 vccd1 vccd1 _13923_/Y sky130_fd_sc_hd__nor2_1
XFILLER_267_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17691_ _22726_/Q _17588_/X _17693_/S vssd1 vssd1 vccd1 vccd1 _17692_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16642_ _16664_/A vssd1 vssd1 vccd1 vccd1 _16651_/S sky130_fd_sc_hd__buf_4
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19430_ _19430_/A vssd1 vssd1 vccd1 vccd1 _23372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13854_ _13851_/Y _13852_/Y _13853_/X vssd1 vssd1 vccd1 vccd1 _13855_/B sky130_fd_sc_hd__o21a_2
XFILLER_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_405 _13880_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_416 _14010_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12805_ _12805_/A _15678_/A vssd1 vssd1 vccd1 vccd1 _13532_/D sky130_fd_sc_hd__nor2_4
X_16573_ _15625_/X _22438_/Q _16579_/S vssd1 vssd1 vccd1 vccd1 _16574_/A sky130_fd_sc_hd__mux2_1
XFILLER_308_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_427 _14521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19361_ _23342_/Q _18801_/X _19361_/S vssd1 vssd1 vccd1 vccd1 _19362_/A sky130_fd_sc_hd__mux2_1
X_13785_ _13736_/B _13835_/A _13782_/X _13830_/B vssd1 vssd1 vccd1 vccd1 _13786_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_438 _23912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_449 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15524_ _15523_/X _22275_/Q _15524_/S vssd1 vssd1 vccd1 vccd1 _15525_/A sky130_fd_sc_hd__mux2_1
X_18312_ _18314_/A _18314_/C _18311_/Y vssd1 vssd1 vccd1 vccd1 _22930_/D sky130_fd_sc_hd__o21a_1
XFILLER_71_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12736_ _12993_/A _12735_/X _12721_/X vssd1 vssd1 vccd1 vccd1 _12736_/X sky130_fd_sc_hd__o21a_1
X_19292_ _19197_/X _23311_/Q _19300_/S vssd1 vssd1 vccd1 vccd1 _19293_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18243_ _18243_/A vssd1 vssd1 vccd1 vccd1 _18253_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_187_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15455_ _15455_/A vssd1 vssd1 vccd1 vccd1 _16034_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_349_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ _12801_/A vssd1 vssd1 vccd1 vccd1 _12667_/X sky130_fd_sc_hd__buf_2
XFILLER_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14406_ _14483_/A vssd1 vssd1 vccd1 vccd1 _20161_/A sky130_fd_sc_hd__buf_4
XFILLER_129_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11618_ _23478_/Q _23574_/Q _22538_/Q _22342_/Q _12043_/S _11613_/X vssd1 vssd1 vccd1
+ vccd1 _11619_/B sky130_fd_sc_hd__mux4_1
X_18174_ _18277_/A vssd1 vssd1 vccd1 vccd1 _18423_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15386_ _15386_/A vssd1 vssd1 vccd1 vccd1 _15386_/Y sky130_fd_sc_hd__inv_2
XFILLER_329_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_318_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12598_ _14368_/A _12602_/A vssd1 vssd1 vccd1 vccd1 _12600_/A sky130_fd_sc_hd__nor2_2
XFILLER_128_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17125_ _21720_/A _17123_/X _17234_/S vssd1 vssd1 vccd1 vccd1 _17125_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14337_ _15132_/S vssd1 vssd1 vccd1 vccd1 _15133_/A sky130_fd_sc_hd__buf_2
XFILLER_305_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11549_ _22483_/Q _22643_/Q _22322_/Q _23458_/Q _11543_/X _13276_/A vssd1 vssd1 vccd1
+ vccd1 _11549_/X sky130_fd_sc_hd__mux4_1
XFILLER_345_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17056_ _16951_/X _17055_/X _17078_/A _16996_/X vssd1 vssd1 vccd1 vccd1 _17056_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14268_ _12235_/B _13242_/B _14348_/A vssd1 vssd1 vccd1 vccd1 _14268_/X sky130_fd_sc_hd__mux2_1
XFILLER_333_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16007_ _14987_/B _13570_/B _15574_/X _16006_/X vssd1 vssd1 vccd1 vccd1 _16007_/X
+ sky130_fd_sc_hd__o211a_1
X_13219_ _22801_/Q _22769_/Q _22670_/Q _22737_/Q _11526_/A _11519_/A vssd1 vssd1 vccd1
+ vccd1 _13219_/X sky130_fd_sc_hd__mux4_1
XFILLER_315_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _14199_/A _14199_/B _14199_/C vssd1 vssd1 vccd1 vccd1 _20549_/A sky130_fd_sc_hd__and3_2
XFILLER_298_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_286_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_340_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_10_0_wb_clk_i clkbuf_3_5_1_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_10_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_257_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_300_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _22830_/Q _17950_/X _17957_/X _17948_/X vssd1 vssd1 vccd1 vccd1 _22830_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_300_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_wb_clk_i clkbuf_opt_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23453_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_273_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16909_ _16908_/X _22550_/Q _16909_/S vssd1 vssd1 vccd1 vccd1 _16910_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17889_ _17908_/A _18021_/B vssd1 vssd1 vccd1 vccd1 _17981_/A sky130_fd_sc_hd__nor2_2
XFILLER_272_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23502_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_122_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19628_ _19684_/A vssd1 vssd1 vccd1 vccd1 _19697_/S sky130_fd_sc_hd__buf_6
XFILLER_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19559_ _19559_/A vssd1 vssd1 vccd1 vccd1 _23429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22570_ _23646_/CLK _22570_/D vssd1 vssd1 vccd1 vccd1 _22570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_278_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21521_ _21517_/Y _21519_/X _21840_/A vssd1 vssd1 vccd1 vccd1 _21521_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_355_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21452_ _21452_/A _21452_/B vssd1 vssd1 vccd1 vccd1 _21452_/X sky130_fd_sc_hd__and2_1
XFILLER_348_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20403_ _20226_/X _16194_/X _20401_/X _20402_/Y vssd1 vssd1 vccd1 vccd1 _20765_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_135_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21383_ _14195_/A _21336_/A _21520_/A vssd1 vssd1 vccd1 vccd1 _21600_/A sky130_fd_sc_hd__a21oi_4
XFILLER_308_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_323_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_336_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_351_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23122_ _23474_/CLK _23122_/D vssd1 vssd1 vccd1 vccd1 _23122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20334_ _20334_/A _20400_/B vssd1 vssd1 vccd1 vccd1 _20336_/B sky130_fd_sc_hd__nor2_1
XFILLER_324_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_323_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20265_ _15408_/A _20261_/X _20267_/B vssd1 vssd1 vccd1 vccd1 _20265_/X sky130_fd_sc_hd__o21a_1
X_23053_ _23367_/CLK _23053_/D vssd1 vssd1 vccd1 vccd1 _23053_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_351_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_295_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22004_ _21515_/B _22002_/X _22003_/Y _21767_/X vssd1 vssd1 vccd1 vccd1 _22004_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_6039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20196_ _20220_/A vssd1 vssd1 vccd1 vccd1 _20196_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput105 dout0[8] vssd1 vssd1 vccd1 vccd1 input105/X sky130_fd_sc_hd__buf_2
Xinput116 dout1[18] vssd1 vssd1 vccd1 vccd1 input116/X sky130_fd_sc_hd__clkbuf_1
XTAP_5327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput127 dout1[28] vssd1 vssd1 vccd1 vccd1 input127/X sky130_fd_sc_hd__clkbuf_1
XTAP_5338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput138 dout1[38] vssd1 vssd1 vccd1 vccd1 input138/X sky130_fd_sc_hd__buf_2
XTAP_5349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput149 dout1[48] vssd1 vssd1 vccd1 vccd1 input149/X sky130_fd_sc_hd__buf_2
XFILLER_236_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22906_ _22929_/CLK _22906_/D vssd1 vssd1 vccd1 vccd1 _22906_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23886_ _23910_/CLK _23886_/D vssd1 vssd1 vccd1 vccd1 _23886_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22837_ _23632_/CLK _22837_/D vssd1 vssd1 vccd1 vccd1 _22837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _13570_/A _13570_/B vssd1 vssd1 vccd1 vccd1 _13570_/Y sky130_fd_sc_hd__nand2_1
X_22768_ _23068_/CLK _22768_/D vssd1 vssd1 vccd1 vccd1 _22768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_339_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_319_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _13359_/B vssd1 vssd1 vccd1 vccd1 _13362_/B sky130_fd_sc_hd__buf_4
XFILLER_157_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21719_ _21719_/A _21845_/A vssd1 vssd1 vccd1 vccd1 _21719_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22699_ _23068_/CLK _22699_/D vssd1 vssd1 vccd1 vccd1 _22699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _19191_/A vssd1 vssd1 vccd1 vccd1 _15240_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_346_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12452_ _23398_/Q _23014_/Q _23366_/Q _23334_/Q _11411_/A _12449_/X vssd1 vssd1 vccd1
+ vccd1 _12452_/X sky130_fd_sc_hd__mux4_2
XFILLER_327_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11403_ _11403_/A vssd1 vssd1 vccd1 vccd1 _11403_/X sky130_fd_sc_hd__buf_2
X_15171_ _15171_/A vssd1 vssd1 vccd1 vccd1 _15995_/A sky130_fd_sc_hd__buf_4
XFILLER_126_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12383_ _12383_/A _12383_/B vssd1 vssd1 vccd1 vccd1 _12383_/X sky130_fd_sc_hd__or2_1
XFILLER_327_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14122_ _22845_/Q _14115_/X _14120_/X _18018_/B vssd1 vssd1 vccd1 vccd1 _14122_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_193_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11334_ _12998_/A vssd1 vssd1 vccd1 vccd1 _13006_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_181_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_326_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_341_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18930_ _18930_/A vssd1 vssd1 vccd1 vccd1 _23165_/D sky130_fd_sc_hd__clkbuf_1
X_14053_ input229/X _14038_/X _14052_/X vssd1 vssd1 vccd1 vccd1 _14053_/X sky130_fd_sc_hd__a21bo_4
XTAP_7230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11265_ _11404_/B vssd1 vssd1 vccd1 vccd1 _12371_/B sky130_fd_sc_hd__clkbuf_2
XTAP_7241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13004_ _11515_/A _13003_/X _12707_/A vssd1 vssd1 vccd1 vccd1 _13004_/X sky130_fd_sc_hd__o21a_1
XTAP_7263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18861_ _18861_/A vssd1 vssd1 vccd1 vccd1 _23136_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11196_ _11196_/A vssd1 vssd1 vccd1 vccd1 _21077_/C sky130_fd_sc_hd__buf_6
XTAP_7296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17812_ _17812_/A vssd1 vssd1 vccd1 vccd1 _22779_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18792_ _18792_/A vssd1 vssd1 vccd1 vccd1 _18792_/X sky130_fd_sc_hd__clkbuf_2
XTAP_6595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14955_ _14953_/Y _14954_/X _15088_/S vssd1 vssd1 vccd1 vccd1 _14955_/X sky130_fd_sc_hd__mux2_1
X_17743_ _22749_/Q _17559_/X _17743_/S vssd1 vssd1 vccd1 vccd1 _17744_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_345_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13906_ _13906_/A _13906_/B vssd1 vssd1 vccd1 vccd1 _13906_/Y sky130_fd_sc_hd__xnor2_4
X_17674_ _22718_/Q _17562_/X _17682_/S vssd1 vssd1 vccd1 vccd1 _17675_/A sky130_fd_sc_hd__mux2_1
X_14886_ _14976_/B _14886_/B vssd1 vssd1 vccd1 vccd1 _21384_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_202 _19969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19413_ _19481_/S vssd1 vssd1 vccd1 vccd1 _19422_/S sky130_fd_sc_hd__buf_6
XINSDIODE2_213 _21300_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13837_ _13830_/Y _13835_/Y _13836_/Y _13730_/X vssd1 vssd1 vccd1 vccd1 _14056_/C
+ sky130_fd_sc_hd__a22o_2
XFILLER_35_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16625_ _22461_/Q _16230_/X _16629_/S vssd1 vssd1 vccd1 vccd1 _16626_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_224 _15057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_235 _15995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_246 _15408_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16556_ _16556_/A vssd1 vssd1 vccd1 vccd1 _22430_/D sky130_fd_sc_hd__clkbuf_1
X_19344_ _23334_/Q _18776_/X _19350_/S vssd1 vssd1 vccd1 vccd1 _19345_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_257 _15606_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13768_ _13768_/A _13771_/B vssd1 vssd1 vccd1 vccd1 _13768_/Y sky130_fd_sc_hd__nand2_1
XINSDIODE2_268 _15656_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_279 _21954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_349_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12719_ _23416_/Q _23032_/Q _23384_/Q _23352_/Q _12029_/X _12009_/X vssd1 vssd1 vccd1
+ vccd1 _12720_/B sky130_fd_sc_hd__mux4_1
XFILLER_231_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15507_ _23795_/Q _14917_/A _14919_/A vssd1 vssd1 vccd1 vccd1 _15507_/X sky130_fd_sc_hd__a21o_1
XFILLER_337_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16487_ _15422_/X _22401_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _16488_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19275_ _19275_/A vssd1 vssd1 vccd1 vccd1 _23303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_349_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13699_ _13765_/A _13699_/B _14089_/A vssd1 vssd1 vccd1 vccd1 _13793_/B sky130_fd_sc_hd__nor3_4
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18226_ _22854_/Q _18216_/X _18225_/X _18219_/X vssd1 vssd1 vccd1 vccd1 _22902_/D
+ sky130_fd_sc_hd__o211a_1
X_15438_ _18305_/A _15000_/A _15001_/A _22959_/Q vssd1 vssd1 vccd1 vccd1 _15438_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_337_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18157_ _18157_/A vssd1 vssd1 vccd1 vccd1 _22888_/D sky130_fd_sc_hd__clkbuf_1
X_15369_ _22989_/Q _15416_/A _15417_/A input217/X vssd1 vssd1 vccd1 vccd1 _21676_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_1_wb_clk_i clkbuf_2_0_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_117_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_317_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17108_ _17073_/X _17106_/X _17107_/X _17078_/X vssd1 vssd1 vccd1 vccd1 _17108_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_117_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18088_ _22867_/Q _18081_/X _18087_/X _18075_/X vssd1 vssd1 vccd1 vccd1 _22867_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17039_ _17039_/A vssd1 vssd1 vccd1 vccd1 _17276_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20050_ _23627_/Q vssd1 vssd1 vccd1 vccd1 _20066_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_286_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_344_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23740_ _23915_/CLK _23740_/D vssd1 vssd1 vccd1 vccd1 _23740_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20952_ _23800_/Q _20939_/X _20951_/X _20948_/X vssd1 vssd1 vccd1 vccd1 _23800_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_260_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23671_ _23704_/CLK _23671_/D vssd1 vssd1 vccd1 vccd1 _23671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_281_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20883_ _21215_/A _20883_/B vssd1 vssd1 vccd1 vccd1 _20884_/A sky130_fd_sc_hd__and2_1
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22622_ _23565_/CLK _22622_/D vssd1 vssd1 vccd1 vccd1 _22622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22553_ _23693_/CLK _22553_/D vssd1 vssd1 vccd1 vccd1 _22553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21504_ _21500_/B _21503_/Y _22171_/B vssd1 vssd1 vccd1 vccd1 _21504_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22484_ _23588_/CLK _22484_/D vssd1 vssd1 vccd1 vccd1 _22484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21435_ _21435_/A _21435_/B vssd1 vssd1 vccd1 vccd1 _21435_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_135_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_352_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21366_ _21479_/A vssd1 vssd1 vccd1 vccd1 _21366_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_218_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23105_ _23489_/CLK _23105_/D vssd1 vssd1 vccd1 vccd1 _23105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_352_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20317_ _23671_/Q _20165_/X _20316_/Y _20285_/X vssd1 vssd1 vccd1 vccd1 _23671_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_311_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21297_ _22257_/B _21297_/B _21297_/C _21297_/D vssd1 vssd1 vccd1 vccd1 _21328_/A
+ sky130_fd_sc_hd__nor4_4
XFILLER_289_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23036_ _23354_/CLK _23036_/D vssd1 vssd1 vccd1 vccd1 _23036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_277_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20248_ _21616_/A _20279_/B vssd1 vssd1 vccd1 vccd1 _20250_/B sky130_fd_sc_hd__and2_1
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20179_ _17172_/A _21340_/A _20197_/S vssd1 vssd1 vccd1 vccd1 _20179_/X sky130_fd_sc_hd__mux2_1
XFILLER_276_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_289_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ _23783_/Q _20160_/A _15068_/C vssd1 vssd1 vccd1 vccd1 _14740_/X sky130_fd_sc_hd__or3_1
XFILLER_29_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11952_ _22469_/Q _22629_/Q _12042_/S vssd1 vssd1 vccd1 vccd1 _11952_/X sky130_fd_sc_hd__mux2_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23938_ _23938_/CLK _23938_/D vssd1 vssd1 vccd1 vccd1 _23938_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_291_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _15488_/A _14669_/X _14671_/S vssd1 vssd1 vccd1 vccd1 _14671_/X sky130_fd_sc_hd__mux2_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _23920_/Q vssd1 vssd1 vccd1 vccd1 _21601_/A sky130_fd_sc_hd__inv_8
X_23869_ _23871_/CLK _23869_/D vssd1 vssd1 vccd1 vccd1 _23869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_264_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16410_ _15324_/X _22367_/Q _16418_/S vssd1 vssd1 vccd1 vccd1 _16411_/A sky130_fd_sc_hd__mux2_1
X_13622_ _13342_/A _13625_/B _13497_/A vssd1 vssd1 vccd1 vccd1 _13623_/B sky130_fd_sc_hd__a21oi_2
XFILLER_305_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17390_ _22122_/A vssd1 vssd1 vccd1 vccd1 _17390_/X sky130_fd_sc_hd__buf_4
XFILLER_60_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16341_ _16341_/A vssd1 vssd1 vccd1 vccd1 _22337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13553_ _13555_/A _13555_/B _16128_/S vssd1 vssd1 vccd1 vccd1 _13554_/B sky130_fd_sc_hd__a21o_1
XFILLER_158_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_347_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_349_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19060_ _16873_/X _23223_/Q _19062_/S vssd1 vssd1 vccd1 vccd1 _19061_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12504_ _11659_/A _12503_/X _11818_/A vssd1 vssd1 vccd1 vccd1 _12504_/X sky130_fd_sc_hd__o21a_1
XFILLER_319_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16272_ _16288_/A vssd1 vssd1 vccd1 vccd1 _16285_/S sky130_fd_sc_hd__buf_2
XFILLER_160_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13484_ _13593_/A _20530_/B vssd1 vssd1 vccd1 vccd1 _19969_/D sky130_fd_sc_hd__and2_4
XFILLER_146_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_328_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18011_ _18118_/A _14115_/X _14125_/Y _22845_/Q vssd1 vssd1 vccd1 vccd1 _18011_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15223_ _23821_/Q _15211_/X _15214_/X _15221_/X _15222_/X vssd1 vssd1 vccd1 vccd1
+ _15223_/X sky130_fd_sc_hd__a221o_2
XFILLER_334_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12435_ _12570_/A _12435_/B vssd1 vssd1 vccd1 vccd1 _12435_/Y sky130_fd_sc_hd__nor2_1
XFILLER_355_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15154_ _18286_/A _14509_/X _14513_/X _22953_/Q vssd1 vssd1 vccd1 vccd1 _15154_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_343_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12366_ _12359_/Y _12361_/Y _12363_/Y _12365_/Y _11242_/A vssd1 vssd1 vccd1 vccd1
+ _12366_/X sky130_fd_sc_hd__o221a_1
Xoutput409 _22563_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[10] sky130_fd_sc_hd__buf_2
XFILLER_181_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14105_ _22892_/Q vssd1 vssd1 vccd1 vccd1 _18188_/B sky130_fd_sc_hd__inv_2
XFILLER_271_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11317_ _11317_/A vssd1 vssd1 vccd1 vccd1 _11457_/B sky130_fd_sc_hd__buf_8
XFILLER_314_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_302_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19962_ _19962_/A vssd1 vssd1 vccd1 vccd1 _19962_/X sky130_fd_sc_hd__clkbuf_4
X_15085_ _14782_/X _14776_/X _15085_/S vssd1 vssd1 vccd1 vccd1 _15085_/X sky130_fd_sc_hd__mux2_1
XFILLER_342_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_330_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12297_ _12350_/A _12296_/X _12365_/A vssd1 vssd1 vccd1 vccd1 _12297_/X sky130_fd_sc_hd__a21o_1
XFILLER_99_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18913_ _18913_/A vssd1 vssd1 vccd1 vccd1 _23157_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_351_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14036_ _13770_/B _14036_/B vssd1 vssd1 vccd1 vccd1 _14036_/X sky130_fd_sc_hd__and2b_1
XTAP_7060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11248_ _11222_/Y _11225_/Y _11237_/Y _11239_/Y _11247_/X vssd1 vssd1 vccd1 vccd1
+ _11249_/C sky130_fd_sc_hd__o221a_1
XTAP_7071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19893_ _19893_/A vssd1 vssd1 vccd1 vccd1 _23578_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18844_ _23131_/Q _18843_/X _18850_/S vssd1 vssd1 vccd1 vccd1 _18845_/A sky130_fd_sc_hd__mux2_1
XTAP_6370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11179_ _12130_/A vssd1 vssd1 vccd1 vccd1 _12983_/A sky130_fd_sc_hd__buf_2
XTAP_6381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_314_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18775_ _18775_/A vssd1 vssd1 vccd1 vccd1 _23109_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15987_ _23807_/Q _14917_/X _15067_/X vssd1 vssd1 vccd1 vccd1 _15987_/X sky130_fd_sc_hd__a21o_1
XTAP_5691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17726_ _22742_/Q _17639_/X _17726_/S vssd1 vssd1 vccd1 vccd1 _17727_/A sky130_fd_sc_hd__mux2_1
XFILLER_282_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14938_ _14898_/X _14900_/X _14929_/X _14935_/X _14937_/X vssd1 vssd1 vccd1 vccd1
+ _14939_/B sky130_fd_sc_hd__o32a_4
XFILLER_250_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17657_ _22254_/A vssd1 vssd1 vccd1 vccd1 _17657_/X sky130_fd_sc_hd__buf_6
X_14869_ _23592_/Q _14450_/X _14455_/X _23624_/Q vssd1 vssd1 vccd1 vccd1 _14869_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_330_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16608_ _16664_/A vssd1 vssd1 vccd1 vccd1 _16677_/S sky130_fd_sc_hd__buf_6
XFILLER_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17588_ _18814_/A vssd1 vssd1 vccd1 vccd1 _17588_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19327_ _19249_/X _23327_/Q _19333_/S vssd1 vssd1 vccd1 vccd1 _19328_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_177_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16539_ _16539_/A vssd1 vssd1 vccd1 vccd1 _22422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_338_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19258_ _19258_/A vssd1 vssd1 vccd1 vccd1 _19258_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_338_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18209_ hold2/X _18202_/X _18208_/X _18206_/X vssd1 vssd1 vccd1 vccd1 _22895_/D sky130_fd_sc_hd__o211a_1
XFILLER_337_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19189_ _19188_/X _23276_/Q _19195_/S vssd1 vssd1 vccd1 vccd1 _19190_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_305_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21220_ _21220_/A vssd1 vssd1 vccd1 vccd1 _21258_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21151_ _21083_/X _20525_/D _21150_/X vssd1 vssd1 vccd1 vccd1 _21151_/X sky130_fd_sc_hd__a21o_1
XFILLER_333_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20102_ _23641_/Q _20106_/A _20101_/X vssd1 vssd1 vccd1 vccd1 _20102_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21082_ _23845_/Q vssd1 vssd1 vccd1 vccd1 _21083_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_132_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20033_ _23622_/Q _23621_/Q vssd1 vssd1 vccd1 vccd1 _20042_/D sky130_fd_sc_hd__and2_1
XFILLER_113_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21984_ _21984_/A vssd1 vssd1 vccd1 vccd1 _21984_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23723_ _23755_/CLK _23723_/D vssd1 vssd1 vccd1 vccd1 _23723_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20935_ _23794_/Q _20925_/X _20933_/X _20934_/X vssd1 vssd1 vccd1 vccd1 _23794_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_242_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23654_ _23700_/CLK _23654_/D vssd1 vssd1 vccd1 vccd1 _23654_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20866_ _20727_/B _20864_/X _20865_/X _23773_/Q vssd1 vssd1 vccd1 vccd1 _20867_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22605_ _23646_/CLK _22605_/D vssd1 vssd1 vccd1 vccd1 _22605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_330_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23585_ _23585_/CLK _23585_/D vssd1 vssd1 vccd1 vccd1 _23585_/Q sky130_fd_sc_hd__dfxtp_1
X_20797_ _20806_/A _20797_/B vssd1 vssd1 vccd1 vccd1 _20798_/A sky130_fd_sc_hd__and2_1
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22536_ _23574_/CLK _22536_/D vssd1 vssd1 vccd1 vccd1 _22536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_317_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22467_ _23567_/CLK _22467_/D vssd1 vssd1 vccd1 vccd1 _22467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12220_ _22364_/Q _22396_/Q _22685_/Q _23052_/Q _11920_/A _11815_/A vssd1 vssd1 vccd1
+ vccd1 _12221_/B sky130_fd_sc_hd__mux4_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21418_ _21418_/A _21418_/B vssd1 vssd1 vccd1 vccd1 _21418_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22398_ _23566_/CLK _22398_/D vssd1 vssd1 vccd1 vccd1 _22398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_335_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12151_ _22789_/Q _22757_/Q _22658_/Q _22725_/Q _11457_/C _12009_/A vssd1 vssd1 vccd1
+ vccd1 _12152_/B sky130_fd_sc_hd__mux4_1
XFILLER_340_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21349_ _21319_/A _21348_/Y _21318_/A vssd1 vssd1 vccd1 vccd1 _21353_/A sky130_fd_sc_hd__o21ai_1
XFILLER_108_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_311_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11102_ _11102_/A vssd1 vssd1 vccd1 vccd1 _11102_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_312_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12082_ _12082_/A _12082_/B vssd1 vssd1 vccd1 vccd1 _12082_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23019_ _23531_/CLK _23019_/D vssd1 vssd1 vccd1 vccd1 _23019_/Q sky130_fd_sc_hd__dfxtp_1
X_15910_ _23709_/Q _14905_/A _15909_/X vssd1 vssd1 vccd1 vccd1 _15910_/X sky130_fd_sc_hd__o21a_4
XFILLER_231_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16890_ _16889_/X _22544_/Q _16893_/S vssd1 vssd1 vccd1 vccd1 _16891_/A sky130_fd_sc_hd__mux2_1
XFILLER_277_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_311_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _23835_/Q _14907_/X _15837_/X _15840_/X _14923_/X vssd1 vssd1 vccd1 vccd1
+ _15841_/X sky130_fd_sc_hd__a221o_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_138_wb_clk_i clkbuf_opt_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23692_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18560_ _16822_/X _23015_/Q _18564_/S vssd1 vssd1 vccd1 vccd1 _18561_/A sky130_fd_sc_hd__mux2_1
X_12984_ _23227_/Q _23195_/Q _23163_/Q _23131_/Q _12820_/S _12749_/A vssd1 vssd1 vccd1
+ vccd1 _12985_/B sky130_fd_sc_hd__mux4_2
XFILLER_224_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15772_ _16034_/A _15338_/B _15771_/X vssd1 vssd1 vccd1 vccd1 _15772_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17511_ _17511_/A vssd1 vssd1 vccd1 vccd1 _22662_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14723_ _22513_/Q _14232_/A _14223_/X _14722_/X vssd1 vssd1 vccd1 vccd1 _14724_/B
+ sky130_fd_sc_hd__o22a_1
X_11935_ _23919_/Q _11935_/B vssd1 vssd1 vccd1 vccd1 _11935_/X sky130_fd_sc_hd__or2_4
X_18491_ _18480_/X _18488_/Y _18490_/X vssd1 vssd1 vccd1 vccd1 _22991_/D sky130_fd_sc_hd__a21oi_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17442_ _17442_/A vssd1 vssd1 vccd1 vccd1 _22632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14654_ _14321_/X _14326_/X _14660_/S vssd1 vssd1 vccd1 vccd1 _14654_/X sky130_fd_sc_hd__mux2_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _23406_/Q _23022_/Q _23374_/Q _23342_/Q _11821_/X _11317_/A vssd1 vssd1 vccd1
+ vccd1 _11866_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13605_ _13605_/A _13605_/B vssd1 vssd1 vccd1 vccd1 _13605_/Y sky130_fd_sc_hd__xnor2_4
X_17373_ _17373_/A vssd1 vssd1 vccd1 vccd1 _22606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14585_ _14936_/A _16186_/A vssd1 vssd1 vccd1 vccd1 _14586_/A sky130_fd_sc_hd__nor2_2
X_11797_ _12378_/A vssd1 vssd1 vccd1 vccd1 _11926_/A sky130_fd_sc_hd__buf_4
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_319_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_300_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19112_ _19112_/A vssd1 vssd1 vccd1 vccd1 _23245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16324_ _16381_/S vssd1 vssd1 vccd1 vccd1 _16333_/S sky130_fd_sc_hd__buf_6
X_13536_ _13536_/A _13536_/B vssd1 vssd1 vccd1 vccd1 _13536_/Y sky130_fd_sc_hd__nand2_1
XFILLER_201_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16255_ _18820_/A vssd1 vssd1 vccd1 vccd1 _16255_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19043_ _16847_/X _23215_/Q _19051_/S vssd1 vssd1 vccd1 vccd1 _19044_/A sky130_fd_sc_hd__mux2_1
XFILLER_319_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13467_ _13467_/A vssd1 vssd1 vccd1 vccd1 _13593_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_174_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_334_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15206_ _22922_/Q _15299_/B vssd1 vssd1 vccd1 vccd1 _15206_/X sky130_fd_sc_hd__and2_1
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12418_ _22359_/Q _22391_/Q _22680_/Q _23047_/Q _12424_/S _12538_/A vssd1 vssd1 vccd1
+ vccd1 _12419_/B sky130_fd_sc_hd__mux4_2
XFILLER_127_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16186_ _16186_/A _16186_/B _16186_/C vssd1 vssd1 vccd1 vccd1 _16186_/X sky130_fd_sc_hd__and3_1
X_13398_ _13579_/A vssd1 vssd1 vccd1 vccd1 _13399_/B sky130_fd_sc_hd__inv_2
XFILLER_182_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15137_ _15131_/Y _15136_/Y _15491_/S vssd1 vssd1 vccd1 vccd1 _15137_/X sky130_fd_sc_hd__mux2_1
XFILLER_343_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12349_ _22296_/Q _23432_/Q _12349_/S vssd1 vssd1 vccd1 vccd1 _12350_/B sky130_fd_sc_hd__mux2_1
XFILLER_331_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19945_ _19975_/D _19971_/B _19944_/Y vssd1 vssd1 vccd1 vccd1 _23597_/D sky130_fd_sc_hd__o21a_1
X_15068_ _23787_/Q _20160_/A _15068_/C vssd1 vssd1 vccd1 vccd1 _15068_/X sky130_fd_sc_hd__or3_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_302_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14019_ _14072_/B _14036_/B _14019_/C vssd1 vssd1 vccd1 vccd1 _14019_/X sky130_fd_sc_hd__and3_1
XFILLER_141_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_325_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19876_ _16252_/X _23571_/Q _19876_/S vssd1 vssd1 vccd1 vccd1 _19877_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_296_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18827_ _18827_/A vssd1 vssd1 vccd1 vccd1 _18827_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_255_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18758_ _18758_/A vssd1 vssd1 vccd1 vccd1 _23103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_255_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_341_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17709_ _22734_/Q _17614_/X _17715_/S vssd1 vssd1 vccd1 vccd1 _17710_/A sky130_fd_sc_hd__mux2_1
XFILLER_247_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18689_ _23073_/Q _17636_/X _18691_/S vssd1 vssd1 vccd1 vccd1 _18690_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20720_ _12841_/Y _20701_/X _20719_/Y vssd1 vssd1 vccd1 vccd1 _20721_/C sky130_fd_sc_hd__a21oi_2
XFILLER_251_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20651_ _12137_/Y _20648_/X _20650_/Y vssd1 vssd1 vccd1 vccd1 _20652_/C sky130_fd_sc_hd__a21oi_1
XFILLER_210_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23370_ _23370_/CLK _23370_/D vssd1 vssd1 vccd1 vccd1 _23370_/Q sky130_fd_sc_hd__dfxtp_1
X_20582_ _17020_/A _20572_/X _20581_/Y vssd1 vssd1 vccd1 vccd1 _20583_/C sky130_fd_sc_hd__a21oi_2
XFILLER_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22321_ _23880_/CLK _22321_/D vssd1 vssd1 vccd1 vccd1 _22321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_326_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_307_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22252_ _23943_/Q _22253_/S _22251_/Y vssd1 vssd1 vccd1 vccd1 _23943_/D sky130_fd_sc_hd__o21a_1
XFILLER_293_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21203_ _21243_/A vssd1 vssd1 vccd1 vccd1 _21227_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_322_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22183_ _22183_/A _22183_/B vssd1 vssd1 vccd1 vccd1 _22183_/X sky130_fd_sc_hd__xor2_4
XFILLER_105_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_333_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_333_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21134_ _21134_/A _21134_/B vssd1 vssd1 vccd1 vccd1 _23861_/D sky130_fd_sc_hd__nor2_1
XFILLER_305_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21065_ _22151_/A _20996_/B _21064_/Y _21061_/X vssd1 vssd1 vccd1 vccd1 _23840_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20016_ _23616_/Q _20016_/B _20016_/C vssd1 vssd1 vccd1 vccd1 _20026_/C sky130_fd_sc_hd__and3_1
XFILLER_47_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21967_ _22234_/A _21967_/B vssd1 vssd1 vccd1 vccd1 _21967_/Y sky130_fd_sc_hd__nor2_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _23408_/Q _23024_/Q _23376_/Q _23344_/Q _11777_/S _11590_/A vssd1 vssd1 vccd1
+ vccd1 _11720_/X sky130_fd_sc_hd__mux4_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23706_ _23706_/CLK _23706_/D vssd1 vssd1 vccd1 vccd1 _23706_/Q sky130_fd_sc_hd__dfxtp_4
X_20918_ _23788_/Q _20911_/X _20917_/X _20906_/X vssd1 vssd1 vccd1 vccd1 _23788_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21898_ _21898_/A _22048_/A vssd1 vssd1 vccd1 vccd1 _21898_/Y sky130_fd_sc_hd__nand2_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23637_ _23637_/CLK _23637_/D vssd1 vssd1 vccd1 vccd1 _23637_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_214_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11651_ _11651_/A vssd1 vssd1 vccd1 vccd1 _11652_/A sky130_fd_sc_hd__buf_6
X_20849_ _20861_/A _20849_/B vssd1 vssd1 vccd1 vccd1 _20850_/A sky130_fd_sc_hd__and2_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14370_ _21335_/A _14524_/B _14370_/C vssd1 vssd1 vccd1 vccd1 _14370_/X sky130_fd_sc_hd__and3_1
X_23568_ _23568_/CLK _23568_/D vssd1 vssd1 vccd1 vccd1 _23568_/Q sky130_fd_sc_hd__dfxtp_1
X_11582_ _11582_/A vssd1 vssd1 vccd1 vccd1 _11957_/A sky130_fd_sc_hd__buf_6
XFILLER_11_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_302_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13321_ _13548_/A _13321_/B vssd1 vssd1 vccd1 vccd1 _13410_/C sky130_fd_sc_hd__xnor2_2
XFILLER_357_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22519_ _22520_/CLK _22519_/D vssd1 vssd1 vccd1 vccd1 _22519_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_344_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23499_ _23563_/CLK _23499_/D vssd1 vssd1 vccd1 vccd1 _23499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_346_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16040_ _17267_/A _16039_/C _23938_/Q vssd1 vssd1 vccd1 vccd1 _16041_/B sky130_fd_sc_hd__a21oi_1
X_13252_ _22805_/Q _22773_/Q _22674_/Q _22741_/Q _11492_/S _11200_/A vssd1 vssd1 vccd1
+ vccd1 _13253_/B sky130_fd_sc_hd__mux4_1
XFILLER_10_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_344_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12203_ _12260_/A _12203_/B _12203_/C vssd1 vssd1 vccd1 vccd1 _13727_/A sky130_fd_sc_hd__or3_4
XFILLER_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13183_ _13176_/X _13178_/X _13180_/X _13182_/X _11277_/A vssd1 vssd1 vccd1 vccd1
+ _13184_/C sky130_fd_sc_hd__a221o_1
XFILLER_89_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12134_ _12134_/A _12134_/B _12134_/C vssd1 vssd1 vccd1 vccd1 _13858_/A sky130_fd_sc_hd__nor3_4
XFILLER_151_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17991_ _17991_/A vssd1 vssd1 vccd1 vccd1 _18005_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_297_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19730_ _19207_/X _23506_/Q _19732_/S vssd1 vssd1 vccd1 vccd1 _19731_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16942_ _16942_/A _21320_/A _16942_/C vssd1 vssd1 vccd1 vccd1 _17145_/A sky130_fd_sc_hd__nor3_2
X_12065_ _12065_/A _15492_/S vssd1 vssd1 vccd1 vccd1 _13351_/A sky130_fd_sc_hd__nor2_2
XFILLER_296_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19661_ _19661_/A vssd1 vssd1 vccd1 vccd1 _23475_/D sky130_fd_sc_hd__clkbuf_1
X_16873_ _19223_/A vssd1 vssd1 vccd1 vccd1 _16873_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_293_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_292_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18612_ _18612_/A vssd1 vssd1 vccd1 vccd1 _23038_/D sky130_fd_sc_hd__clkbuf_1
X_15824_ _15823_/X _22282_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15825_/A sky130_fd_sc_hd__mux2_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19592_ _19592_/A vssd1 vssd1 vccd1 vccd1 _23444_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18543_ _18537_/B _18550_/C _18542_/Y _18203_/C vssd1 vssd1 vccd1 vccd1 _18544_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ _22283_/Q _23099_/Q _23515_/Q _22444_/Q _12921_/S _12749_/X vssd1 vssd1 vccd1
+ vccd1 _12968_/B sky130_fd_sc_hd__mux4_1
X_15755_ _22934_/Q _16168_/B vssd1 vssd1 vccd1 vccd1 _15755_/X sky130_fd_sc_hd__and2_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ _19169_/A vssd1 vssd1 vccd1 vccd1 _14706_/X sky130_fd_sc_hd__buf_2
X_11918_ _12321_/A vssd1 vssd1 vccd1 vccd1 _12397_/A sky130_fd_sc_hd__clkbuf_4
X_18474_ _18467_/X _18473_/Y _18463_/X vssd1 vssd1 vccd1 vccd1 _22985_/D sky130_fd_sc_hd__a21oi_1
XFILLER_261_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15686_ _23607_/Q _14732_/X _14734_/X _23639_/Q vssd1 vssd1 vccd1 vccd1 _15686_/X
+ sky130_fd_sc_hd__o22a_2
X_12898_ _22798_/Q _22766_/Q _22667_/Q _22734_/Q _12792_/X _12793_/X vssd1 vssd1 vccd1
+ vccd1 _12898_/X sky130_fd_sc_hd__mux4_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _17425_/A vssd1 vssd1 vccd1 vccd1 _22624_/D sky130_fd_sc_hd__clkbuf_1
X_14637_ _14305_/X _14308_/Y _14651_/A vssd1 vssd1 vccd1 vccd1 _14637_/X sky130_fd_sc_hd__mux2_1
X_11849_ _11853_/A _11849_/B vssd1 vssd1 vccd1 vccd1 _11849_/Y sky130_fd_sc_hd__nor2_1
XFILLER_221_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17356_ _22599_/Q input193/X _17358_/S vssd1 vssd1 vccd1 vccd1 _17357_/A sky130_fd_sc_hd__mux2_1
X_14568_ _14568_/A vssd1 vssd1 vccd1 vccd1 _15367_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_220_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_35_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23068_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_348_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_335_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16307_ _22324_/Q _16306_/X _16307_/S vssd1 vssd1 vccd1 vccd1 _16308_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_307_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13519_ _13942_/A _15198_/A vssd1 vssd1 vccd1 vccd1 _13935_/A sky130_fd_sc_hd__or2_2
X_14499_ _14755_/A _14456_/X _14494_/X _14498_/X vssd1 vssd1 vccd1 vccd1 _14499_/X
+ sky130_fd_sc_hd__o22a_1
X_17287_ input99/X input63/X _17314_/S vssd1 vssd1 vccd1 vccd1 _17287_/X sky130_fd_sc_hd__mux2_8
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19026_ _19026_/A vssd1 vssd1 vccd1 vccd1 _23207_/D sky130_fd_sc_hd__clkbuf_1
X_16238_ _16238_/A vssd1 vssd1 vccd1 vccd1 _22302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_350_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16169_ _23620_/Q _15589_/A _15590_/A _23652_/Q vssd1 vssd1 vccd1 vccd1 _16169_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_6_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_331_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_330_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_303_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19928_ _23593_/Q _19926_/A _18012_/X vssd1 vssd1 vccd1 vccd1 _19929_/B sky130_fd_sc_hd__o21ai_1
XFILLER_287_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19859_ _16227_/X _23563_/Q _19865_/S vssd1 vssd1 vccd1 vccd1 _19860_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22870_ _23632_/CLK _22870_/D vssd1 vssd1 vccd1 vccd1 _22870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21821_ _21821_/A _21821_/B vssd1 vssd1 vccd1 vccd1 _21822_/B sky130_fd_sc_hd__xnor2_1
XFILLER_243_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21752_ _21801_/C _21752_/B vssd1 vssd1 vccd1 vccd1 _21752_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_212_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20703_ _13454_/A _20692_/X _20702_/X vssd1 vssd1 vccd1 vccd1 _20703_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_357_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21683_ _21683_/A vssd1 vssd1 vccd1 vccd1 _21683_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23422_ _23422_/CLK _23422_/D vssd1 vssd1 vccd1 vccd1 _23422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_357_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20634_ _13951_/B _20632_/X _20633_/X vssd1 vssd1 vccd1 vccd1 _20635_/C sky130_fd_sc_hd__o21a_1
XFILLER_221_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23353_ _23545_/CLK _23353_/D vssd1 vssd1 vccd1 vccd1 _23353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_339_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20565_ _20662_/A vssd1 vssd1 vccd1 vccd1 _20732_/A sky130_fd_sc_hd__buf_2
XFILLER_138_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22304_ _23568_/CLK _22304_/D vssd1 vssd1 vccd1 vccd1 _22304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_354_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23284_ _23414_/CLK _23284_/D vssd1 vssd1 vccd1 vccd1 _23284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20496_ _21333_/A _21333_/B vssd1 vssd1 vccd1 vccd1 _20500_/A sky130_fd_sc_hd__xor2_2
XFILLER_106_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22235_ _22218_/A _22223_/A _17315_/X vssd1 vssd1 vccd1 vccd1 _22235_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_316_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22166_ _22166_/A _22171_/A vssd1 vssd1 vccd1 vccd1 _22166_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21117_ _21121_/A _21117_/B vssd1 vssd1 vccd1 vccd1 _23854_/D sky130_fd_sc_hd__nor2_1
XFILLER_132_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22097_ _17267_/A _21867_/X _22096_/X _21865_/X vssd1 vssd1 vccd1 vccd1 _22100_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21048_ _23834_/Q _21048_/B vssd1 vssd1 vccd1 vccd1 _21048_/X sky130_fd_sc_hd__or2_1
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13870_ _11452_/B _13836_/B _13721_/B vssd1 vssd1 vccd1 vccd1 _13871_/B sky130_fd_sc_hd__a21oi_1
XFILLER_86_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12821_ _11587_/A _12820_/X _12683_/A vssd1 vssd1 vccd1 vccd1 _12821_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22999_ _23592_/CLK _22999_/D vssd1 vssd1 vccd1 vccd1 _22999_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12752_ _11587_/A _12751_/X _12130_/A vssd1 vssd1 vccd1 vccd1 _12752_/X sky130_fd_sc_hd__a21o_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15540_ _15011_/A _14380_/Y _15538_/Y _15539_/Y vssd1 vssd1 vccd1 vccd1 _15540_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_199_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_349_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11703_ _11703_/A vssd1 vssd1 vccd1 vccd1 _11839_/A sky130_fd_sc_hd__buf_6
X_15471_ _22991_/Q _15620_/A _15621_/A input219/X vssd1 vssd1 vccd1 vccd1 _21741_/A
+ sky130_fd_sc_hd__a22o_4
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12683_ _12683_/A vssd1 vssd1 vccd1 vccd1 _12836_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_231_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _22900_/Q _14394_/A _14164_/A _22593_/Q vssd1 vssd1 vccd1 vccd1 _16942_/A
+ sky130_fd_sc_hd__a22o_2
X_17210_ input91/X input56/X _17266_/S vssd1 vssd1 vccd1 vccd1 _17210_/X sky130_fd_sc_hd__mux2_8
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11634_ _12383_/A vssd1 vssd1 vccd1 vccd1 _12401_/A sky130_fd_sc_hd__buf_4
X_18190_ _18162_/A _18167_/X _18118_/A vssd1 vssd1 vccd1 vccd1 _18191_/D sky130_fd_sc_hd__o21ai_1
XFILLER_230_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17141_ _17255_/A vssd1 vssd1 vccd1 vccd1 _17141_/X sky130_fd_sc_hd__buf_2
X_14353_ _14665_/S vssd1 vssd1 vccd1 vccd1 _14840_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_344_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11565_ _11565_/A vssd1 vssd1 vccd1 vccd1 _11566_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_11_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_357_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13304_ _13318_/A _13319_/A _13319_/B _11555_/A _11557_/A vssd1 vssd1 vccd1 vccd1
+ _13316_/B sky130_fd_sc_hd__o32a_1
X_17072_ _22810_/Q _17244_/B _17244_/C vssd1 vssd1 vccd1 vccd1 _17073_/A sky130_fd_sc_hd__and3_1
XFILLER_196_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14284_ _14331_/S vssd1 vssd1 vccd1 vccd1 _14646_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_7_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11496_ _23234_/Q _23202_/Q _23170_/Q _23138_/Q _11432_/X _11435_/X vssd1 vssd1 vccd1
+ vccd1 _11497_/B sky130_fd_sc_hd__mux4_1
XFILLER_344_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13235_ _13242_/A _13241_/A vssd1 vssd1 vccd1 vccd1 _13237_/A sky130_fd_sc_hd__and2_1
X_16023_ _23808_/Q _15219_/X _14606_/X vssd1 vssd1 vccd1 vccd1 _16023_/X sky130_fd_sc_hd__a21o_1
XFILLER_171_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13166_ _22286_/Q _23102_/Q _23518_/Q _22447_/Q _11532_/X _11544_/A vssd1 vssd1 vccd1
+ vccd1 _13167_/B sky130_fd_sc_hd__mux4_2
XFILLER_313_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_298_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12117_ _12117_/A _12117_/B vssd1 vssd1 vccd1 vccd1 _12117_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_153_wb_clk_i _23945_/CLK vssd1 vssd1 vccd1 vccd1 _23911_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_112_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17974_ _22835_/Q _17965_/X _17973_/X _17963_/X vssd1 vssd1 vccd1 vccd1 _22835_/D
+ sky130_fd_sc_hd__o211a_1
X_13097_ _22383_/Q _22415_/Q _22704_/Q _23071_/Q _13034_/S _13096_/X vssd1 vssd1 vccd1
+ vccd1 _13097_/X sky130_fd_sc_hd__mux4_2
XFILLER_151_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19713_ _19181_/X _23498_/Q _19721_/S vssd1 vssd1 vccd1 vccd1 _19714_/A sky130_fd_sc_hd__mux2_1
X_12048_ _22371_/Q _22403_/Q _22692_/Q _23059_/Q _11972_/X _11973_/X vssd1 vssd1 vccd1
+ vccd1 _12048_/X sky130_fd_sc_hd__mux4_1
X_16925_ _22809_/Q _17241_/B vssd1 vssd1 vccd1 vccd1 _17000_/A sky130_fd_sc_hd__nand2_1
XFILLER_78_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19644_ _19644_/A vssd1 vssd1 vccd1 vccd1 _23467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_293_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16856_ _16856_/A vssd1 vssd1 vccd1 vccd1 _22533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_281_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_348_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15807_ _23802_/Q _15219_/A _14919_/A vssd1 vssd1 vccd1 vccd1 _15807_/X sky130_fd_sc_hd__a21o_1
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19575_ _23437_/Q _19191_/A _19577_/S vssd1 vssd1 vccd1 vccd1 _19576_/A sky130_fd_sc_hd__mux2_1
XFILLER_281_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16787_ _16787_/A vssd1 vssd1 vccd1 vccd1 _22512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13999_ _14000_/A _14097_/A vssd1 vssd1 vccd1 vccd1 _13999_/Y sky130_fd_sc_hd__nor2_4
XFILLER_225_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18526_ _23005_/Q _18530_/B vssd1 vssd1 vccd1 vccd1 _18526_/Y sky130_fd_sc_hd__nand2_1
X_15738_ _15738_/A vssd1 vssd1 vccd1 vccd1 _15738_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_80_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18457_ _18451_/X _18455_/Y _22260_/A vssd1 vssd1 vccd1 vccd1 _22978_/D sky130_fd_sc_hd__a21oi_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15669_ _15668_/X _22278_/Q _15750_/S vssd1 vssd1 vccd1 vccd1 _15670_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17408_ _22617_/Q _16217_/X _17410_/S vssd1 vssd1 vccd1 vccd1 _17409_/A sky130_fd_sc_hd__mux2_1
X_18388_ _22956_/Q _18386_/B _18387_/Y vssd1 vssd1 vccd1 vccd1 _22956_/D sky130_fd_sc_hd__o21a_1
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_336_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17339_ _22591_/Q input208/X _17347_/S vssd1 vssd1 vccd1 vccd1 _17340_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_336_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20350_ _20226_/X _22032_/A _20349_/X vssd1 vssd1 vccd1 vccd1 _21165_/A sky130_fd_sc_hd__a21oi_4
XFILLER_128_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19009_ _19009_/A vssd1 vssd1 vccd1 vccd1 _23200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20281_ _20275_/A _20279_/Y _20220_/A vssd1 vssd1 vccd1 vccd1 _20281_/X sky130_fd_sc_hd__o21a_1
XFILLER_143_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_288_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22020_ _21993_/B _21995_/B _21993_/A vssd1 vssd1 vccd1 vccd1 _22024_/A sky130_fd_sc_hd__o21bai_1
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_350_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_289_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22922_ _22923_/CLK _22922_/D vssd1 vssd1 vccd1 vccd1 _22922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22853_ _22908_/CLK _22853_/D vssd1 vssd1 vccd1 vccd1 _22853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21804_ _21800_/X _21804_/B _21804_/C vssd1 vssd1 vccd1 vccd1 _21812_/B sky130_fd_sc_hd__and3b_2
X_22784_ _23144_/CLK _22784_/D vssd1 vssd1 vccd1 vccd1 _22784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21735_ _23826_/Q _21734_/Y _22083_/A vssd1 vssd1 vccd1 vccd1 _21735_/X sky130_fd_sc_hd__mux2_1
XFILLER_358_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21666_ _23824_/Q _23758_/Q vssd1 vssd1 vccd1 vccd1 _21667_/B sky130_fd_sc_hd__nand2_1
XFILLER_200_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23405_ _23565_/CLK _23405_/D vssd1 vssd1 vccd1 vccd1 _23405_/Q sky130_fd_sc_hd__dfxtp_1
X_20617_ _20724_/A vssd1 vssd1 vccd1 vccd1 _20617_/X sky130_fd_sc_hd__clkbuf_2
X_21597_ _14195_/X _21518_/X _21517_/B _15277_/B vssd1 vssd1 vccd1 vccd1 _21597_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_338_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ _12721_/A vssd1 vssd1 vccd1 vccd1 _11537_/A sky130_fd_sc_hd__clkbuf_4
X_23336_ _23368_/CLK _23336_/D vssd1 vssd1 vccd1 vccd1 _23336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20548_ _14970_/S _13481_/B _13455_/Y vssd1 vssd1 vccd1 vccd1 _20632_/A sky130_fd_sc_hd__a21oi_4
XFILLER_327_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_353_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_327_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_342_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23267_ _23555_/CLK _23267_/D vssd1 vssd1 vccd1 vccd1 _23267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11281_ _11818_/A vssd1 vssd1 vccd1 vccd1 _11282_/A sky130_fd_sc_hd__buf_2
XFILLER_353_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20479_ _20731_/A _20467_/X _20478_/X _20472_/X vssd1 vssd1 vccd1 vccd1 _23710_/D
+ sky130_fd_sc_hd__o211a_1
X_13020_ _20327_/A vssd1 vssd1 vccd1 vccd1 _13020_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22218_ _22218_/A _22218_/B vssd1 vssd1 vccd1 vccd1 _22222_/A sky130_fd_sc_hd__or2_1
XFILLER_152_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23198_ _23550_/CLK _23198_/D vssd1 vssd1 vccd1 vccd1 _23198_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_350_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22149_ _23841_/Q _23775_/Q vssd1 vssd1 vccd1 vccd1 _22150_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14971_ _14882_/A _14939_/X _14959_/Y _14822_/X _14970_/X vssd1 vssd1 vccd1 vccd1
+ _14971_/X sky130_fd_sc_hd__a32o_2
XTAP_6799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16710_ _16710_/A vssd1 vssd1 vccd1 vccd1 _22491_/D sky130_fd_sc_hd__clkbuf_1
X_13922_ _21500_/A vssd1 vssd1 vccd1 vccd1 _13923_/B sky130_fd_sc_hd__buf_6
XFILLER_248_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17690_ _17690_/A vssd1 vssd1 vccd1 vccd1 _22725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_1_wb_clk_i clkbuf_3_2_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 INSDIODE2_358/DIODE
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_63_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16641_ _16641_/A vssd1 vssd1 vccd1 vccd1 _22468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13853_ _13056_/B _13836_/B _13746_/X vssd1 vssd1 vccd1 vccd1 _13853_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_406 _13880_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12804_ _13534_/A _13534_/B vssd1 vssd1 vccd1 vccd1 _15678_/A sky130_fd_sc_hd__nor2_2
XFILLER_16_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_417 _14054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19360_ _19360_/A vssd1 vssd1 vccd1 vccd1 _23341_/D sky130_fd_sc_hd__clkbuf_1
X_16572_ _16572_/A vssd1 vssd1 vccd1 vccd1 _22437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_428 _14521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13784_ _13821_/A _14006_/C vssd1 vssd1 vccd1 vccd1 _13830_/B sky130_fd_sc_hd__or2_1
XINSDIODE2_439 _23915_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_308_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18311_ _18314_/A _18314_/C _18292_/X vssd1 vssd1 vccd1 vccd1 _18311_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15523_ _19210_/A vssd1 vssd1 vccd1 vccd1 _15523_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _22473_/Q _22633_/Q _22312_/Q _23448_/Q _12733_/X _12734_/X vssd1 vssd1 vccd1
+ vccd1 _12735_/X sky130_fd_sc_hd__mux4_1
X_19291_ _19337_/S vssd1 vssd1 vccd1 vccd1 _19300_/S sky130_fd_sc_hd__buf_4
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _18242_/A vssd1 vssd1 vccd1 vccd1 _18242_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_231_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_337_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _13349_/A _13349_/B _13611_/A vssd1 vssd1 vccd1 vccd1 _13350_/A sky130_fd_sc_hd__a21oi_4
X_15454_ _13385_/Y _16131_/B _15453_/Y _13439_/A vssd1 vssd1 vccd1 vccd1 _15454_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_231_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11617_ _11890_/A vssd1 vssd1 vccd1 vccd1 _12117_/A sky130_fd_sc_hd__clkbuf_4
X_14405_ _14473_/A _14446_/B vssd1 vssd1 vccd1 vccd1 _14483_/A sky130_fd_sc_hd__or2_4
XFILLER_169_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18173_ _18187_/A _18167_/X _18195_/B _18118_/A vssd1 vssd1 vccd1 vccd1 _18173_/X
+ sky130_fd_sc_hd__o211a_1
X_15385_ _14953_/A _14949_/X _15385_/S vssd1 vssd1 vccd1 vccd1 _15386_/A sky130_fd_sc_hd__mux2_1
X_12597_ _11884_/B _21422_/A _12596_/Y vssd1 vssd1 vccd1 vccd1 _12602_/A sky130_fd_sc_hd__o21ai_4
XFILLER_317_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_345_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17124_ _17222_/B vssd1 vssd1 vccd1 vccd1 _17234_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_128_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11548_ _13073_/A _11548_/B vssd1 vssd1 vccd1 vccd1 _11548_/X sky130_fd_sc_hd__or2_1
X_14336_ _15084_/S _15192_/B _14848_/A vssd1 vssd1 vccd1 vccd1 _14336_/X sky130_fd_sc_hd__o21a_1
XFILLER_344_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_333_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17055_ _13923_/B _17054_/X _17087_/S vssd1 vssd1 vccd1 vccd1 _17055_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14267_ _14281_/A vssd1 vssd1 vccd1 vccd1 _14348_/A sky130_fd_sc_hd__buf_2
X_11479_ _22807_/Q _22775_/Q _22676_/Q _22743_/Q _21771_/A _15616_/A vssd1 vssd1 vccd1
+ vccd1 _11480_/B sky130_fd_sc_hd__mux4_1
XFILLER_171_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13218_ _13218_/A _13218_/B vssd1 vssd1 vccd1 vccd1 _13218_/X sky130_fd_sc_hd__or2_1
X_16006_ _15752_/X _16002_/X _16004_/Y _16005_/X vssd1 vssd1 vccd1 vccd1 _16006_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_315_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14198_ _14195_/X _14198_/B _14198_/C _14198_/D vssd1 vssd1 vccd1 vccd1 _14199_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_313_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _13149_/A _13149_/B vssd1 vssd1 vccd1 vccd1 _13149_/Y sky130_fd_sc_hd__nor2_1
XFILLER_286_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _22829_/Q _17956_/X _17939_/X input275/X _17951_/X vssd1 vssd1 vccd1 vccd1
+ _17957_/X sky130_fd_sc_hd__a221o_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16908_ _19258_/A vssd1 vssd1 vccd1 vccd1 _16908_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_254_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17888_ _14125_/Y _18191_/A _18018_/A vssd1 vssd1 vccd1 vccd1 _18021_/B sky130_fd_sc_hd__o21ai_4
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19627_ _19627_/A _19843_/A vssd1 vssd1 vccd1 vccd1 _19684_/A sky130_fd_sc_hd__or2_4
XFILLER_253_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16839_ _16838_/X _22528_/Q _16845_/S vssd1 vssd1 vccd1 vccd1 _16840_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19558_ _23429_/Q _19163_/A _19566_/S vssd1 vssd1 vccd1 vccd1 _19559_/A sky130_fd_sc_hd__mux2_1
XFILLER_253_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23507_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18509_ _22998_/Q _18518_/B vssd1 vssd1 vccd1 vccd1 _18509_/Y sky130_fd_sc_hd__nand2_1
XFILLER_202_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19489_ _19489_/A vssd1 vssd1 vccd1 vccd1 _23398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_278_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21520_ _21520_/A vssd1 vssd1 vccd1 vccd1 _21840_/A sky130_fd_sc_hd__buf_2
XFILLER_179_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21451_ _21451_/A _21451_/B vssd1 vssd1 vccd1 vccd1 _21454_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_308_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20402_ _20355_/A _20400_/Y _20174_/A vssd1 vssd1 vccd1 vccd1 _20402_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_193_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21382_ _21382_/A vssd1 vssd1 vccd1 vccd1 _21520_/A sky130_fd_sc_hd__buf_2
XFILLER_175_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_351_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23121_ _23537_/CLK _23121_/D vssd1 vssd1 vccd1 vccd1 _23121_/Q sky130_fd_sc_hd__dfxtp_1
X_20333_ _20333_/A vssd1 vssd1 vccd1 vccd1 _20333_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_324_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23052_ _23500_/CLK _23052_/D vssd1 vssd1 vccd1 vccd1 _23052_/Q sky130_fd_sc_hd__dfxtp_1
X_20264_ _20264_/A _20368_/B vssd1 vssd1 vccd1 vccd1 _20267_/B sky130_fd_sc_hd__or2_1
XFILLER_350_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_332_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22003_ _22003_/A _22224_/B vssd1 vssd1 vccd1 vccd1 _22003_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_289_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20195_ _20146_/X _20579_/A _20194_/X _18547_/X vssd1 vssd1 vccd1 vccd1 _23656_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_331_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput106 dout0[9] vssd1 vssd1 vccd1 vccd1 input106/X sky130_fd_sc_hd__buf_2
Xinput117 dout1[19] vssd1 vssd1 vccd1 vccd1 input117/X sky130_fd_sc_hd__clkbuf_1
XTAP_5328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput128 dout1[29] vssd1 vssd1 vccd1 vccd1 input128/X sky130_fd_sc_hd__clkbuf_1
XTAP_5339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput139 dout1[39] vssd1 vssd1 vccd1 vccd1 input139/X sky130_fd_sc_hd__clkbuf_2
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22905_ _22929_/CLK _22905_/D vssd1 vssd1 vccd1 vccd1 _22905_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23885_ _23888_/CLK _23885_/D vssd1 vssd1 vccd1 vccd1 _23885_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_186_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22836_ _23632_/CLK _22836_/D vssd1 vssd1 vccd1 vccd1 _22836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_260_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22767_ _22801_/CLK _22767_/D vssd1 vssd1 vccd1 vccd1 _22767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_347_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12520_ _23911_/Q _20499_/B _12520_/S vssd1 vssd1 vccd1 vccd1 _13359_/B sky130_fd_sc_hd__mux2_1
XFILLER_213_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21718_ _21716_/X _21717_/X _21598_/X vssd1 vssd1 vccd1 vccd1 _21718_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_40_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22698_ _23068_/CLK _22698_/D vssd1 vssd1 vccd1 vccd1 _22698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_297_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12463_/A _12451_/B vssd1 vssd1 vccd1 vccd1 _12451_/Y sky130_fd_sc_hd__nor2_1
XFILLER_338_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21649_ _21649_/A vssd1 vssd1 vccd1 vccd1 _21649_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11402_ _11402_/A vssd1 vssd1 vccd1 vccd1 _11403_/A sky130_fd_sc_hd__buf_2
XFILLER_327_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15170_ _15170_/A vssd1 vssd1 vccd1 vccd1 _22268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12382_ _22360_/Q _22392_/Q _22681_/Q _23048_/Q _12209_/X _12210_/X vssd1 vssd1 vccd1
+ vccd1 _12383_/B sky130_fd_sc_hd__mux4_1
XFILLER_326_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14121_ _22888_/Q _14110_/B _14121_/C _14121_/D vssd1 vssd1 vccd1 vccd1 _18018_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_299_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23319_ _23543_/CLK _23319_/D vssd1 vssd1 vccd1 vccd1 _23319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_327_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11333_ _11986_/A vssd1 vssd1 vccd1 vccd1 _12998_/A sky130_fd_sc_hd__buf_4
XFILLER_153_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_299_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14052_ _14064_/A _14052_/B _14052_/C vssd1 vssd1 vccd1 vccd1 _14052_/X sky130_fd_sc_hd__or3_1
XTAP_7220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11264_ _14371_/A _14371_/B _11263_/Y _13459_/A vssd1 vssd1 vccd1 vccd1 _11404_/B
+ sky130_fd_sc_hd__o211a_2
XTAP_7231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_7242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13003_ _22379_/Q _22411_/Q _22700_/Q _23067_/Q _11532_/A _11533_/A vssd1 vssd1 vccd1
+ vccd1 _13003_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18860_ _23136_/Q _18859_/X _18866_/S vssd1 vssd1 vccd1 vccd1 _18861_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XTAP_7275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11195_ _11195_/A vssd1 vssd1 vccd1 vccd1 _11196_/A sky130_fd_sc_hd__buf_6
XFILLER_122_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17811_ _22779_/Q _17553_/X _17815_/S vssd1 vssd1 vccd1 vccd1 _17812_/A sky130_fd_sc_hd__mux2_1
XTAP_6563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18791_ _18791_/A vssd1 vssd1 vccd1 vccd1 _23114_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17742_ _17742_/A vssd1 vssd1 vccd1 vccd1 _22748_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_294_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14954_ _14347_/X _14325_/X _15018_/S vssd1 vssd1 vccd1 vccd1 _14954_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_291_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13905_ _13933_/A _14085_/A vssd1 vssd1 vccd1 vccd1 _13905_/Y sky130_fd_sc_hd__nor2_4
XFILLER_63_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17673_ _17730_/S vssd1 vssd1 vccd1 vccd1 _17682_/S sky130_fd_sc_hd__buf_6
X_14885_ _17020_/A _21339_/B vssd1 vssd1 vccd1 vccd1 _14886_/B sky130_fd_sc_hd__and2_1
XFILLER_303_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19412_ _19468_/A vssd1 vssd1 vccd1 vccd1 _19481_/S sky130_fd_sc_hd__buf_6
XINSDIODE2_203 _19969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16624_ _16624_/A vssd1 vssd1 vccd1 vccd1 _22460_/D sky130_fd_sc_hd__clkbuf_1
X_13836_ _13836_/A _13836_/B vssd1 vssd1 vccd1 vccd1 _13836_/Y sky130_fd_sc_hd__nand2_1
XINSDIODE2_214 _14548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_225 _17052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_236 _15995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_247 _15408_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19343_ _19343_/A vssd1 vssd1 vccd1 vccd1 _23333_/D sky130_fd_sc_hd__clkbuf_1
X_16555_ _15240_/X _22430_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _16556_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_258 _21890_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13767_ _13807_/A _13767_/B vssd1 vssd1 vccd1 vccd1 _13767_/Y sky130_fd_sc_hd__nor2_1
XINSDIODE2_269 _18827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15506_ _23731_/Q _23861_/Q _16138_/S vssd1 vssd1 vccd1 vccd1 _15506_/X sky130_fd_sc_hd__mux2_1
XFILLER_349_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12718_ _23320_/Q _23288_/Q _23256_/Q _23544_/Q _12716_/X _12717_/X vssd1 vssd1 vccd1
+ vccd1 _12718_/X sky130_fd_sc_hd__mux4_2
XFILLER_241_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19274_ _19172_/X _23303_/Q _19278_/S vssd1 vssd1 vccd1 vccd1 _19275_/A sky130_fd_sc_hd__mux2_1
XFILLER_338_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16486_ _16486_/A vssd1 vssd1 vccd1 vccd1 _22400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13698_ _13765_/C vssd1 vssd1 vccd1 vccd1 _14089_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_309_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_321_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18225_ _22902_/Q _18227_/B vssd1 vssd1 vccd1 vccd1 _18225_/X sky130_fd_sc_hd__or2_1
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15437_ _22927_/Q vssd1 vssd1 vccd1 vccd1 _18305_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_175_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12649_ _12641_/Y _12643_/Y _12645_/Y _12648_/Y _11217_/A vssd1 vssd1 vccd1 vccd1
+ _12660_/B sky130_fd_sc_hd__o221a_1
XFILLER_176_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18156_ _18159_/A _18156_/B vssd1 vssd1 vccd1 vccd1 _18157_/A sky130_fd_sc_hd__and2_1
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15368_ _14804_/A _15330_/Y _15367_/Y _15162_/X vssd1 vssd1 vccd1 vccd1 _15368_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_345_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17107_ _17262_/A vssd1 vssd1 vccd1 vccd1 _17107_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14319_ _14316_/X _14651_/B _14664_/S vssd1 vssd1 vccd1 vccd1 _14319_/X sky130_fd_sc_hd__mux2_1
X_18087_ _22866_/Q _18082_/X _18083_/X _22999_/Q _18084_/X vssd1 vssd1 vccd1 vccd1
+ _18087_/X sky130_fd_sc_hd__a221o_1
XFILLER_183_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15299_ _22924_/Q _15299_/B vssd1 vssd1 vccd1 vccd1 _15299_/X sky130_fd_sc_hd__and2_1
XFILLER_132_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17038_ _17091_/A vssd1 vssd1 vccd1 vccd1 _17038_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_320_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_314_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_286_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18989_ _18989_/A vssd1 vssd1 vccd1 vccd1 _23191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20951_ _21916_/A _20950_/X _20695_/B _20940_/X vssd1 vssd1 vccd1 vccd1 _20951_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_66_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23670_ _23684_/CLK _23670_/D vssd1 vssd1 vccd1 vccd1 _23670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20882_ _20757_/B _20810_/A _20811_/A _23778_/Q vssd1 vssd1 vccd1 vccd1 _20883_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22621_ _23368_/CLK _22621_/D vssd1 vssd1 vccd1 vccd1 _22621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22552_ _23556_/CLK _22552_/D vssd1 vssd1 vccd1 vccd1 _22552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_356_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21503_ _21503_/A _21503_/B vssd1 vssd1 vccd1 vccd1 _21503_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_328_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22483_ _23585_/CLK _22483_/D vssd1 vssd1 vccd1 vccd1 _22483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21434_ _21401_/A _21404_/B _21400_/Y vssd1 vssd1 vccd1 vccd1 _21435_/B sky130_fd_sc_hd__o21a_1
XFILLER_355_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_308_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_324_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_323_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21365_ _14713_/A _21305_/X _21364_/Y _21281_/X vssd1 vssd1 vccd1 vccd1 _23913_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_352_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_324_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23104_ _23584_/CLK _23104_/D vssd1 vssd1 vccd1 vccd1 _23104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20316_ _20323_/A _21149_/A vssd1 vssd1 vccd1 vccd1 _20316_/Y sky130_fd_sc_hd__nand2_1
XFILLER_323_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21296_ _21293_/Y _21321_/B _21677_/A vssd1 vssd1 vccd1 vccd1 _21297_/D sky130_fd_sc_hd__a21oi_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_311_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_296_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23035_ _23419_/CLK _23035_/D vssd1 vssd1 vccd1 vccd1 _23035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_305_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20247_ _20213_/X _20622_/A _20245_/X _20246_/X vssd1 vssd1 vccd1 vccd1 _23662_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_304_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_324_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20178_ _23654_/Q _20165_/X _20177_/Y _18547_/X vssd1 vssd1 vccd1 vccd1 _23654_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_277_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_291_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11951_ _12754_/A _11951_/B vssd1 vssd1 vccd1 vccd1 _11951_/Y sky130_fd_sc_hd__nor2_1
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23937_ _23938_/CLK _23937_/D vssd1 vssd1 vccd1 vccd1 _23937_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_123_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ _15387_/S vssd1 vssd1 vccd1 vccd1 _14671_/S sky130_fd_sc_hd__buf_2
X_11882_ _11683_/A _11868_/X _11881_/Y _12634_/A vssd1 vssd1 vccd1 vccd1 _21596_/A
+ sky130_fd_sc_hd__a211o_4
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23868_ _23871_/CLK _23868_/D vssd1 vssd1 vccd1 vccd1 _23868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13621_ _13621_/A _13621_/B _13621_/C vssd1 vssd1 vccd1 vccd1 _13625_/B sky130_fd_sc_hd__nand3_4
X_22819_ _23551_/CLK _22819_/D vssd1 vssd1 vccd1 vccd1 _22819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23799_ _23942_/CLK _23799_/D vssd1 vssd1 vccd1 vccd1 _23799_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_60_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16340_ _15422_/X _22337_/Q _16344_/S vssd1 vssd1 vccd1 vccd1 _16341_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13552_ _13318_/A _13565_/A _13565_/B _13551_/X vssd1 vssd1 vccd1 vccd1 _13555_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_305_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12503_ _23461_/Q _23557_/Q _22521_/Q _22325_/Q _12501_/X _12502_/X vssd1 vssd1 vccd1
+ vccd1 _12503_/X sky130_fd_sc_hd__mux4_2
X_16271_ _18836_/A vssd1 vssd1 vccd1 vccd1 _16271_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13483_ _13570_/A _14820_/A _14821_/B vssd1 vssd1 vccd1 vccd1 _14206_/A sky130_fd_sc_hd__a21o_1
XFILLER_9_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18010_ _18018_/A vssd1 vssd1 vccd1 vccd1 _18118_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15222_ _15222_/A vssd1 vssd1 vccd1 vccd1 _15222_/X sky130_fd_sc_hd__buf_2
X_12434_ _22263_/Q _23079_/Q _23495_/Q _22424_/Q _11699_/A _11840_/A vssd1 vssd1 vccd1
+ vccd1 _12435_/B sky130_fd_sc_hd__mux4_1
XFILLER_328_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_327_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15153_ _22921_/Q vssd1 vssd1 vccd1 vccd1 _18286_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12365_ _12365_/A _12365_/B vssd1 vssd1 vccd1 vccd1 _12365_/Y sky130_fd_sc_hd__nor2_1
XFILLER_299_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_343_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14104_ _22893_/Q vssd1 vssd1 vccd1 vccd1 _18188_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_303_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11316_ _11800_/A vssd1 vssd1 vccd1 vccd1 _11317_/A sky130_fd_sc_hd__clkbuf_4
X_19961_ _23602_/Q _19957_/B _19960_/Y vssd1 vssd1 vccd1 vccd1 _23602_/D sky130_fd_sc_hd__o21a_1
X_15084_ _14627_/X _15083_/X _15084_/S vssd1 vssd1 vccd1 vccd1 _15252_/A sky130_fd_sc_hd__mux2_1
X_12296_ _22298_/Q _23434_/Q _12556_/A vssd1 vssd1 vccd1 vccd1 _12296_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_287_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18912_ _23157_/Q _18824_/X _18918_/S vssd1 vssd1 vccd1 vccd1 _18913_/A sky130_fd_sc_hd__mux2_1
XFILLER_314_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14035_ input219/X _14027_/X _14034_/X vssd1 vssd1 vccd1 vccd1 _14035_/X sky130_fd_sc_hd__a21o_4
XTAP_7050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11247_ _11247_/A vssd1 vssd1 vccd1 vccd1 _11247_/X sky130_fd_sc_hd__buf_4
XFILLER_180_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19892_ _16275_/X _23578_/Q _19898_/S vssd1 vssd1 vccd1 vccd1 _19893_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_351_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18843_ _18843_/A vssd1 vssd1 vccd1 vccd1 _18843_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11178_ _11961_/A vssd1 vssd1 vccd1 vccd1 _12130_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_311_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_267_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_310_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18774_ _23109_/Q _18769_/X _18786_/S vssd1 vssd1 vccd1 vccd1 _18775_/A sky130_fd_sc_hd__mux2_1
XTAP_5670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15986_ _23743_/Q _23873_/Q _16103_/S vssd1 vssd1 vccd1 vccd1 _15986_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17725_ _17725_/A vssd1 vssd1 vccd1 vccd1 _22741_/D sky130_fd_sc_hd__clkbuf_1
X_14937_ _15003_/A vssd1 vssd1 vccd1 vccd1 _14937_/X sky130_fd_sc_hd__buf_2
XFILLER_76_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17656_ _21185_/A vssd1 vssd1 vccd1 vccd1 _22254_/A sky130_fd_sc_hd__buf_8
X_14868_ _22917_/Q _14868_/B vssd1 vssd1 vccd1 vccd1 _14868_/X sky130_fd_sc_hd__and2_1
XFILLER_36_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16607_ _19267_/A _19555_/A vssd1 vssd1 vccd1 vccd1 _16664_/A sky130_fd_sc_hd__nor2_4
XFILLER_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13819_ _13893_/A vssd1 vssd1 vccd1 vccd1 _13861_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17587_ _17587_/A vssd1 vssd1 vccd1 vccd1 _22690_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14799_ _14682_/X _14757_/X _14759_/Y _14798_/Y vssd1 vssd1 vccd1 vccd1 _14799_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_259_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19326_ _19326_/A vssd1 vssd1 vccd1 vccd1 _23326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16538_ _14534_/X _22422_/Q _16546_/S vssd1 vssd1 vccd1 vccd1 _16539_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_337_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19257_ _19257_/A vssd1 vssd1 vccd1 vccd1 _23297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16469_ _14984_/X _22393_/Q _16469_/S vssd1 vssd1 vccd1 vccd1 _16470_/A sky130_fd_sc_hd__mux2_1
X_18208_ _22895_/Q _18214_/B vssd1 vssd1 vccd1 vccd1 _18208_/X sky130_fd_sc_hd__or2_1
XFILLER_339_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19188_ _19188_/A vssd1 vssd1 vccd1 vccd1 _19188_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_306_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_346_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_318_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_346_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18139_ _18139_/A vssd1 vssd1 vccd1 vccd1 _22884_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_318_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_306_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21150_ _21150_/A vssd1 vssd1 vccd1 vccd1 _21150_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_305_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_321_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_321_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20101_ _20790_/A vssd1 vssd1 vccd1 vccd1 _20101_/X sky130_fd_sc_hd__buf_12
X_21081_ _21081_/A _21308_/C vssd1 vssd1 vccd1 vccd1 _21301_/D sky130_fd_sc_hd__and2_2
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20032_ _23621_/Q _20040_/C _23622_/Q vssd1 vssd1 vccd1 vccd1 _20035_/B sky130_fd_sc_hd__a21oi_1
XFILLER_291_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_287_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21983_ _21975_/A _21714_/A _21967_/Y _21982_/X _18135_/X vssd1 vssd1 vccd1 vccd1
+ _23932_/D sky130_fd_sc_hd__o221a_1
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23722_ _23755_/CLK _23722_/D vssd1 vssd1 vccd1 vccd1 _23722_/Q sky130_fd_sc_hd__dfxtp_1
X_20934_ _20948_/A vssd1 vssd1 vccd1 vccd1 _20934_/X sky130_fd_sc_hd__buf_4
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23653_ _23700_/CLK _23653_/D vssd1 vssd1 vccd1 vccd1 _23653_/Q sky130_fd_sc_hd__dfxtp_1
X_20865_ _20865_/A vssd1 vssd1 vccd1 vccd1 _20865_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22604_ _23646_/CLK _22604_/D vssd1 vssd1 vccd1 vccd1 _22604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23584_ _23584_/CLK _23584_/D vssd1 vssd1 vccd1 vccd1 _23584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_356_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20796_ _20601_/B _20791_/X _20792_/X _23754_/Q vssd1 vssd1 vccd1 vccd1 _20797_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_329_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22535_ _23507_/CLK _22535_/D vssd1 vssd1 vccd1 vccd1 _22535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_356_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22466_ _23568_/CLK _22466_/D vssd1 vssd1 vccd1 vccd1 _22466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_356_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21417_ _21417_/A _21417_/B vssd1 vssd1 vccd1 vccd1 _21418_/B sky130_fd_sc_hd__xnor2_1
XFILLER_120_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22397_ _23565_/CLK _22397_/D vssd1 vssd1 vccd1 vccd1 _22397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12150_ _12007_/A _12149_/X _11631_/A vssd1 vssd1 vccd1 vccd1 _12150_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21348_ _23912_/Q _21348_/B vssd1 vssd1 vccd1 vccd1 _21348_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_351_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_335_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11101_ _16679_/A _22519_/Q vssd1 vssd1 vccd1 vccd1 _11102_/A sky130_fd_sc_hd__and2b_1
XFILLER_297_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12081_ _22274_/Q _23090_/Q _23506_/Q _22435_/Q _11700_/X _11839_/A vssd1 vssd1 vccd1
+ vccd1 _12082_/B sky130_fd_sc_hd__mux4_1
XFILLER_150_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21279_ _21076_/A _21199_/B _21278_/Y _21270_/X vssd1 vssd1 vccd1 vccd1 _23908_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23018_ _23466_/CLK _23018_/D vssd1 vssd1 vccd1 vccd1 _23018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_311_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ _23771_/Q _14911_/X _14913_/X _15838_/X _15839_/X vssd1 vssd1 vccd1 vccd1
+ _15840_/X sky130_fd_sc_hd__a221o_2
XFILLER_94_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_292_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _13322_/C _14793_/A _15770_/Y _13328_/A vssd1 vssd1 vccd1 vccd1 _15771_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_92_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12983_ _12983_/A _12983_/B vssd1 vssd1 vccd1 vccd1 _12983_/X sky130_fd_sc_hd__or2_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _22662_/Q _16259_/X _17516_/S vssd1 vssd1 vccd1 vccd1 _17511_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14722_ input160/X input125/X _14967_/S vssd1 vssd1 vccd1 vccd1 _14722_/X sky130_fd_sc_hd__mux2_8
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18490_ _18516_/A vssd1 vssd1 vccd1 vccd1 _18490_/X sky130_fd_sc_hd__buf_2
XFILLER_218_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _11275_/A _11924_/X _11933_/X _12156_/A vssd1 vssd1 vccd1 vccd1 _20234_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_233_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _22632_/Q _16265_/X _17443_/S vssd1 vssd1 vccd1 vccd1 _17442_/A sky130_fd_sc_hd__mux2_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14653_ _14653_/A vssd1 vssd1 vccd1 vccd1 _14653_/Y sky130_fd_sc_hd__inv_2
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _11914_/A _11865_/B vssd1 vssd1 vccd1 vccd1 _11865_/Y sky130_fd_sc_hd__nor2_1
XFILLER_261_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_107_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23583_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13604_ _13604_/A _13633_/A vssd1 vssd1 vccd1 vccd1 _13605_/B sky130_fd_sc_hd__nor2_2
X_17372_ _22606_/Q input200/X _17380_/S vssd1 vssd1 vccd1 vccd1 _17373_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14584_ _13706_/A _14572_/X _14577_/X _14583_/X vssd1 vssd1 vccd1 vccd1 _21204_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_32_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11796_ _12485_/A vssd1 vssd1 vccd1 vccd1 _12378_/A sky130_fd_sc_hd__buf_2
X_19111_ _23245_/Q _18798_/X _19113_/S vssd1 vssd1 vccd1 vccd1 _19112_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16323_ _16323_/A vssd1 vssd1 vccd1 vccd1 _22329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_319_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13535_ _13536_/A _13536_/B vssd1 vssd1 vccd1 vccd1 _13535_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19042_ _19088_/S vssd1 vssd1 vccd1 vccd1 _19051_/S sky130_fd_sc_hd__buf_4
XFILLER_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16254_ _16254_/A vssd1 vssd1 vccd1 vccd1 _22307_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_335_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13466_ _23946_/Q _23945_/Q vssd1 vssd1 vccd1 vccd1 _13467_/A sky130_fd_sc_hd__and2_1
XFILLER_328_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15205_ _15903_/B vssd1 vssd1 vccd1 vccd1 _15299_/B sky130_fd_sc_hd__buf_2
X_12417_ _12463_/A vssd1 vssd1 vccd1 vccd1 _12570_/A sky130_fd_sc_hd__buf_2
X_16185_ _14250_/A _13554_/A _16183_/X _16184_/Y vssd1 vssd1 vccd1 vccd1 _16186_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_154_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13397_ _13592_/A _13397_/B vssd1 vssd1 vccd1 vccd1 _13400_/C sky130_fd_sc_hd__xnor2_4
XFILLER_315_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15136_ _15136_/A vssd1 vssd1 vccd1 vccd1 _15136_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_303_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12348_ _12423_/A _12348_/B vssd1 vssd1 vccd1 vccd1 _12348_/Y sky130_fd_sc_hd__nand2_1
XFILLER_287_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19944_ _19950_/A _19944_/B vssd1 vssd1 vccd1 vccd1 _19944_/Y sky130_fd_sc_hd__nor2_1
X_12279_ _22460_/Q _22620_/Q _22299_/Q _23435_/Q _11455_/A _11733_/A vssd1 vssd1 vccd1
+ vccd1 _12279_/X sky130_fd_sc_hd__mux4_1
X_15067_ _15067_/A vssd1 vssd1 vccd1 vccd1 _15067_/X sky130_fd_sc_hd__buf_4
XFILLER_141_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_302_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_302_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14018_ _14012_/X _13722_/B _14013_/X input242/X vssd1 vssd1 vccd1 vccd1 _14018_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_296_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19875_ _19875_/A vssd1 vssd1 vccd1 vccd1 _23570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18826_ _18826_/A vssd1 vssd1 vccd1 vccd1 _23125_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_295_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18757_ _16899_/X _23103_/Q _18763_/S vssd1 vssd1 vccd1 vccd1 _18758_/A sky130_fd_sc_hd__mux2_1
XFILLER_209_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15969_ _21448_/B vssd1 vssd1 vccd1 vccd1 _21078_/B sky130_fd_sc_hd__buf_6
XFILLER_286_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17708_ _17708_/A vssd1 vssd1 vccd1 vccd1 _22733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18688_ _18688_/A vssd1 vssd1 vccd1 vccd1 _23072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17639_ _18865_/A vssd1 vssd1 vccd1 vccd1 _17639_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_208_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20650_ _15081_/A _20642_/X _20649_/X vssd1 vssd1 vccd1 vccd1 _20650_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_210_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_338_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19309_ _19223_/X _23319_/Q _19311_/S vssd1 vssd1 vccd1 vccd1 _19310_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20581_ _14196_/A _20773_/A _20574_/X vssd1 vssd1 vccd1 vccd1 _20581_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22320_ _23422_/CLK _22320_/D vssd1 vssd1 vccd1 vccd1 _22320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_286_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_338_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_325_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_307_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22251_ _14200_/Y _22253_/S _18268_/A vssd1 vssd1 vccd1 vccd1 _22251_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_353_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_293_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_307_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21202_ _21242_/A vssd1 vssd1 vccd1 vccd1 _21202_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22182_ _22182_/A _22182_/B vssd1 vssd1 vccd1 vccd1 _22183_/B sky130_fd_sc_hd__nand2_2
XFILLER_321_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21133_ _23861_/Q _21123_/X _21124_/X _20661_/A vssd1 vssd1 vccd1 vccd1 _21134_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_133_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21064_ _21177_/A _21064_/B vssd1 vssd1 vccd1 vccd1 _21064_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20015_ _20041_/A _20015_/B _20031_/C vssd1 vssd1 vccd1 vccd1 _23616_/D sky130_fd_sc_hd__nor3_1
XFILLER_286_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_321_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_5_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23563_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_234_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21966_ _23802_/Q _21683_/X _21965_/X _21660_/X vssd1 vssd1 vccd1 vccd1 _21967_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_261_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23705_ _23706_/CLK _23705_/D vssd1 vssd1 vccd1 vccd1 _23705_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_242_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20917_ _13931_/B _20908_/X _20613_/B _20912_/X vssd1 vssd1 vccd1 vccd1 _20917_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21897_ _17180_/X _21612_/X _21895_/X _21896_/X vssd1 vssd1 vccd1 vccd1 _23929_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_200_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23528_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_348_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11650_ _12216_/A vssd1 vssd1 vccd1 vccd1 _11651_/A sky130_fd_sc_hd__buf_2
X_23636_ _23637_/CLK _23636_/D vssd1 vssd1 vccd1 vccd1 _23636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20848_ _20695_/B _20846_/X _20847_/X _23768_/Q vssd1 vssd1 vccd1 vccd1 _20849_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11581_ _12291_/A vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__buf_2
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23567_ _23567_/CLK _23567_/D vssd1 vssd1 vccd1 vccd1 _23567_/Q sky130_fd_sc_hd__dfxtp_1
X_20779_ _20779_/A _20779_/B _20888_/C vssd1 vssd1 vccd1 vccd1 _20779_/X sky130_fd_sc_hd__or3_1
XFILLER_357_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13320_ _13403_/A _13403_/B _13319_/X vssd1 vssd1 vccd1 vccd1 _13321_/B sky130_fd_sc_hd__o21a_1
X_22518_ _23692_/CLK _22518_/D vssd1 vssd1 vccd1 vccd1 _22518_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23498_ _23530_/CLK _23498_/D vssd1 vssd1 vccd1 vccd1 _23498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_314_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_346_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22449_ _23584_/CLK _22449_/D vssd1 vssd1 vccd1 vccd1 _22449_/Q sky130_fd_sc_hd__dfxtp_1
X_13251_ _13399_/A _13239_/X _13250_/Y vssd1 vssd1 vccd1 vccd1 _13403_/A sky130_fd_sc_hd__a21oi_4
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12202_ _12189_/Y _12195_/Y _12198_/Y _12201_/Y _11242_/A vssd1 vssd1 vccd1 vccd1
+ _12203_/C sky130_fd_sc_hd__o221a_1
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_325_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_313_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13182_ _13117_/A _13181_/X _11352_/A vssd1 vssd1 vccd1 vccd1 _13182_/X sky130_fd_sc_hd__o21a_1
XFILLER_313_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_313_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12133_ _12126_/Y _12128_/Y _12130_/Y _12132_/Y _11244_/A vssd1 vssd1 vccd1 vccd1
+ _12134_/C sky130_fd_sc_hd__o221a_1
XFILLER_89_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_340_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ _18052_/A vssd1 vssd1 vccd1 vccd1 _17990_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_297_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16941_ _16941_/A _16941_/B vssd1 vssd1 vccd1 vccd1 _16943_/C sky130_fd_sc_hd__nor2_1
X_12064_ _12168_/A _12168_/B vssd1 vssd1 vccd1 vccd1 _15492_/S sky130_fd_sc_hd__and2b_2
XFILLER_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19660_ _19210_/X _23475_/Q _19660_/S vssd1 vssd1 vccd1 vccd1 _19661_/A sky130_fd_sc_hd__mux2_1
X_16872_ _16872_/A vssd1 vssd1 vccd1 vccd1 _22538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18611_ _16895_/X _23038_/Q _18619_/S vssd1 vssd1 vccd1 vccd1 _18612_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15823_ _19233_/A vssd1 vssd1 vccd1 vccd1 _15823_/X sky130_fd_sc_hd__buf_2
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19591_ _23444_/Q _19213_/A _19599_/S vssd1 vssd1 vccd1 vccd1 _19592_/A sky130_fd_sc_hd__mux2_1
XFILLER_253_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_292_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ _18542_/A vssd1 vssd1 vccd1 vccd1 _18542_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _15633_/X _15381_/Y _15578_/A vssd1 vssd1 vccd1 vccd1 _15754_/X sky130_fd_sc_hd__a21bo_2
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_90 _11627_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12966_ _13328_/A _13604_/A vssd1 vssd1 vccd1 vccd1 _13322_/C sky130_fd_sc_hd__or2_2
XFILLER_205_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _18776_/A vssd1 vssd1 vccd1 vccd1 _19169_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18473_ _22985_/Q _18478_/B vssd1 vssd1 vccd1 vccd1 _18473_/Y sky130_fd_sc_hd__nand2_1
XFILLER_233_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _22785_/Q _22753_/Q _22654_/Q _22721_/Q _11648_/A _11653_/A vssd1 vssd1 vccd1
+ vccd1 _11917_/X sky130_fd_sc_hd__mux4_1
X_15685_ _22964_/Q _16070_/A vssd1 vssd1 vccd1 vccd1 _15685_/X sky130_fd_sc_hd__or2_1
XFILLER_73_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _12897_/A _12897_/B vssd1 vssd1 vccd1 vccd1 _12897_/X sky130_fd_sc_hd__or2_1
XFILLER_221_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17424_ _22624_/Q _16239_/X _17432_/S vssd1 vssd1 vccd1 vccd1 _17425_/A sky130_fd_sc_hd__mux2_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14636_ _14633_/X _14634_/X _14845_/S vssd1 vssd1 vccd1 vccd1 _14636_/X sky130_fd_sc_hd__mux2_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11848_ _23310_/Q _23278_/Q _23246_/Q _23534_/Q _11770_/A _11621_/A vssd1 vssd1 vccd1
+ vccd1 _11849_/B sky130_fd_sc_hd__mux4_1
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _17355_/A vssd1 vssd1 vccd1 vccd1 _22598_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14567_ _16980_/A _14713_/C vssd1 vssd1 vccd1 vccd1 _14567_/Y sky130_fd_sc_hd__xnor2_2
X_11779_ _22787_/Q _22755_/Q _22656_/Q _22723_/Q _11595_/A _11566_/A vssd1 vssd1 vccd1
+ vccd1 _11779_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16306_ _18871_/A vssd1 vssd1 vccd1 vccd1 _16306_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_186_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13518_ _13518_/A _13518_/B vssd1 vssd1 vccd1 vccd1 _13518_/Y sky130_fd_sc_hd__nand2_1
XFILLER_347_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17286_ _22580_/Q _17255_/X _17240_/X _17285_/X vssd1 vssd1 vccd1 vccd1 _22580_/D
+ sky130_fd_sc_hd__a211o_1
X_14498_ _14748_/A vssd1 vssd1 vccd1 vccd1 _14498_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_335_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19025_ _16822_/X _23207_/Q _19029_/S vssd1 vssd1 vccd1 vccd1 _19026_/A sky130_fd_sc_hd__mux2_1
X_16237_ _22302_/Q _16236_/X _16237_/S vssd1 vssd1 vccd1 vccd1 _16238_/A sky130_fd_sc_hd__mux2_1
X_13449_ _23946_/Q _23945_/Q vssd1 vssd1 vccd1 vccd1 _13473_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_75_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23419_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_322_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16168_ _16168_/A _16168_/B vssd1 vssd1 vccd1 vccd1 _16168_/X sky130_fd_sc_hd__and2_1
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_318_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_318_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_303_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15119_ _15119_/A _15119_/B vssd1 vssd1 vccd1 vccd1 _15532_/A sky130_fd_sc_hd__and2_1
XFILLER_170_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_287_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16099_ _22943_/Q _14752_/X _14753_/X _22975_/Q vssd1 vssd1 vccd1 vccd1 _16099_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_330_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19927_ _23593_/Q _23592_/Q _19927_/C vssd1 vssd1 vccd1 vccd1 _19934_/C sky130_fd_sc_hd__and3_1
XFILLER_303_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19858_ _19858_/A vssd1 vssd1 vccd1 vccd1 _23562_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18809_ _23120_/Q _18808_/X _18818_/S vssd1 vssd1 vccd1 vccd1 _18810_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19789_ _23532_/Q _19188_/A _19793_/S vssd1 vssd1 vccd1 vccd1 _19790_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21820_ _21787_/A _21786_/B _21786_/A vssd1 vssd1 vccd1 vccd1 _21821_/B sky130_fd_sc_hd__o21ba_1
XFILLER_71_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21751_ _21724_/A _21727_/B _21724_/B vssd1 vssd1 vccd1 vccd1 _21752_/B sky130_fd_sc_hd__o21ba_2
XFILLER_70_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20702_ _20733_/A vssd1 vssd1 vccd1 vccd1 _20702_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_180_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21682_ _15329_/A _21479_/X _21664_/Y _21680_/X _21681_/X vssd1 vssd1 vccd1 vccd1
+ _23922_/D sky130_fd_sc_hd__o221a_1
XFILLER_52_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_339_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23421_ _23547_/CLK _23421_/D vssd1 vssd1 vccd1 vccd1 _23421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_260_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20633_ _14538_/X _20617_/X _20598_/X vssd1 vssd1 vccd1 vccd1 _20633_/X sky130_fd_sc_hd__a21o_1
XFILLER_354_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23352_ _23544_/CLK _23352_/D vssd1 vssd1 vccd1 vccd1 _23352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20564_ _20724_/A vssd1 vssd1 vccd1 vccd1 _20564_/X sky130_fd_sc_hd__buf_2
XFILLER_353_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22303_ _23047_/CLK _22303_/D vssd1 vssd1 vccd1 vccd1 _22303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23283_ _23510_/CLK _23283_/D vssd1 vssd1 vccd1 vccd1 _23283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_307_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20495_ _12493_/X _14567_/Y _21443_/A vssd1 vssd1 vccd1 vccd1 _21333_/B sky130_fd_sc_hd__mux2_1
XFILLER_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22234_ _22234_/A _22234_/B vssd1 vssd1 vccd1 vccd1 _22234_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22165_ _22165_/A _22171_/A vssd1 vssd1 vccd1 vccd1 _22167_/A sky130_fd_sc_hd__nor2_1
XTAP_6904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21116_ _23854_/Q _21110_/X _21111_/X _21013_/A vssd1 vssd1 vccd1 vccd1 _21117_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_160_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22096_ _20368_/A _21900_/B _16004_/B _22046_/X vssd1 vssd1 vccd1 vccd1 _22096_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_121_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21047_ _21047_/A vssd1 vssd1 vccd1 vccd1 _21047_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12820_ _22477_/Q _22637_/Q _12820_/S vssd1 vssd1 vccd1 vccd1 _12820_/X sky130_fd_sc_hd__mux2_1
XFILLER_234_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22998_ _23592_/CLK _22998_/D vssd1 vssd1 vccd1 vccd1 _22998_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_290_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _22472_/Q _22632_/Q _12751_/S vssd1 vssd1 vccd1 vccd1 _12751_/X sky130_fd_sc_hd__mux2_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21949_ _21949_/A _21954_/A vssd1 vssd1 vccd1 vccd1 _21951_/A sky130_fd_sc_hd__nand2_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _11702_/A vssd1 vssd1 vccd1 vccd1 _11703_/A sky130_fd_sc_hd__buf_4
XFILLER_70_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_349_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _21720_/A _15375_/X _15468_/Y _15469_/X vssd1 vssd1 vccd1 vccd1 _15470_/X
+ sky130_fd_sc_hd__a22o_2
X_12682_ _12926_/A _12682_/B vssd1 vssd1 vccd1 vccd1 _12682_/Y sky130_fd_sc_hd__nor2_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14421_ _21526_/A _14550_/A _14421_/S vssd1 vssd1 vccd1 vccd1 _14451_/B sky130_fd_sc_hd__mux2_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23619_ _23624_/CLK _23619_/D vssd1 vssd1 vccd1 vccd1 _23619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _12485_/A vssd1 vssd1 vccd1 vccd1 _12383_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_357_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17140_ _22567_/Q _17091_/X _17131_/X _17139_/X vssd1 vssd1 vccd1 vccd1 _22567_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_357_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14352_ _14635_/A vssd1 vssd1 vccd1 vccd1 _14665_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_168_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11564_ _12458_/A vssd1 vssd1 vccd1 vccd1 _11565_/A sky130_fd_sc_hd__buf_6
XFILLER_329_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ _13318_/A _13403_/A _13403_/B vssd1 vssd1 vccd1 vccd1 _13316_/A sky130_fd_sc_hd__or3_1
X_17071_ input77/X input105/X _17084_/S vssd1 vssd1 vccd1 vccd1 _17071_/X sky130_fd_sc_hd__mux2_8
XFILLER_317_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11495_ _11418_/X _11492_/X _11494_/X vssd1 vssd1 vccd1 vccd1 _11495_/Y sky130_fd_sc_hd__a21oi_1
X_14283_ _11557_/B _14791_/A _14343_/S vssd1 vssd1 vccd1 vccd1 _14283_/X sky130_fd_sc_hd__mux2_2
XFILLER_155_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16022_ _23744_/Q _23874_/Q _16022_/S vssd1 vssd1 vccd1 vccd1 _16022_/X sky130_fd_sc_hd__mux2_1
XFILLER_304_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13234_ _13214_/Y _20353_/A _13234_/S vssd1 vssd1 vccd1 vccd1 _13241_/A sky130_fd_sc_hd__mux2_2
XFILLER_344_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_298_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13165_ _23936_/Q vssd1 vssd1 vccd1 vccd1 _13165_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_313_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_312_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_298_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12116_ _23217_/Q _23185_/Q _23153_/Q _23121_/Q _12043_/S _11613_/X vssd1 vssd1 vccd1
+ vccd1 _12117_/B sky130_fd_sc_hd__mux4_1
XFILLER_111_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17973_ _22834_/Q _17972_/X _17959_/X input265/X _17966_/X vssd1 vssd1 vccd1 vccd1
+ _17973_/X sky130_fd_sc_hd__a221o_1
X_13096_ _13096_/A vssd1 vssd1 vccd1 vccd1 _13096_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_301_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12047_ _12047_/A _12047_/B vssd1 vssd1 vccd1 vccd1 _12047_/Y sky130_fd_sc_hd__nor2_1
X_16924_ _13662_/B _22421_/Q _17325_/B vssd1 vssd1 vccd1 vccd1 _17241_/B sky130_fd_sc_hd__and3b_2
X_19712_ _19769_/S vssd1 vssd1 vccd1 vccd1 _19721_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_238_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_193_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23496_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16855_ _16854_/X _22533_/Q _16861_/S vssd1 vssd1 vccd1 vccd1 _16856_/A sky130_fd_sc_hd__mux2_1
X_19643_ _19185_/X _23467_/Q _19649_/S vssd1 vssd1 vccd1 vccd1 _19644_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_322_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_122_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23624_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15806_ _23738_/Q _23868_/Q _15806_/S vssd1 vssd1 vccd1 vccd1 _15806_/X sky130_fd_sc_hd__mux2_1
XFILLER_219_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19574_ _19574_/A vssd1 vssd1 vccd1 vccd1 _23436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_253_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16786_ _16795_/A _16786_/B vssd1 vssd1 vccd1 vccd1 _16787_/A sky130_fd_sc_hd__or2_1
X_13998_ _14000_/A _14095_/A vssd1 vssd1 vccd1 vccd1 _13998_/Y sky130_fd_sc_hd__nor2_4
XFILLER_207_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18525_ _18520_/X _18524_/Y _18516_/X vssd1 vssd1 vccd1 vccd1 _23004_/D sky130_fd_sc_hd__a21oi_1
XFILLER_280_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15737_ _14592_/X _15725_/X _15736_/X vssd1 vssd1 vccd1 vccd1 _15738_/A sky130_fd_sc_hd__o21ai_4
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12949_ _12949_/A _12949_/B vssd1 vssd1 vccd1 vccd1 _12949_/X sky130_fd_sc_hd__or2_1
XFILLER_222_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18456_ _18476_/A vssd1 vssd1 vccd1 vccd1 _22260_/A sky130_fd_sc_hd__buf_6
XFILLER_244_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15668_ _19220_/A vssd1 vssd1 vccd1 vccd1 _15668_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_179_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17407_ _17407_/A vssd1 vssd1 vccd1 vccd1 _22616_/D sky130_fd_sc_hd__clkbuf_1
X_14619_ _14431_/X _14590_/X _14616_/X _14618_/X _14518_/X vssd1 vssd1 vccd1 vccd1
+ _14619_/X sky130_fd_sc_hd__o32a_4
X_18387_ _18403_/A _18392_/C vssd1 vssd1 vccd1 vccd1 _18387_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15599_ _23797_/Q _14742_/X _15067_/X vssd1 vssd1 vccd1 vccd1 _15599_/X sky130_fd_sc_hd__a21o_1
XFILLER_202_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17338_ _17882_/S vssd1 vssd1 vccd1 vccd1 _17347_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_187_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_336_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_335_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17269_ _17269_/A vssd1 vssd1 vccd1 vccd1 _17269_/Y sky130_fd_sc_hd__inv_2
X_19008_ _16902_/X _23200_/Q _19012_/S vssd1 vssd1 vccd1 vccd1 _19009_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_347_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20280_ _17134_/A _20295_/A _20279_/Y vssd1 vssd1 vccd1 vccd1 _20280_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_128_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_288_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_290_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_288_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22921_ _22923_/CLK _22921_/D vssd1 vssd1 vccd1 vccd1 _22921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22852_ _23426_/CLK _22852_/D vssd1 vssd1 vccd1 vccd1 _22852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21803_ _21803_/A _21803_/B vssd1 vssd1 vccd1 vccd1 _21804_/C sky130_fd_sc_hd__nand2_1
XFILLER_225_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22783_ _23369_/CLK _22783_/D vssd1 vssd1 vccd1 vccd1 _22783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21734_ _21734_/A _21734_/B vssd1 vssd1 vccd1 vccd1 _21734_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_224_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_358_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21665_ _23824_/Q _23758_/Q vssd1 vssd1 vccd1 vccd1 _21667_/A sky130_fd_sc_hd__or2_1
XFILLER_240_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23404_ _23950_/A _23404_/D vssd1 vssd1 vccd1 vccd1 _23404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20616_ _20616_/A _20631_/B vssd1 vssd1 vccd1 vccd1 _20620_/B sky130_fd_sc_hd__nor2_2
XFILLER_326_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21596_ _21596_/A _21716_/B vssd1 vssd1 vccd1 vccd1 _21596_/X sky130_fd_sc_hd__or2_1
XFILLER_177_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20547_ _20547_/A _20936_/A vssd1 vssd1 vccd1 vccd1 _20558_/A sky130_fd_sc_hd__nor2_2
X_23335_ _23367_/CLK _23335_/D vssd1 vssd1 vccd1 vccd1 _23335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_353_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11280_ _11280_/A vssd1 vssd1 vccd1 vccd1 _11818_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_125_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_326_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23266_ _23554_/CLK _23266_/D vssd1 vssd1 vccd1 vccd1 _23266_/Q sky130_fd_sc_hd__dfxtp_1
X_20478_ _23710_/Q _20487_/B vssd1 vssd1 vccd1 vccd1 _20478_/X sky130_fd_sc_hd__or2_1
XFILLER_342_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22217_ _22217_/A _22224_/A vssd1 vssd1 vccd1 vccd1 _22218_/B sky130_fd_sc_hd__nor2_1
X_23197_ _23419_/CLK _23197_/D vssd1 vssd1 vccd1 vccd1 _23197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22148_ _23841_/Q _23775_/Q vssd1 vssd1 vccd1 vccd1 _22148_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_350_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput390 _14057_/X vssd1 vssd1 vccd1 vccd1 din0[24] sky130_fd_sc_hd__buf_2
XFILLER_105_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14970_ _14961_/X _14969_/Y _14970_/S vssd1 vssd1 vccd1 vccd1 _14970_/X sky130_fd_sc_hd__mux2_4
X_22079_ _23838_/Q _23772_/Q vssd1 vssd1 vccd1 vccd1 _22081_/A sky130_fd_sc_hd__and2_1
XFILLER_0_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13921_ _23917_/Q vssd1 vssd1 vccd1 vccd1 _21500_/A sky130_fd_sc_hd__buf_2
XFILLER_247_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16640_ _22468_/Q _16252_/X _16640_/S vssd1 vssd1 vccd1 vccd1 _16641_/A sky130_fd_sc_hd__mux2_1
X_13852_ _13852_/A _13864_/B vssd1 vssd1 vccd1 vccd1 _13852_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12803_ _13534_/A _13534_/B vssd1 vssd1 vccd1 vccd1 _12805_/A sky130_fd_sc_hd__and2_2
XINSDIODE2_407 _13880_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16571_ _15570_/X _22437_/Q _16579_/S vssd1 vssd1 vccd1 vccd1 _16572_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13783_ _15576_/A vssd1 vssd1 vccd1 vccd1 _13821_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_418 _14054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_290_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_429 _22887_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18310_ _22929_/Q _18306_/C _18309_/Y vssd1 vssd1 vccd1 vccd1 _22929_/D sky130_fd_sc_hd__o21a_1
XFILLER_27_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15522_ _18817_/A vssd1 vssd1 vccd1 vccd1 _19210_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12734_/X sky130_fd_sc_hd__buf_4
XFILLER_203_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19290_ _19290_/A vssd1 vssd1 vccd1 vccd1 _23310_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _22860_/Q _18229_/X _18240_/X _18232_/X vssd1 vssd1 vccd1 vccd1 _22908_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_188_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _15453_/A _16131_/B vssd1 vssd1 vccd1 vccd1 _15453_/Y sky130_fd_sc_hd__nor2_1
X_12665_ _12665_/A _15582_/A vssd1 vssd1 vccd1 vccd1 _13611_/A sky130_fd_sc_hd__nor2_2
XFILLER_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_318_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14404_ _14457_/A _14404_/B vssd1 vssd1 vccd1 vccd1 _14446_/B sky130_fd_sc_hd__or2_2
X_18172_ _18172_/A _18171_/X vssd1 vssd1 vccd1 vccd1 _18195_/B sky130_fd_sc_hd__or2b_1
XFILLER_318_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11616_ _11834_/A vssd1 vssd1 vccd1 vccd1 _11890_/A sky130_fd_sc_hd__buf_4
XFILLER_30_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_329_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15384_ _15011_/A _14856_/Y _15253_/X vssd1 vssd1 vccd1 vccd1 _15384_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_318_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12596_ _17033_/A _12596_/B vssd1 vssd1 vccd1 vccd1 _12596_/Y sky130_fd_sc_hd__nand2_1
X_17123_ _23474_/Q _17113_/X _17114_/X _17094_/X _17122_/Y vssd1 vssd1 vccd1 vccd1
+ _17123_/X sky130_fd_sc_hd__a32o_1
X_14335_ _14325_/X _14333_/Y _15132_/S vssd1 vssd1 vccd1 vccd1 _15192_/B sky130_fd_sc_hd__mux2_4
X_11547_ _22806_/Q _22774_/Q _22675_/Q _22742_/Q _11543_/X _13276_/A vssd1 vssd1 vccd1
+ vccd1 _11548_/B sky130_fd_sc_hd__mux4_1
XFILLER_345_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_344_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17054_ _13440_/A _17053_/X _17144_/A vssd1 vssd1 vccd1 vccd1 _17054_/X sky130_fd_sc_hd__mux2_1
X_14266_ _20205_/A _20139_/A vssd1 vssd1 vccd1 vccd1 _14281_/A sky130_fd_sc_hd__nand2_4
X_11478_ _21848_/A _11477_/X _11288_/X vssd1 vssd1 vccd1 vccd1 _11478_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_326_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_344_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16005_ _16005_/A vssd1 vssd1 vccd1 vccd1 _16005_/X sky130_fd_sc_hd__clkbuf_2
X_13217_ _23229_/Q _23197_/Q _23165_/Q _23133_/Q _11517_/A _11527_/A vssd1 vssd1 vccd1
+ vccd1 _13218_/B sky130_fd_sc_hd__mux4_2
XFILLER_332_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14197_ _11068_/Y _11095_/C _20532_/A _14196_/Y _20532_/D vssd1 vssd1 vccd1 vccd1
+ _14198_/D sky130_fd_sc_hd__o41a_1
XFILLER_298_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13148_ _23230_/Q _23198_/Q _23166_/Q _23134_/Q _13190_/S _13096_/X vssd1 vssd1 vccd1
+ vccd1 _13149_/B sky130_fd_sc_hd__mux4_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17956_ _17956_/A vssd1 vssd1 vccd1 vccd1 _17956_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_285_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _13249_/A _14276_/B vssd1 vssd1 vccd1 vccd1 _13080_/A sky130_fd_sc_hd__nand2_1
XFILLER_257_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16907_ _16907_/A vssd1 vssd1 vccd1 vccd1 _22549_/D sky130_fd_sc_hd__clkbuf_1
X_17887_ _22883_/Q vssd1 vssd1 vccd1 vccd1 _18018_/A sky130_fd_sc_hd__buf_2
XFILLER_294_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_293_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19626_ _19626_/A vssd1 vssd1 vccd1 vccd1 _23460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16838_ _19188_/A vssd1 vssd1 vccd1 vccd1 _16838_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16769_ _16769_/A vssd1 vssd1 vccd1 vccd1 _22507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19557_ _19625_/S vssd1 vssd1 vccd1 vccd1 _19566_/S sky130_fd_sc_hd__buf_4
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18508_ _18521_/A vssd1 vssd1 vccd1 vccd1 _18518_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_222_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19488_ _19169_/X _23398_/Q _19494_/S vssd1 vssd1 vccd1 vccd1 _19489_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18439_ _22974_/Q _18440_/C _18438_/Y vssd1 vssd1 vccd1 vccd1 _22974_/D sky130_fd_sc_hd__o21a_1
XFILLER_278_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_90_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23581_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21450_ _21485_/A _21485_/B vssd1 vssd1 vccd1 vccd1 _21451_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20401_ _16179_/X _20169_/X _20400_/Y vssd1 vssd1 vccd1 vccd1 _20401_/X sky130_fd_sc_hd__a21o_1
XFILLER_358_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_309_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21381_ _22130_/B vssd1 vssd1 vccd1 vccd1 _21381_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_335_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23120_ _23474_/CLK _23120_/D vssd1 vssd1 vccd1 vccd1 _23120_/Q sky130_fd_sc_hd__dfxtp_1
X_20332_ _20272_/X _20700_/A _20331_/X _20324_/X vssd1 vssd1 vccd1 vccd1 _23673_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_190_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_351_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_323_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23051_ _23369_/CLK _23051_/D vssd1 vssd1 vccd1 vccd1 _23051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_323_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20263_ _20387_/B vssd1 vssd1 vccd1 vccd1 _20368_/B sky130_fd_sc_hd__clkbuf_1
XTAP_6008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22002_ _22002_/A _22002_/B vssd1 vssd1 vccd1 vccd1 _22002_/X sky130_fd_sc_hd__xor2_2
XFILLER_350_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20194_ _23656_/Q _20223_/B vssd1 vssd1 vccd1 vccd1 _20194_/X sky130_fd_sc_hd__or2_1
XFILLER_89_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_304_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput107 dout1[0] vssd1 vssd1 vccd1 vccd1 input107/X sky130_fd_sc_hd__clkbuf_1
XTAP_5329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput118 dout1[1] vssd1 vssd1 vccd1 vccd1 input118/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput129 dout1[2] vssd1 vssd1 vccd1 vccd1 input129/X sky130_fd_sc_hd__clkbuf_1
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22904_ _22929_/CLK _22904_/D vssd1 vssd1 vccd1 vccd1 _22904_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23884_ _23926_/CLK _23884_/D vssd1 vssd1 vccd1 vccd1 _23884_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22835_ _23632_/CLK _22835_/D vssd1 vssd1 vccd1 vccd1 _22835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_353_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22766_ _23068_/CLK _22766_/D vssd1 vssd1 vccd1 vccd1 _22766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21717_ _13432_/A _13432_/B _21517_/B _15431_/X vssd1 vssd1 vccd1 vccd1 _21717_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22697_ _23450_/CLK _22697_/D vssd1 vssd1 vccd1 vccd1 _22697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _23302_/Q _23270_/Q _23238_/Q _23526_/Q _12537_/S _12449_/X vssd1 vssd1 vccd1
+ vccd1 _12451_/B sky130_fd_sc_hd__mux4_2
X_21648_ _21648_/A _21716_/B vssd1 vssd1 vccd1 vccd1 _21649_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11401_ _11401_/A vssd1 vssd1 vccd1 vccd1 _11402_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_338_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12381_ _12374_/X _12376_/X _12378_/X _12380_/X _11375_/A vssd1 vssd1 vccd1 vccd1
+ _12391_/B sky130_fd_sc_hd__a221o_1
XFILLER_138_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_327_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21579_ _22093_/A _21579_/B vssd1 vssd1 vccd1 vccd1 _21579_/Y sky130_fd_sc_hd__nand2_1
XFILLER_326_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14120_ _17908_/A _18009_/C _22844_/Q vssd1 vssd1 vccd1 vccd1 _14120_/X sky130_fd_sc_hd__and3b_1
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23318_ _23542_/CLK _23318_/D vssd1 vssd1 vccd1 vccd1 _23318_/Q sky130_fd_sc_hd__dfxtp_1
X_11332_ _12105_/A vssd1 vssd1 vccd1 vccd1 _11986_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_165_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_338_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_354_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_354_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_330_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14051_ _14074_/B vssd1 vssd1 vccd1 vccd1 _14064_/A sky130_fd_sc_hd__clkbuf_1
XTAP_7210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23249_ _23537_/CLK _23249_/D vssd1 vssd1 vccd1 vccd1 _23249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11263_ _12345_/B _14132_/D _11382_/B _13412_/A vssd1 vssd1 vccd1 vccd1 _11263_/Y
+ sky130_fd_sc_hd__nand4_1
XTAP_7221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13002_ _13006_/A _13002_/B vssd1 vssd1 vccd1 vccd1 _13002_/X sky130_fd_sc_hd__or2_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_295_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11194_ _11584_/A vssd1 vssd1 vccd1 vccd1 _11195_/A sky130_fd_sc_hd__buf_4
XTAP_7265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17810_ _17810_/A vssd1 vssd1 vccd1 vccd1 _22778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18790_ _23114_/Q _18788_/X _18802_/S vssd1 vssd1 vccd1 vccd1 _18791_/A sky130_fd_sc_hd__mux2_1
XFILLER_294_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17741_ _22748_/Q _17556_/X _17743_/S vssd1 vssd1 vccd1 vccd1 _17742_/A sky130_fd_sc_hd__mux2_1
XTAP_5863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14953_ _14953_/A vssd1 vssd1 vccd1 vccd1 _14953_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_43_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13904_ _17020_/A _14865_/A _13931_/A vssd1 vssd1 vccd1 vccd1 _14085_/A sky130_fd_sc_hd__mux2_8
X_17672_ _17672_/A vssd1 vssd1 vccd1 vccd1 _22717_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14884_ _17020_/A _21339_/B vssd1 vssd1 vccd1 vccd1 _14976_/B sky130_fd_sc_hd__nor2_1
XFILLER_345_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19411_ _19699_/B _19483_/B vssd1 vssd1 vccd1 vccd1 _19468_/A sky130_fd_sc_hd__nor2_8
X_16623_ _22460_/Q _16227_/X _16629_/S vssd1 vssd1 vccd1 vccd1 _16624_/A sky130_fd_sc_hd__mux2_1
X_13835_ _13835_/A _13875_/C vssd1 vssd1 vccd1 vccd1 _13835_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_204 _19969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_215 _14619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_226 _17052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_237 _15995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16554_ _16554_/A vssd1 vssd1 vccd1 vccd1 _22429_/D sky130_fd_sc_hd__clkbuf_1
X_19342_ _23333_/Q _18769_/X _19350_/S vssd1 vssd1 vccd1 vccd1 _19343_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_248 _15408_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13766_ _13874_/A _13815_/B _13864_/A _13721_/B vssd1 vssd1 vccd1 vccd1 _13767_/B
+ sky130_fd_sc_hd__o22a_4
XFILLER_204_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_259 _21890_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_349_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15505_ _23667_/Q _16137_/B vssd1 vssd1 vccd1 vccd1 _15505_/X sky130_fd_sc_hd__or2_1
X_12717_ _12717_/A vssd1 vssd1 vccd1 vccd1 _12717_/X sky130_fd_sc_hd__buf_6
X_19273_ _19273_/A vssd1 vssd1 vccd1 vccd1 _23302_/D sky130_fd_sc_hd__clkbuf_1
X_16485_ _15372_/X _22400_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _16486_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13697_ _13697_/A vssd1 vssd1 vccd1 vccd1 _13697_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_349_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18224_ _22853_/Q _18216_/X _18223_/X _18219_/X vssd1 vssd1 vccd1 vccd1 _22901_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15436_ _15832_/A vssd1 vssd1 vccd1 vccd1 _15436_/X sky130_fd_sc_hd__clkbuf_2
XPHY_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12648_ _12759_/A _12647_/X _12687_/A vssd1 vssd1 vccd1 vccd1 _12648_/Y sky130_fd_sc_hd__o21ai_1
XPHY_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18155_ _14119_/B _22881_/Q _18158_/S vssd1 vssd1 vccd1 vccd1 _18156_/B sky130_fd_sc_hd__mux2_1
XFILLER_200_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_318_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15367_ _15367_/A _15367_/B vssd1 vssd1 vccd1 vccd1 _15367_/Y sky130_fd_sc_hd__nor2_1
XFILLER_306_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12579_ _12590_/A _12578_/X _11282_/A vssd1 vssd1 vccd1 vccd1 _12579_/X sky130_fd_sc_hd__o21a_1
XFILLER_346_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17106_ _15329_/A _17105_/X _17137_/S vssd1 vssd1 vccd1 vccd1 _17106_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_345_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_318_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14318_ _14369_/A vssd1 vssd1 vccd1 vccd1 _14664_/S sky130_fd_sc_hd__buf_2
XFILLER_332_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18086_ _22866_/Q _18081_/X _18085_/X _18075_/X vssd1 vssd1 vccd1 vccd1 _22866_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15298_ _14682_/X _15290_/X _15297_/X vssd1 vssd1 vccd1 vccd1 _15298_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_305_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17037_ _22557_/Q _16922_/X _17028_/X _17036_/X vssd1 vssd1 vccd1 vccd1 _22557_/D
+ sky130_fd_sc_hd__a211o_1
X_14249_ _14244_/X _14248_/Y _15830_/A vssd1 vssd1 vccd1 vccd1 _21199_/A sky130_fd_sc_hd__mux2_4
XFILLER_132_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_286_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_313_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18988_ _16873_/X _23191_/Q _18990_/S vssd1 vssd1 vccd1 vccd1 _18989_/A sky130_fd_sc_hd__mux2_1
XFILLER_286_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_301_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17939_ _17959_/A vssd1 vssd1 vccd1 vccd1 _17939_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20950_ _20966_/A vssd1 vssd1 vccd1 vccd1 _20950_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_242_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19609_ _19609_/A vssd1 vssd1 vccd1 vccd1 _23452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20881_ _20881_/A vssd1 vssd1 vccd1 vccd1 _21215_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22620_ _23563_/CLK _22620_/D vssd1 vssd1 vccd1 vccd1 _22620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_289_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22551_ _23459_/CLK _22551_/D vssd1 vssd1 vccd1 vccd1 _22551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21502_ _21472_/A _21468_/Y _21472_/C _21470_/B vssd1 vssd1 vccd1 vccd1 _21503_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_179_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_356_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22482_ _23585_/CLK _22482_/D vssd1 vssd1 vccd1 vccd1 _22482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21433_ _21472_/A _21432_/Y vssd1 vssd1 vccd1 vccd1 _21435_/A sky130_fd_sc_hd__or2b_1
XFILLER_148_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_324_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21364_ _21942_/A _21347_/X _21363_/X vssd1 vssd1 vccd1 vccd1 _21364_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_238_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23103_ _23551_/CLK _23103_/D vssd1 vssd1 vccd1 vccd1 _23103_/Q sky130_fd_sc_hd__dfxtp_1
X_20315_ _20174_/X _20312_/X _20313_/Y _20314_/Y _20147_/X vssd1 vssd1 vccd1 vccd1
+ _21149_/A sky130_fd_sc_hd__o32a_4
XFILLER_101_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21295_ _16936_/C _21295_/B vssd1 vssd1 vccd1 vccd1 _21321_/B sky130_fd_sc_hd__and2b_4
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_323_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_351_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23034_ _23354_/CLK _23034_/D vssd1 vssd1 vccd1 vccd1 _23034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_289_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20246_ _20324_/A vssd1 vssd1 vccd1 vccd1 _20246_/X sky130_fd_sc_hd__buf_2
XFILLER_150_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_332_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_324_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20177_ _20177_/A _20996_/A vssd1 vssd1 vccd1 vccd1 _20177_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_296_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_320_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_291_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11950_ _22792_/Q _22760_/Q _22661_/Q _22728_/Q _12675_/A _12746_/A vssd1 vssd1 vccd1
+ vccd1 _11951_/B sky130_fd_sc_hd__mux4_1
XFILLER_218_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23936_ _23936_/CLK _23936_/D vssd1 vssd1 vccd1 vccd1 _23936_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_340_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23867_ _23874_/CLK _23867_/D vssd1 vssd1 vccd1 vccd1 _23867_/Q sky130_fd_sc_hd__dfxtp_1
X_11881_ _11630_/A _11871_/X _11875_/X _11880_/X _11683_/A vssd1 vssd1 vccd1 vccd1
+ _11881_/Y sky130_fd_sc_hd__a311oi_2
XFILLER_264_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13620_ _23925_/Q _13587_/A _15479_/B _13451_/A vssd1 vssd1 vccd1 vccd1 _13963_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_22818_ _22822_/CLK _22818_/D vssd1 vssd1 vccd1 vccd1 _22818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23798_ _23942_/CLK _23798_/D vssd1 vssd1 vccd1 vccd1 _23798_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_201_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13551_ _11558_/B _16054_/A _11558_/A vssd1 vssd1 vccd1 vccd1 _13551_/X sky130_fd_sc_hd__o21ba_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22749_ _23054_/CLK _22749_/D vssd1 vssd1 vccd1 vccd1 _22749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12502_ _23895_/Q vssd1 vssd1 vccd1 vccd1 _12502_/X sky130_fd_sc_hd__buf_2
X_16270_ _16270_/A vssd1 vssd1 vccd1 vccd1 _22312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_347_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13482_ _23946_/Q _20530_/B vssd1 vssd1 vccd1 vccd1 _14821_/B sky130_fd_sc_hd__nand2_2
XFILLER_41_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15221_ _23757_/Q _15215_/X _15216_/X _15218_/X _15220_/X vssd1 vssd1 vccd1 vccd1
+ _15221_/X sky130_fd_sc_hd__a221o_1
XFILLER_157_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12433_ _12421_/A _12432_/X _11844_/A vssd1 vssd1 vccd1 vccd1 _12433_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_200_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15152_ _22953_/Q _15151_/Y _15360_/A vssd1 vssd1 vccd1 vccd1 _15152_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12364_ _22264_/Q _23080_/Q _23496_/Q _22425_/Q _11413_/A _12425_/A vssd1 vssd1 vccd1
+ vccd1 _12365_/B sky130_fd_sc_hd__mux4_2
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14103_ _18187_/A vssd1 vssd1 vccd1 vccd1 _18126_/S sky130_fd_sc_hd__clkbuf_2
X_11315_ _11815_/A vssd1 vssd1 vccd1 vccd1 _11800_/A sky130_fd_sc_hd__buf_6
XFILLER_343_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19960_ _19981_/A _19960_/B vssd1 vssd1 vccd1 vccd1 _19960_/Y sky130_fd_sc_hd__nor2_1
X_15083_ _14778_/A _14772_/X _15129_/S vssd1 vssd1 vccd1 vccd1 _15083_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12295_ _22459_/Q _22619_/Q _12554_/S vssd1 vssd1 vccd1 vccd1 _12295_/X sky130_fd_sc_hd__mux2_1
X_18911_ _18911_/A vssd1 vssd1 vccd1 vccd1 _23156_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_268_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14034_ _13767_/B _14049_/A vssd1 vssd1 vccd1 vccd1 _14034_/X sky130_fd_sc_hd__and2b_1
XTAP_7040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_302_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11246_ _11246_/A vssd1 vssd1 vccd1 vccd1 _11247_/A sky130_fd_sc_hd__buf_6
XTAP_7051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19891_ _19891_/A vssd1 vssd1 vccd1 vccd1 _23577_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_351_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18842_ _18842_/A vssd1 vssd1 vccd1 vccd1 _23130_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11177_ _12082_/A vssd1 vssd1 vccd1 vccd1 _11961_/A sky130_fd_sc_hd__clkbuf_4
XTAP_6361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18773_ _18872_/S vssd1 vssd1 vccd1 vccd1 _18786_/S sky130_fd_sc_hd__buf_6
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15985_ _23679_/Q _15985_/B vssd1 vssd1 vccd1 vccd1 _15985_/X sky130_fd_sc_hd__or2_2
XFILLER_295_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14936_ _14936_/A vssd1 vssd1 vccd1 vccd1 _15003_/A sky130_fd_sc_hd__clkbuf_4
X_17724_ _22741_/Q _17636_/X _17726_/S vssd1 vssd1 vccd1 vccd1 _17725_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23588_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_180_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17655_ _17655_/A _17655_/B vssd1 vssd1 vccd1 vccd1 _17655_/Y sky130_fd_sc_hd__nand2_1
X_14867_ _13367_/D _14940_/B _14865_/Y _15010_/A vssd1 vssd1 vccd1 vccd1 _14867_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_90_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16606_ _16606_/A vssd1 vssd1 vccd1 vccd1 _22453_/D sky130_fd_sc_hd__clkbuf_1
X_13818_ _13818_/A vssd1 vssd1 vccd1 vccd1 _13818_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_223_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17586_ _22690_/Q _17585_/X _17592_/S vssd1 vssd1 vccd1 vccd1 _17587_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14798_ _14794_/A _14761_/X _14770_/Y _14797_/Y vssd1 vssd1 vccd1 vccd1 _14798_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_211_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19325_ _19245_/X _23326_/Q _19333_/S vssd1 vssd1 vccd1 vccd1 _19326_/A sky130_fd_sc_hd__mux2_1
X_16537_ _16605_/S vssd1 vssd1 vccd1 vccd1 _16546_/S sky130_fd_sc_hd__buf_8
XFILLER_73_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13749_ _14216_/A vssd1 vssd1 vccd1 vccd1 _15576_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19256_ _19255_/X _23297_/Q _19259_/S vssd1 vssd1 vccd1 vccd1 _19257_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16468_ _16468_/A vssd1 vssd1 vccd1 vccd1 _22392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18207_ hold1/X _18202_/X _18205_/X _18206_/X vssd1 vssd1 vccd1 vccd1 _22894_/D sky130_fd_sc_hd__o211a_1
X_15419_ _15519_/A vssd1 vssd1 vccd1 vccd1 _15708_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_192_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19187_ _19187_/A vssd1 vssd1 vccd1 vccd1 _23275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16399_ _15044_/X _22362_/Q _16407_/S vssd1 vssd1 vccd1 vccd1 _16400_/A sky130_fd_sc_hd__mux2_1
XFILLER_339_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18138_ _18138_/A _22122_/A vssd1 vssd1 vccd1 vccd1 _18139_/A sky130_fd_sc_hd__and2_1
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_345_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18069_ _18099_/A vssd1 vssd1 vccd1 vccd1 _18069_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20100_ _20120_/A _20100_/B _20106_/A vssd1 vssd1 vccd1 vccd1 _23640_/D sky130_fd_sc_hd__nor3_1
XFILLER_305_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21080_ _21080_/A _21080_/B vssd1 vssd1 vccd1 vccd1 _21308_/C sky130_fd_sc_hd__nor2_2
XFILLER_299_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_320_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20031_ _23620_/Q _23619_/Q _20031_/C _20031_/D vssd1 vssd1 vccd1 vccd1 _20040_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_258_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_286_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_302_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_301_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21982_ _21377_/X _21973_/X _21981_/Y vssd1 vssd1 vccd1 vccd1 _21982_/X sky130_fd_sc_hd__a21o_1
XFILLER_261_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23721_ _23856_/CLK _23721_/D vssd1 vssd1 vccd1 vccd1 _23721_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_328_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20933_ _21737_/A _20922_/X _20658_/B _20926_/X vssd1 vssd1 vccd1 vccd1 _20933_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23652_ _23652_/CLK _23652_/D vssd1 vssd1 vccd1 vccd1 _23652_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20864_ _20864_/A vssd1 vssd1 vccd1 vccd1 _20864_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_263_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22603_ _23649_/CLK _22603_/D vssd1 vssd1 vccd1 vccd1 _22603_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_53_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23583_ _23583_/CLK _23583_/D vssd1 vssd1 vccd1 vccd1 _23583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20795_ _20795_/A vssd1 vssd1 vccd1 vccd1 _23753_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22534_ _23503_/CLK _22534_/D vssd1 vssd1 vccd1 vccd1 _22534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_319_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22465_ _23568_/CLK _22465_/D vssd1 vssd1 vccd1 vccd1 _22465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_337_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_325_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_309_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21416_ _21416_/A _21415_/Y vssd1 vssd1 vccd1 vccd1 _21417_/B sky130_fd_sc_hd__or2b_1
XFILLER_5_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22396_ _23500_/CLK _22396_/D vssd1 vssd1 vccd1 vccd1 _22396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21347_ _23783_/Q _21814_/B _21345_/X _21346_/X vssd1 vssd1 vccd1 vccd1 _21347_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_163_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_352_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_311_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11100_ _22520_/Q vssd1 vssd1 vccd1 vccd1 _16679_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_296_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12080_ _11582_/A _12079_/X _11780_/X vssd1 vssd1 vccd1 vccd1 _12080_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21278_ _21278_/A _21283_/B vssd1 vssd1 vccd1 vccd1 _21278_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23017_ _23560_/CLK _23017_/D vssd1 vssd1 vccd1 vccd1 _23017_/Q sky130_fd_sc_hd__dfxtp_1
X_20229_ _15155_/X _20154_/X _20228_/Y vssd1 vssd1 vccd1 vccd1 _20229_/X sky130_fd_sc_hd__a21bo_1
XFILLER_270_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_292_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15770_ _13604_/A _15460_/B _14259_/A vssd1 vssd1 vccd1 vccd1 _15770_/Y sky130_fd_sc_hd__a21oi_1
X_12982_ _22379_/Q _22411_/Q _22700_/Q _23067_/Q _12820_/S _12749_/A vssd1 vssd1 vccd1
+ vccd1 _12983_/B sky130_fd_sc_hd__mux4_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _13789_/A _15286_/A _14720_/Y _15113_/A _15180_/A vssd1 vssd1 vccd1 vccd1
+ _14721_/X sky130_fd_sc_hd__o221a_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _11284_/A _11926_/X _11928_/X _11932_/X _11826_/A vssd1 vssd1 vccd1 vccd1
+ _11933_/X sky130_fd_sc_hd__a311o_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23919_ _23935_/CLK _23919_/D vssd1 vssd1 vccd1 vccd1 _23919_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_206_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _17440_/A vssd1 vssd1 vccd1 vccd1 _22631_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _14660_/S _14320_/X _14651_/Y vssd1 vssd1 vccd1 vccd1 _14653_/A sky130_fd_sc_hd__a21oi_4
XFILLER_45_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _23310_/Q _23278_/Q _23246_/Q _23534_/Q _11648_/A _11653_/A vssd1 vssd1 vccd1
+ vccd1 _11865_/B sky130_fd_sc_hd__mux4_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13603_ _13603_/A vssd1 vssd1 vccd1 vccd1 _13603_/X sky130_fd_sc_hd__buf_4
XFILLER_26_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _17371_/A vssd1 vssd1 vccd1 vccd1 _17380_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14583_ _15113_/A _14580_/Y _15244_/A _13789_/A _13706_/A vssd1 vssd1 vccd1 vccd1
+ _14583_/X sky130_fd_sc_hd__o221a_1
XFILLER_232_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11795_ _12135_/A _13752_/A _11794_/X vssd1 vssd1 vccd1 vccd1 _11939_/A sky130_fd_sc_hd__a21oi_2
XFILLER_25_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_347_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19110_ _19110_/A vssd1 vssd1 vccd1 vccd1 _23244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16322_ _14984_/X _22329_/Q _16322_/S vssd1 vssd1 vccd1 vccd1 _16323_/A sky130_fd_sc_hd__mux2_1
XFILLER_347_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13534_ _13534_/A _13534_/B vssd1 vssd1 vccd1 vccd1 _13534_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_319_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19041_ _19041_/A vssd1 vssd1 vccd1 vccd1 _23214_/D sky130_fd_sc_hd__clkbuf_1
X_16253_ _22307_/Q _16252_/X _16253_/S vssd1 vssd1 vccd1 vccd1 _16254_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13465_ _16980_/A _13587_/A _13476_/A _13473_/B vssd1 vssd1 vccd1 vccd1 _14216_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_201_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15204_ _14839_/X _15194_/X _15199_/X _15203_/Y vssd1 vssd1 vccd1 vccd1 _15204_/X
+ sky130_fd_sc_hd__o211a_2
X_12416_ _14791_/A vssd1 vssd1 vccd1 vccd1 _13364_/A sky130_fd_sc_hd__clkinv_4
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16184_ _14762_/A _14367_/X _14382_/X _15455_/A vssd1 vssd1 vccd1 vccd1 _16184_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_138_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_327_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13396_ _13323_/A _13601_/A _13027_/X vssd1 vssd1 vccd1 vccd1 _13397_/B sky130_fd_sc_hd__o21ai_2
XFILLER_343_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_315_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15135_ _15084_/S _15132_/X _15133_/Y _15134_/X vssd1 vssd1 vccd1 vccd1 _15136_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_342_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12347_ _22457_/Q _22617_/Q _12349_/S vssd1 vssd1 vccd1 vccd1 _12348_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_342_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19943_ _19975_/D _19971_/B vssd1 vssd1 vccd1 vccd1 _19944_/B sky130_fd_sc_hd__and2_1
XFILLER_299_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15066_ _23819_/Q _15066_/B _20986_/A vssd1 vssd1 vccd1 vccd1 _15066_/X sky130_fd_sc_hd__or3_1
X_12278_ _12410_/A _12278_/B vssd1 vssd1 vccd1 vccd1 _12278_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14017_ _13715_/A _14083_/A _13810_/B _14058_/A input241/X vssd1 vssd1 vccd1 vccd1
+ _14017_/X sky130_fd_sc_hd__a32o_4
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11229_ _11229_/A vssd1 vssd1 vccd1 vccd1 _11230_/A sky130_fd_sc_hd__buf_4
X_19874_ _16249_/X _23570_/Q _19876_/S vssd1 vssd1 vccd1 vccd1 _19875_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18825_ _23125_/Q _18824_/X _18834_/S vssd1 vssd1 vccd1 vccd1 _18826_/A sky130_fd_sc_hd__mux2_1
XTAP_6180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_295_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18756_ _18756_/A vssd1 vssd1 vccd1 vccd1 _23102_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15968_ _14987_/B _13575_/B _15574_/X _15967_/X vssd1 vssd1 vccd1 vccd1 _15968_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_271_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17707_ _22733_/Q _17610_/X _17715_/S vssd1 vssd1 vccd1 vccd1 _17708_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14919_ _14919_/A vssd1 vssd1 vccd1 vccd1 _14919_/X sky130_fd_sc_hd__buf_2
X_18687_ _23072_/Q _17633_/X _18691_/S vssd1 vssd1 vccd1 vccd1 _18688_/A sky130_fd_sc_hd__mux2_1
X_15899_ _15898_/X _22284_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15900_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17638_ _17638_/A vssd1 vssd1 vccd1 vccd1 _22706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17569_ _18795_/A vssd1 vssd1 vccd1 vccd1 _17569_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_210_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_338_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19308_ _19308_/A vssd1 vssd1 vccd1 vccd1 _23318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20580_ _20580_/A _20891_/A vssd1 vssd1 vccd1 vccd1 _20583_/B sky130_fd_sc_hd__nor2_2
XFILLER_149_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19239_ _19239_/A vssd1 vssd1 vccd1 vccd1 _19239_/X sky130_fd_sc_hd__buf_2
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22250_ _22246_/Y _22257_/A _22249_/X _21297_/C vssd1 vssd1 vccd1 vccd1 _22253_/S
+ sky130_fd_sc_hd__a31o_1
XFILLER_306_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21201_ _21214_/S vssd1 vssd1 vccd1 vccd1 _21242_/A sky130_fd_sc_hd__buf_2
X_22181_ _22205_/A _22181_/B vssd1 vssd1 vccd1 vccd1 _22182_/B sky130_fd_sc_hd__or2_1
XFILLER_191_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21132_ _21134_/A _21132_/B vssd1 vssd1 vccd1 vccd1 _23860_/D sky130_fd_sc_hd__nor2_1
XFILLER_133_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21063_ _23840_/Q vssd1 vssd1 vccd1 vccd1 _22151_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_302_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20014_ _23616_/Q _23615_/Q _20014_/C _20014_/D vssd1 vssd1 vccd1 vccd1 _20031_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_274_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_287_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_301_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21965_ _22038_/B _21965_/B vssd1 vssd1 vccd1 vccd1 _21965_/X sky130_fd_sc_hd__xor2_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23704_ _23704_/CLK _23704_/D vssd1 vssd1 vccd1 vccd1 _23704_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20916_ _23787_/Q _20911_/X _20915_/X _20906_/X vssd1 vssd1 vccd1 vccd1 _23787_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21896_ _22122_/A vssd1 vssd1 vccd1 vccd1 _21896_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23635_ _23637_/CLK _23635_/D vssd1 vssd1 vccd1 vccd1 _23635_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20847_ _20865_/A vssd1 vssd1 vccd1 vccd1 _20847_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_357_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23566_ _23566_/CLK _23566_/D vssd1 vssd1 vccd1 vccd1 _23566_/Q sky130_fd_sc_hd__dfxtp_1
X_11580_ _12421_/A vssd1 vssd1 vccd1 vccd1 _12291_/A sky130_fd_sc_hd__buf_4
XFILLER_356_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20778_ _23749_/Q _20786_/B _20777_/X _20763_/X vssd1 vssd1 vccd1 vccd1 _23749_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_211_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_357_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22517_ _23700_/CLK _22517_/D vssd1 vssd1 vccd1 vccd1 _22517_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_356_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23497_ _23529_/CLK _23497_/D vssd1 vssd1 vccd1 vccd1 _23497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13250_ _13561_/A _13247_/Y _13249_/Y vssd1 vssd1 vccd1 vccd1 _13250_/Y sky130_fd_sc_hd__o21ai_1
X_22448_ _23551_/CLK _22448_/D vssd1 vssd1 vccd1 vccd1 _22448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12201_ _12307_/A _12201_/B vssd1 vssd1 vccd1 vccd1 _12201_/Y sky130_fd_sc_hd__nor2_1
X_13181_ _22479_/Q _22639_/Q _22318_/Q _23454_/Q _11543_/A _13127_/X vssd1 vssd1 vccd1
+ vccd1 _13181_/X sky130_fd_sc_hd__mux4_2
XFILLER_159_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_324_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22379_ _23451_/CLK _22379_/D vssd1 vssd1 vccd1 vccd1 _22379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_325_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_313_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12132_ _12117_/A _12131_/X _11965_/A vssd1 vssd1 vccd1 vccd1 _12132_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_108_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16940_ _22712_/Q vssd1 vssd1 vccd1 vccd1 _16940_/X sky130_fd_sc_hd__buf_4
XFILLER_150_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12063_ _12168_/B _12168_/A vssd1 vssd1 vccd1 vccd1 _12065_/A sky130_fd_sc_hd__and2b_1
XFILLER_2_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16871_ _16870_/X _22538_/Q _16877_/S vssd1 vssd1 vccd1 vccd1 _16872_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18610_ _18610_/A vssd1 vssd1 vccd1 vccd1 _18619_/S sky130_fd_sc_hd__buf_4
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_293_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15822_ _18840_/A vssd1 vssd1 vccd1 vccd1 _19233_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_237_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19590_ _19612_/A vssd1 vssd1 vccd1 vccd1 _19599_/S sky130_fd_sc_hd__buf_4
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18541_ _18549_/A _18549_/B _23010_/Q _18098_/A _18550_/C vssd1 vssd1 vccd1 vccd1
+ _18542_/A sky130_fd_sc_hd__o41a_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15753_ _15753_/A _15790_/C vssd1 vssd1 vccd1 vccd1 _15753_/Y sky130_fd_sc_hd__xnor2_4
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12965_ _12965_/A vssd1 vssd1 vccd1 vccd1 _13604_/A sky130_fd_sc_hd__buf_2
XINSDIODE2_80 _21771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_91 _11627_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11916_ _12097_/A _11916_/B vssd1 vssd1 vccd1 vccd1 _11916_/X sky130_fd_sc_hd__or2_1
X_14704_ _12494_/X _14530_/X _14699_/X _21348_/B _14703_/X vssd1 vssd1 vccd1 vccd1
+ _18776_/A sky130_fd_sc_hd__a32o_4
X_18472_ _18467_/X _18471_/Y _18463_/X vssd1 vssd1 vccd1 vccd1 _22984_/D sky130_fd_sc_hd__a21oi_1
X_15684_ _22932_/Q _15000_/X _15001_/X _22964_/Q vssd1 vssd1 vccd1 vccd1 _15684_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_233_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _23226_/Q _23194_/Q _23162_/Q _23130_/Q _12792_/X _12793_/X vssd1 vssd1 vccd1
+ vccd1 _12897_/B sky130_fd_sc_hd__mux4_2
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _17469_/S vssd1 vssd1 vccd1 vccd1 _17432_/S sky130_fd_sc_hd__buf_4
X_14635_ _14635_/A vssd1 vssd1 vccd1 vccd1 _14845_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11847_ _11780_/X _11832_/Y _11834_/Y _11846_/X _11215_/A vssd1 vssd1 vccd1 vccd1
+ _11857_/B sky130_fd_sc_hd__o311a_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _22598_/Q input192/X _17358_/S vssd1 vssd1 vccd1 vccd1 _17355_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _14568_/A vssd1 vssd1 vccd1 vccd1 _14804_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_347_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11778_ _11949_/A _11778_/B vssd1 vssd1 vccd1 vccd1 _11778_/Y sky130_fd_sc_hd__nand2_1
X_16305_ _16305_/A vssd1 vssd1 vccd1 vccd1 _22323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13517_ _12234_/X _12287_/A _13516_/X _12236_/B vssd1 vssd1 vccd1 vccd1 _13935_/C
+ sky130_fd_sc_hd__o31ai_2
X_17285_ _17242_/X _17277_/X _17284_/X _17237_/X vssd1 vssd1 vccd1 vccd1 _17285_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_158_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14497_ _14497_/A vssd1 vssd1 vccd1 vccd1 _14748_/A sky130_fd_sc_hd__buf_2
XFILLER_159_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_307_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19024_ _19024_/A vssd1 vssd1 vccd1 vccd1 _23206_/D sky130_fd_sc_hd__clkbuf_1
X_16236_ _18801_/A vssd1 vssd1 vccd1 vccd1 _16236_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13448_ _23905_/Q _21448_/B _13448_/C vssd1 vssd1 vccd1 vccd1 _14175_/B sky130_fd_sc_hd__or3_2
XFILLER_316_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_316_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16167_ _22945_/Q vssd1 vssd1 vccd1 vccd1 _16168_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13379_ _13373_/X _13379_/B _13379_/C vssd1 vssd1 vccd1 vccd1 _13386_/B sky130_fd_sc_hd__nand3b_1
XFILLER_331_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15118_ _22510_/Q _13688_/A _14235_/A _15117_/X vssd1 vssd1 vccd1 vccd1 _15119_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
X_16098_ _14384_/X _14790_/X _16096_/X _16097_/X vssd1 vssd1 vccd1 vccd1 _16098_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_336_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_336_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_287_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19926_ _19926_/A _19926_/B vssd1 vssd1 vccd1 vccd1 _23592_/D sky130_fd_sc_hd__nor2_1
XFILLER_272_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15049_ _23917_/Q _23916_/Q _15049_/C vssd1 vssd1 vccd1 vccd1 _15159_/B sky130_fd_sc_hd__and3_1
XFILLER_253_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_287_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_44_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23538_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_296_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19857_ _16223_/X _23562_/Q _19865_/S vssd1 vssd1 vccd1 vccd1 _19858_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18808_ _18808_/A vssd1 vssd1 vccd1 vccd1 _18808_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19788_ _19788_/A vssd1 vssd1 vccd1 vccd1 _23531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_284_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18739_ _16873_/X _23095_/Q _18741_/S vssd1 vssd1 vccd1 vccd1 _18740_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21750_ _21779_/A _21779_/B vssd1 vssd1 vccd1 vccd1 _21801_/C sky130_fd_sc_hd__xor2_4
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20701_ _20732_/A vssd1 vssd1 vccd1 vccd1 _20701_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_196_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21681_ _21681_/A vssd1 vssd1 vccd1 vccd1 _21681_/X sky130_fd_sc_hd__buf_2
XFILLER_211_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23420_ _23420_/CLK _23420_/D vssd1 vssd1 vccd1 vccd1 _23420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_297_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20632_ _20632_/A vssd1 vssd1 vccd1 vccd1 _20632_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_338_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23351_ _23446_/CLK _23351_/D vssd1 vssd1 vccd1 vccd1 _23351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20563_ _20632_/A vssd1 vssd1 vccd1 vccd1 _20563_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_354_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_353_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22302_ _23566_/CLK _22302_/D vssd1 vssd1 vccd1 vccd1 _22302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_326_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23282_ _23538_/CLK _23282_/D vssd1 vssd1 vccd1 vccd1 _23282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_354_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20494_ _14546_/X _14195_/A _21336_/A _20493_/Y vssd1 vssd1 vccd1 vccd1 _21333_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_4_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22233_ _23812_/Q _21683_/X _22232_/Y _21660_/X vssd1 vssd1 vccd1 vccd1 _22234_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_117_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_307_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22164_ _23809_/Q _22130_/B _22163_/X _22129_/A vssd1 vssd1 vccd1 vccd1 _22164_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21115_ _21121_/A _21115_/B vssd1 vssd1 vccd1 vccd1 _23853_/D sky130_fd_sc_hd__nor2_1
XTAP_6938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22095_ _22116_/A _21984_/X _22094_/X _21896_/X vssd1 vssd1 vccd1 vccd1 _23936_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21046_ _20700_/A _21027_/X _21045_/X _21037_/X vssd1 vssd1 vccd1 vccd1 _23833_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_332_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22997_ _23009_/CLK _22997_/D vssd1 vssd1 vccd1 vccd1 _22997_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_234_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12750_ _22311_/Q _23447_/Q _12750_/S vssd1 vssd1 vccd1 vccd1 _12750_/X sky130_fd_sc_hd__mux2_1
XFILLER_243_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21948_ _23833_/Q _21947_/Y _22083_/A vssd1 vssd1 vccd1 vccd1 _21948_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11701_/A vssd1 vssd1 vccd1 vccd1 _11702_/A sky130_fd_sc_hd__buf_4
XFILLER_231_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12681_ _23224_/Q _23192_/Q _23160_/Q _23128_/Q _12680_/X _11166_/A vssd1 vssd1 vccd1
+ vccd1 _12682_/B sky130_fd_sc_hd__mux4_2
XFILLER_203_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21879_ _21879_/A _21879_/B vssd1 vssd1 vccd1 vccd1 _21879_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _22902_/Q _14394_/X _14164_/X _22595_/Q vssd1 vssd1 vccd1 vccd1 _14550_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23618_ _23624_/CLK _23618_/D vssd1 vssd1 vccd1 vccd1 _23618_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_187_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _12506_/A vssd1 vssd1 vccd1 vccd1 _12485_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14351_ _14349_/X _14350_/X _14351_/S vssd1 vssd1 vccd1 vccd1 _14354_/A sky130_fd_sc_hd__mux2_1
XFILLER_357_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23549_ _23549_/CLK _23549_/D vssd1 vssd1 vccd1 vccd1 _23549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_317_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11563_ _11701_/A vssd1 vssd1 vccd1 vccd1 _12458_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_357_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13302_ _13565_/A vssd1 vssd1 vccd1 vccd1 _13403_/B sky130_fd_sc_hd__clkbuf_2
X_17070_ _17070_/A vssd1 vssd1 vccd1 vccd1 _17070_/X sky130_fd_sc_hd__buf_2
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14282_ _13502_/A _13300_/B _14317_/S vssd1 vssd1 vccd1 vccd1 _14282_/X sky130_fd_sc_hd__mux2_1
XFILLER_356_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11494_ _11196_/A _11493_/X _13051_/A vssd1 vssd1 vccd1 vccd1 _11494_/X sky130_fd_sc_hd__a21o_1
XFILLER_171_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16021_ _23680_/Q _16021_/B vssd1 vssd1 vccd1 vccd1 _16021_/X sky130_fd_sc_hd__or2_1
X_13233_ _11278_/A _13223_/X _13232_/X _13184_/A vssd1 vssd1 vccd1 vccd1 _20353_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_7_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_313_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_313_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13164_ _21448_/B _13185_/S _11403_/A _13163_/Y vssd1 vssd1 vccd1 vccd1 _13187_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_312_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_313_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12115_ _12656_/A _12115_/B vssd1 vssd1 vccd1 vccd1 _12115_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17972_ _18052_/A vssd1 vssd1 vccd1 vccd1 _17972_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_312_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13095_ _13095_/A _13095_/B vssd1 vssd1 vccd1 vccd1 _13095_/Y sky130_fd_sc_hd__nor2_1
XFILLER_312_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19711_ _19711_/A vssd1 vssd1 vccd1 vccd1 _23497_/D sky130_fd_sc_hd__clkbuf_1
X_12046_ _23219_/Q _23187_/Q _23155_/Q _23123_/Q _12042_/S _12671_/A vssd1 vssd1 vccd1
+ vccd1 _12047_/B sky130_fd_sc_hd__mux4_1
X_16923_ _22613_/Q _16927_/A vssd1 vssd1 vccd1 vccd1 _17325_/B sky130_fd_sc_hd__or2_2
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_306_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19642_ _19642_/A vssd1 vssd1 vccd1 vccd1 _23466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16854_ _19204_/A vssd1 vssd1 vccd1 vccd1 _16854_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_226_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_322_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _23674_/Q _15905_/B vssd1 vssd1 vccd1 vccd1 _15805_/X sky130_fd_sc_hd__or2_1
XFILLER_322_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19573_ _23436_/Q _19188_/A _19577_/S vssd1 vssd1 vccd1 vccd1 _19574_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13997_ _14000_/A _14093_/A vssd1 vssd1 vccd1 vccd1 _13997_/Y sky130_fd_sc_hd__nor2_4
X_16785_ _22512_/Q _16783_/X _16784_/X input27/X vssd1 vssd1 vccd1 vccd1 _16786_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_292_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18524_ _23004_/Q _18530_/B vssd1 vssd1 vccd1 vccd1 _18524_/Y sky130_fd_sc_hd__nand2_1
XFILLER_283_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_2_0_wb_clk_i _23945_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_12948_ _22474_/Q _22634_/Q _22313_/Q _23449_/Q _12024_/X _12025_/X vssd1 vssd1 vccd1
+ vccd1 _12949_/B sky130_fd_sc_hd__mux4_1
X_15736_ _15724_/X _14588_/A _15726_/X _15735_/Y _15558_/A vssd1 vssd1 vccd1 vccd1
+ _15736_/X sky130_fd_sc_hd__a221o_1
XFILLER_206_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_162_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23877_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18455_ _22978_/Q _18465_/B vssd1 vssd1 vccd1 vccd1 _18455_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15667_ _18827_/A vssd1 vssd1 vccd1 vccd1 _19220_/A sky130_fd_sc_hd__clkbuf_2
X_12879_ _12886_/A _12878_/X _12700_/X vssd1 vssd1 vccd1 vccd1 _12879_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17406_ _22616_/Q _16214_/X _17410_/S vssd1 vssd1 vccd1 vccd1 _17407_/A sky130_fd_sc_hd__mux2_1
X_14618_ _18263_/B _14509_/X _14513_/X _22947_/Q vssd1 vssd1 vccd1 vccd1 _14618_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18386_ _22956_/Q _18386_/B vssd1 vssd1 vccd1 vccd1 _18392_/C sky130_fd_sc_hd__and2_4
X_15598_ _23733_/Q _23863_/Q _16103_/S vssd1 vssd1 vccd1 vccd1 _15598_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17337_ _17371_/A vssd1 vssd1 vccd1 vccd1 _17882_/S sky130_fd_sc_hd__clkbuf_2
X_14549_ _14548_/X _21320_/A _14557_/A vssd1 vssd1 vccd1 vccd1 _16457_/B sky130_fd_sc_hd__mux2_1
XFILLER_308_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_336_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_308_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_335_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17268_ _17268_/A vssd1 vssd1 vccd1 vccd1 _17268_/X sky130_fd_sc_hd__buf_2
XFILLER_135_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19007_ _19007_/A vssd1 vssd1 vccd1 vccd1 _23199_/D sky130_fd_sc_hd__clkbuf_1
X_16219_ _16219_/A vssd1 vssd1 vccd1 vccd1 _22296_/D sky130_fd_sc_hd__clkbuf_1
X_17199_ _17255_/A vssd1 vssd1 vccd1 vccd1 _17199_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_347_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_288_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19909_ _16300_/X _23586_/Q _19909_/S vssd1 vssd1 vccd1 vccd1 _19910_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_331_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22920_ _22956_/CLK _22920_/D vssd1 vssd1 vccd1 vccd1 _22920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_290_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22851_ _23426_/CLK _22851_/D vssd1 vssd1 vccd1 vccd1 _22851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21802_ _21548_/A _21548_/B _21690_/X _21803_/B vssd1 vssd1 vccd1 vccd1 _21804_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22782_ _23144_/CLK _22782_/D vssd1 vssd1 vccd1 vccd1 _22782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21733_ _21733_/A _21733_/B vssd1 vssd1 vccd1 vccd1 _21734_/B sky130_fd_sc_hd__nor2_1
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21664_ _21661_/X _21662_/Y _22234_/A vssd1 vssd1 vccd1 vccd1 _21664_/Y sky130_fd_sc_hd__a21oi_1
X_23403_ _23531_/CLK _23403_/D vssd1 vssd1 vccd1 vccd1 _23403_/Q sky130_fd_sc_hd__dfxtp_1
X_20615_ _20615_/A vssd1 vssd1 vccd1 vccd1 _20616_/A sky130_fd_sc_hd__inv_2
XFILLER_354_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_339_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21595_ _21515_/B _21593_/Y _21594_/Y _21327_/X vssd1 vssd1 vccd1 vccd1 _21595_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_138_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23334_ _23526_/CLK _23334_/D vssd1 vssd1 vccd1 vccd1 _23334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20546_ _20891_/A vssd1 vssd1 vccd1 vccd1 _20936_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_137_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23265_ _23553_/CLK _23265_/D vssd1 vssd1 vccd1 vccd1 _23265_/Q sky130_fd_sc_hd__dfxtp_1
X_20477_ _20723_/A _20467_/X _20476_/X _20472_/X vssd1 vssd1 vccd1 vccd1 _23709_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_180_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22216_ _22216_/A _22224_/A vssd1 vssd1 vccd1 vccd1 _22218_/A sky130_fd_sc_hd__and2_1
XFILLER_341_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23196_ _23545_/CLK _23196_/D vssd1 vssd1 vccd1 vccd1 _23196_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22147_ _22139_/A _21984_/X _22146_/X _22122_/X vssd1 vssd1 vccd1 vccd1 _23938_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput380 _14040_/X vssd1 vssd1 vccd1 vccd1 din0[15] sky130_fd_sc_hd__buf_2
XTAP_6746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput391 _14060_/X vssd1 vssd1 vccd1 vccd1 din0[25] sky130_fd_sc_hd__buf_2
XTAP_6757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22078_ _22057_/B _22059_/B _22057_/A vssd1 vssd1 vccd1 vccd1 _22082_/A sky130_fd_sc_hd__o21bai_1
XTAP_6779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13920_ _13920_/A _13920_/B vssd1 vssd1 vccd1 vccd1 _15078_/A sky130_fd_sc_hd__xnor2_4
X_21029_ _20654_/A _21027_/X _21028_/X _21023_/X vssd1 vssd1 vccd1 vccd1 _23826_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_281_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_274_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13851_ _13851_/A _13863_/B vssd1 vssd1 vccd1 vccd1 _13851_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12802_ _23929_/Q _13234_/S _12801_/X vssd1 vssd1 vccd1 vccd1 _13534_/B sky130_fd_sc_hd__o21ai_2
XFILLER_290_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16570_ _16592_/A vssd1 vssd1 vccd1 vccd1 _16579_/S sky130_fd_sc_hd__buf_6
XFILLER_216_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13782_ _12661_/B _13836_/B _13781_/X vssd1 vssd1 vccd1 vccd1 _13782_/X sky130_fd_sc_hd__a21o_1
XINSDIODE2_408 _14007_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_419 _14060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12733_ _12733_/A vssd1 vssd1 vccd1 vccd1 _12733_/X sky130_fd_sc_hd__buf_6
XFILLER_231_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15521_ _14210_/X _21766_/A _15520_/X vssd1 vssd1 vccd1 vccd1 _18817_/A sky130_fd_sc_hd__o21a_4
XFILLER_349_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18240_ _22908_/Q _18240_/B vssd1 vssd1 vccd1 vccd1 _18240_/X sky130_fd_sc_hd__or2_1
X_15452_ _15003_/A _15438_/X _15451_/X vssd1 vssd1 vccd1 vccd1 _17122_/A sky130_fd_sc_hd__o21ai_4
XFILLER_204_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12664_ _12664_/A _12636_/A vssd1 vssd1 vccd1 vccd1 _15582_/A sky130_fd_sc_hd__nor2b_2
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14403_ _15826_/A _16936_/B _20191_/A vssd1 vssd1 vccd1 vccd1 _14404_/B sky130_fd_sc_hd__mux2_1
XFILLER_129_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11615_ _12656_/A _11615_/B vssd1 vssd1 vccd1 vccd1 _11615_/X sky130_fd_sc_hd__or2_1
X_18171_ _22890_/Q _22891_/Q vssd1 vssd1 vccd1 vccd1 _18171_/X sky130_fd_sc_hd__and2b_1
X_15383_ _14968_/Y _15181_/A _15183_/A _15382_/Y vssd1 vssd1 vccd1 vccd1 _21235_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_168_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12595_ _23915_/Q vssd1 vssd1 vccd1 vccd1 _17033_/A sky130_fd_sc_hd__inv_6
XFILLER_204_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17122_ _17122_/A vssd1 vssd1 vccd1 vccd1 _17122_/Y sky130_fd_sc_hd__inv_2
X_14334_ _14952_/S vssd1 vssd1 vccd1 vccd1 _15132_/S sky130_fd_sc_hd__buf_2
X_11546_ _13064_/A _11545_/X _11288_/A vssd1 vssd1 vccd1 vccd1 _11546_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17053_ _23467_/Q _16987_/X _16988_/X _17042_/X _17052_/Y vssd1 vssd1 vccd1 vccd1
+ _17053_/X sky130_fd_sc_hd__a32o_1
XFILLER_143_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14265_ _14368_/A vssd1 vssd1 vccd1 vccd1 _14848_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_344_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11477_ _22387_/Q _22419_/Q _22708_/Q _23075_/Q _11461_/X _11462_/X vssd1 vssd1 vccd1
+ vccd1 _11477_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16004_ _16004_/A _16004_/B vssd1 vssd1 vccd1 vccd1 _16004_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13216_ _13216_/A _13216_/B vssd1 vssd1 vccd1 vccd1 _13216_/X sky130_fd_sc_hd__or2_1
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14196_ _14196_/A _14196_/B vssd1 vssd1 vccd1 vccd1 _14196_/Y sky130_fd_sc_hd__nand2_1
XFILLER_354_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13147_ _11169_/A _13144_/X _13146_/X vssd1 vssd1 vccd1 vccd1 _13147_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_286_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ _22829_/Q _17950_/X _17954_/X _17948_/X vssd1 vssd1 vccd1 vccd1 _22829_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _22140_/A _20374_/A _13296_/B vssd1 vssd1 vccd1 vccd1 _14276_/B sky130_fd_sc_hd__mux2_4
XFILLER_112_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12029_ _12029_/A vssd1 vssd1 vccd1 vccd1 _12029_/X sky130_fd_sc_hd__buf_6
X_16906_ _16905_/X _22549_/Q _16909_/S vssd1 vssd1 vccd1 vccd1 _16907_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17886_ _18142_/A _18172_/A vssd1 vssd1 vccd1 vccd1 _18191_/A sky130_fd_sc_hd__nor2_2
XFILLER_39_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19625_ _23460_/Q _19264_/A _19625_/S vssd1 vssd1 vccd1 vccd1 _19626_/A sky130_fd_sc_hd__mux2_1
X_16837_ _16837_/A vssd1 vssd1 vccd1 vccd1 _22527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19556_ _19612_/A vssd1 vssd1 vccd1 vccd1 _19625_/S sky130_fd_sc_hd__buf_6
XFILLER_280_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16768_ _16777_/A _16768_/B vssd1 vssd1 vccd1 vccd1 _16769_/A sky130_fd_sc_hd__or2_1
XFILLER_53_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18507_ _18520_/A vssd1 vssd1 vccd1 vccd1 _18507_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15719_ _13599_/X _16031_/S _15718_/Y _15636_/A vssd1 vssd1 vccd1 vccd1 _15723_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_280_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19487_ _19487_/A vssd1 vssd1 vccd1 vccd1 _23397_/D sky130_fd_sc_hd__clkbuf_1
X_16699_ _16699_/A vssd1 vssd1 vccd1 vccd1 _22488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18438_ _18441_/A _18438_/B vssd1 vssd1 vccd1 vccd1 _18438_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_349_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_355_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18369_ _22950_/Q _18369_/B vssd1 vssd1 vccd1 vccd1 _18375_/C sky130_fd_sc_hd__and2_1
XFILLER_348_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20400_ _20400_/A _20400_/B vssd1 vssd1 vccd1 vccd1 _20400_/Y sky130_fd_sc_hd__nor2_1
XFILLER_193_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21380_ _21560_/A vssd1 vssd1 vccd1 vccd1 _22130_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_309_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20331_ _23673_/Q _20338_/B vssd1 vssd1 vccd1 vccd1 _20331_/X sky130_fd_sc_hd__or2_1
XFILLER_135_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_289_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23050_ _23500_/CLK _23050_/D vssd1 vssd1 vccd1 vccd1 _23050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_351_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20262_ _20262_/A vssd1 vssd1 vccd1 vccd1 _20387_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_350_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22001_ _21978_/A _21977_/B _21977_/A vssd1 vssd1 vccd1 vccd1 _22002_/B sky130_fd_sc_hd__a21bo_1
XTAP_6009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_289_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20193_ _20187_/X _20189_/X _20190_/Y _21406_/A _20192_/X vssd1 vssd1 vccd1 vccd1
+ _20579_/A sky130_fd_sc_hd__a32o_4
XFILLER_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput108 dout1[10] vssd1 vssd1 vccd1 vccd1 input108/X sky130_fd_sc_hd__clkbuf_1
XFILLER_248_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput119 dout1[20] vssd1 vssd1 vccd1 vccd1 input119/X sky130_fd_sc_hd__clkbuf_1
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22903_ _22908_/CLK _22903_/D vssd1 vssd1 vccd1 vccd1 _22903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23883_ _23926_/CLK _23883_/D vssd1 vssd1 vccd1 vccd1 _23883_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_99_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22834_ _23632_/CLK _22834_/D vssd1 vssd1 vccd1 vccd1 _22834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22765_ _23068_/CLK _22765_/D vssd1 vssd1 vccd1 vccd1 _22765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21716_ _21716_/A _21716_/B vssd1 vssd1 vccd1 vccd1 _21716_/X sky130_fd_sc_hd__or2_1
XFILLER_80_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22696_ _23446_/CLK _22696_/D vssd1 vssd1 vccd1 vccd1 _22696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_358_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_346_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_327_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21647_ _21077_/D _21646_/X _21865_/A vssd1 vssd1 vccd1 vccd1 _21653_/A sky130_fd_sc_hd__mux2_1
XFILLER_355_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11400_ _11400_/A vssd1 vssd1 vccd1 vccd1 _11401_/A sky130_fd_sc_hd__buf_2
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12380_ _11330_/A _12379_/X _11679_/A vssd1 vssd1 vccd1 vccd1 _12380_/X sky130_fd_sc_hd__o21a_1
XFILLER_166_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21578_ _21569_/X _21574_/Y _21576_/Y _21577_/X vssd1 vssd1 vccd1 vccd1 _21579_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_166_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_338_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23317_ _23541_/CLK _23317_/D vssd1 vssd1 vccd1 vccd1 _23317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11331_ _11863_/A vssd1 vssd1 vccd1 vccd1 _12105_/A sky130_fd_sc_hd__buf_4
X_20529_ _21191_/A _13479_/X _15180_/A _20528_/X vssd1 vssd1 vccd1 vccd1 _20781_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_315_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14050_ _14049_/X _13817_/B _14041_/X input228/X vssd1 vssd1 vccd1 vccd1 _14050_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_153_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23248_ _23537_/CLK _23248_/D vssd1 vssd1 vccd1 vccd1 _23248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11262_ _23892_/Q _23891_/Q vssd1 vssd1 vccd1 vccd1 _13412_/A sky130_fd_sc_hd__or2b_1
XTAP_7211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13001_ _23227_/Q _23195_/Q _23163_/Q _23131_/Q _12733_/X _12734_/X vssd1 vssd1 vccd1
+ vccd1 _13002_/B sky130_fd_sc_hd__mux4_2
XTAP_7233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11193_ _12071_/A vssd1 vssd1 vccd1 vccd1 _11584_/A sky130_fd_sc_hd__clkbuf_4
X_23179_ _23531_/CLK _23179_/D vssd1 vssd1 vccd1 vccd1 _23179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17740_ _17740_/A vssd1 vssd1 vccd1 vccd1 _22747_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14952_ _14333_/A _14303_/X _14952_/S vssd1 vssd1 vccd1 vccd1 _14953_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13903_ _13903_/A _13903_/B vssd1 vssd1 vccd1 vccd1 _14865_/A sky130_fd_sc_hd__xor2_4
XFILLER_48_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17671_ _22717_/Q _17559_/X _17671_/S vssd1 vssd1 vccd1 vccd1 _17672_/A sky130_fd_sc_hd__mux2_1
X_14883_ _14822_/X _14834_/X _14880_/X _14882_/X vssd1 vssd1 vccd1 vccd1 _14883_/X
+ sky130_fd_sc_hd__a22o_1
X_19410_ _19410_/A vssd1 vssd1 vccd1 vccd1 _23364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16622_ _16622_/A vssd1 vssd1 vccd1 vccd1 _22459_/D sky130_fd_sc_hd__clkbuf_1
X_13834_ _13834_/A vssd1 vssd1 vccd1 vccd1 _13875_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_262_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_205 _14228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_216 _14619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_227 _17052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19341_ _19409_/S vssd1 vssd1 vccd1 vccd1 _19350_/S sky130_fd_sc_hd__buf_6
XFILLER_188_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13765_ _13765_/A _13765_/B _13765_/C _13777_/B vssd1 vssd1 vccd1 vccd1 _13864_/A
+ sky130_fd_sc_hd__or4_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16553_ _15168_/X _22429_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _16554_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_238 _15204_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_249 _21720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15504_ _19976_/B _15589_/A _15590_/A _23635_/Q vssd1 vssd1 vccd1 vccd1 _15504_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12716_ _12716_/A vssd1 vssd1 vccd1 vccd1 _12716_/X sky130_fd_sc_hd__buf_6
XFILLER_149_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19272_ _19169_/X _23302_/Q _19278_/S vssd1 vssd1 vccd1 vccd1 _19273_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16484_ _16484_/A vssd1 vssd1 vccd1 vccd1 _22399_/D sky130_fd_sc_hd__clkbuf_1
X_13696_ _13715_/A _13985_/B _14006_/C vssd1 vssd1 vccd1 vccd1 _13697_/A sky130_fd_sc_hd__and3_4
XFILLER_94_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18223_ _22901_/Q _18227_/B vssd1 vssd1 vccd1 vccd1 _18223_/X sky130_fd_sc_hd__or2_1
XPHY_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12647_ _22373_/Q _22405_/Q _22694_/Q _23061_/Q _12680_/A _11973_/X vssd1 vssd1 vccd1
+ vccd1 _12647_/X sky130_fd_sc_hd__mux4_2
X_15435_ _15031_/Y _15181_/A _15183_/A _15434_/Y vssd1 vssd1 vccd1 vccd1 _21238_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_87_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_318_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18154_ _18154_/A vssd1 vssd1 vccd1 vccd1 _22887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15366_ _14570_/X _21233_/A _15364_/Y _15365_/X vssd1 vssd1 vccd1 vccd1 _15367_/B
+ sky130_fd_sc_hd__o22a_1
X_12578_ _23465_/Q _23561_/Q _22525_/Q _22329_/Q _12324_/X _12325_/X vssd1 vssd1 vccd1
+ vccd1 _12578_/X sky130_fd_sc_hd__mux4_1
XFILLER_318_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17105_ _14535_/X _17104_/X _17116_/S vssd1 vssd1 vccd1 vccd1 _17105_/X sky130_fd_sc_hd__mux2_1
X_11529_ _13073_/A _11529_/B vssd1 vssd1 vccd1 vccd1 _11529_/X sky130_fd_sc_hd__or2_1
X_14317_ _14307_/B _13525_/B _14317_/S vssd1 vssd1 vccd1 vccd1 _14651_/B sky130_fd_sc_hd__mux2_1
X_18085_ _22865_/Q _18082_/X _18083_/X _22998_/Q _18084_/X vssd1 vssd1 vccd1 vccd1
+ _18085_/X sky130_fd_sc_hd__a221o_1
XFILLER_318_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15297_ _13528_/B _15082_/X _15296_/X vssd1 vssd1 vccd1 vccd1 _15297_/X sky130_fd_sc_hd__o21a_1
XFILLER_345_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_305_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17036_ _17000_/X _17029_/X _17035_/X _17012_/X vssd1 vssd1 vccd1 vccd1 _17036_/X
+ sky130_fd_sc_hd__o211a_2
X_14248_ _22487_/Q _13692_/A _14245_/X _14247_/X _14072_/A vssd1 vssd1 vccd1 vccd1
+ _14248_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_172_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14179_ _14179_/A vssd1 vssd1 vccd1 vccd1 _16118_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_301_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_298_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_313_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_286_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18987_ _18987_/A vssd1 vssd1 vccd1 vccd1 _23190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17938_ _17956_/A vssd1 vssd1 vccd1 vccd1 _17938_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_239_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17869_ _17869_/A vssd1 vssd1 vccd1 vccd1 _22805_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19608_ _23452_/Q _19239_/A _19610_/S vssd1 vssd1 vccd1 vccd1 _19609_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20880_ _20880_/A vssd1 vssd1 vccd1 vccd1 _23777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19539_ _19539_/A vssd1 vssd1 vccd1 vccd1 _23421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22550_ _23489_/CLK _22550_/D vssd1 vssd1 vccd1 vccd1 _22550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_329_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21501_ _21513_/A _21501_/B vssd1 vssd1 vccd1 vccd1 _21503_/A sky130_fd_sc_hd__and2b_1
XFILLER_166_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_355_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22481_ _23456_/CLK _22481_/D vssd1 vssd1 vccd1 vccd1 _22481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21432_ _23915_/Q _21437_/A vssd1 vssd1 vccd1 vccd1 _21432_/Y sky130_fd_sc_hd__nand2_1
XFILLER_348_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_296_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21363_ _21327_/X _21355_/X _21361_/X _22093_/A vssd1 vssd1 vccd1 vccd1 _21363_/X
+ sky130_fd_sc_hd__o211a_1
X_23102_ _23582_/CLK _23102_/D vssd1 vssd1 vccd1 vccd1 _23102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20314_ _21888_/B vssd1 vssd1 vccd1 vccd1 _20314_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput90 dout0[52] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21294_ _21294_/A _21294_/B _21294_/C vssd1 vssd1 vccd1 vccd1 _21295_/B sky130_fd_sc_hd__nor3_1
XFILLER_116_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23033_ _23419_/CLK _23033_/D vssd1 vssd1 vccd1 vccd1 _23033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_289_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20245_ _23662_/Q _20277_/B vssd1 vssd1 vccd1 vccd1 _20245_/X sky130_fd_sc_hd__or2_1
XFILLER_332_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_331_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_320_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20176_ _16940_/X _17653_/A _20172_/Y _20175_/X vssd1 vssd1 vccd1 vccd1 _20996_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_254_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_320_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23935_ _23935_/CLK _23935_/D vssd1 vssd1 vccd1 vccd1 _23935_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_340_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23866_ _23866_/CLK _23866_/D vssd1 vssd1 vccd1 vccd1 _23866_/Q sky130_fd_sc_hd__dfxtp_1
X_11880_ _11863_/A _11876_/X _11879_/X _11680_/A vssd1 vssd1 vccd1 vccd1 _11880_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22817_ _22822_/CLK _22817_/D vssd1 vssd1 vccd1 vccd1 _22817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23797_ _23810_/CLK _23797_/D vssd1 vssd1 vccd1 vccd1 _23797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13550_ _13647_/A _23940_/Q _13490_/X _13549_/Y vssd1 vssd1 vccd1 vccd1 _13686_/A
+ sky130_fd_sc_hd__o211a_1
X_22748_ _23048_/CLK _22748_/D vssd1 vssd1 vccd1 vccd1 _22748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_337_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12501_ _23894_/Q vssd1 vssd1 vccd1 vccd1 _12501_/X sky130_fd_sc_hd__clkbuf_4
X_13481_ _13879_/B _13481_/B vssd1 vssd1 vccd1 vccd1 _20530_/B sky130_fd_sc_hd__nand2_4
X_22679_ _23496_/CLK _22679_/D vssd1 vssd1 vccd1 vccd1 _22679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15220_ _23789_/Q _15219_/X _14919_/X vssd1 vssd1 vccd1 vccd1 _15220_/X sky130_fd_sc_hd__a21o_1
X_12432_ _23399_/Q _23015_/Q _23367_/Q _23335_/Q _12424_/S _12538_/A vssd1 vssd1 vccd1
+ vccd1 _12432_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_343_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15151_ _14936_/A _15141_/X _15147_/Y _15150_/X vssd1 vssd1 vccd1 vccd1 _15151_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12363_ _12196_/A _12362_/X _11229_/A vssd1 vssd1 vccd1 vccd1 _12363_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14102_ _18178_/B vssd1 vssd1 vccd1 vccd1 _18187_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_295_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11314_ _12476_/A vssd1 vssd1 vccd1 vccd1 _11815_/A sky130_fd_sc_hd__clkbuf_4
X_15082_ _15583_/A vssd1 vssd1 vccd1 vccd1 _15082_/X sky130_fd_sc_hd__buf_4
XFILLER_299_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12294_ _12567_/A _12293_/X _11229_/A vssd1 vssd1 vccd1 vccd1 _12294_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_342_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18910_ _23156_/Q _18820_/X _18918_/S vssd1 vssd1 vccd1 vccd1 _18911_/A sky130_fd_sc_hd__mux2_1
XFILLER_342_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14033_ input218/X _14027_/X _14032_/X vssd1 vssd1 vccd1 vccd1 _14033_/X sky130_fd_sc_hd__a21bo_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11245_ _11559_/A vssd1 vssd1 vccd1 vccd1 _11246_/A sky130_fd_sc_hd__buf_2
XFILLER_106_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19890_ _16271_/X _23577_/Q _19898_/S vssd1 vssd1 vccd1 vccd1 _19891_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18841_ _23130_/Q _18840_/X _18850_/S vssd1 vssd1 vccd1 vccd1 _18842_/A sky130_fd_sc_hd__mux2_1
XTAP_7074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ _12307_/A vssd1 vssd1 vccd1 vccd1 _12082_/A sky130_fd_sc_hd__buf_6
XTAP_6351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_310_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18772_ _18853_/A vssd1 vssd1 vccd1 vccd1 _18872_/S sky130_fd_sc_hd__buf_6
XTAP_6395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15984_ _20016_/B _15589_/X _15590_/X _23647_/Q vssd1 vssd1 vccd1 vccd1 _15984_/X
+ sky130_fd_sc_hd__o22a_2
XTAP_5650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17723_ _17723_/A vssd1 vssd1 vccd1 vccd1 _22740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_314_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14935_ _18275_/A _14932_/X _14934_/X _22950_/Q vssd1 vssd1 vccd1 vccd1 _14935_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17654_ _21301_/B _17653_/B _17653_/Y _17390_/X vssd1 vssd1 vccd1 vccd1 _22711_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14866_ _14866_/A vssd1 vssd1 vccd1 vccd1 _15010_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_291_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_330_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16605_ _16197_/X _22453_/Q _16605_/S vssd1 vssd1 vccd1 vccd1 _16606_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13817_ _13855_/A _13817_/B vssd1 vssd1 vccd1 vccd1 _13818_/A sky130_fd_sc_hd__and2_1
X_17585_ _18811_/A vssd1 vssd1 vccd1 vccd1 _17585_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14797_ _14839_/A _14790_/X _14796_/X vssd1 vssd1 vccd1 vccd1 _14797_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_330_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19324_ _19324_/A vssd1 vssd1 vccd1 vccd1 _19333_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_69_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23480_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_251_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16536_ _16592_/A vssd1 vssd1 vccd1 vccd1 _16605_/S sky130_fd_sc_hd__buf_6
XFILLER_259_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13748_ _13974_/B _13748_/B vssd1 vssd1 vccd1 vccd1 _13748_/Y sky130_fd_sc_hd__nor2_2
XFILLER_189_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19255_ _19255_/A vssd1 vssd1 vccd1 vccd1 _19255_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16467_ _14893_/X _22392_/Q _16469_/S vssd1 vssd1 vccd1 vccd1 _16468_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13679_ _17029_/S _13679_/B vssd1 vssd1 vccd1 vccd1 _13679_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18206_ _18245_/A vssd1 vssd1 vccd1 vccd1 _18206_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_319_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15418_ _22990_/Q _15620_/A _15621_/A input218/X vssd1 vssd1 vccd1 vccd1 _21708_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19186_ _19185_/X _23275_/Q _19195_/S vssd1 vssd1 vccd1 vccd1 _19187_/A sky130_fd_sc_hd__mux2_1
X_16398_ _16455_/S vssd1 vssd1 vccd1 vccd1 _16407_/S sky130_fd_sc_hd__buf_6
XFILLER_191_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18137_ _18138_/A _22884_/Q _18135_/X _18136_/Y vssd1 vssd1 vccd1 vccd1 _22883_/D
+ sky130_fd_sc_hd__o211a_1
X_15349_ _22925_/Q _14932_/X _14934_/X _15351_/A vssd1 vssd1 vccd1 vccd1 _15349_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_333_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18068_ _18098_/A vssd1 vssd1 vccd1 vccd1 _18068_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_176_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17019_ _14196_/A _17018_/X _17317_/S vssd1 vssd1 vccd1 vccd1 _17019_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20030_ _23621_/Q _20042_/C _20029_/Y vssd1 vssd1 vccd1 vccd1 _23621_/D sky130_fd_sc_hd__o21a_1
XFILLER_302_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_302_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21981_ _21981_/A _21981_/B vssd1 vssd1 vccd1 vccd1 _21981_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23720_ _23851_/CLK _23720_/D vssd1 vssd1 vccd1 vccd1 _23720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20932_ _23793_/Q _20925_/X _20931_/X _20920_/X vssd1 vssd1 vccd1 vccd1 _23793_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_215_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23651_ _23651_/CLK _23651_/D vssd1 vssd1 vccd1 vccd1 _23651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20863_ _20881_/A vssd1 vssd1 vccd1 vccd1 _20879_/A sky130_fd_sc_hd__clkbuf_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22602_ _23649_/CLK _22602_/D vssd1 vssd1 vccd1 vccd1 _22602_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_23_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23582_ _23582_/CLK _23582_/D vssd1 vssd1 vccd1 vccd1 _23582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20794_ _20806_/A _20794_/B vssd1 vssd1 vccd1 vccd1 _20795_/A sky130_fd_sc_hd__and2_1
XFILLER_329_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22533_ _23504_/CLK _22533_/D vssd1 vssd1 vccd1 vccd1 _22533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_356_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_328_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22464_ _23567_/CLK _22464_/D vssd1 vssd1 vccd1 vccd1 _22464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_356_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_337_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21415_ _23817_/Q _23751_/Q vssd1 vssd1 vccd1 vccd1 _21415_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22395_ _23563_/CLK _22395_/D vssd1 vssd1 vccd1 vccd1 _22395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_309_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_309_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_324_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21346_ _21346_/A vssd1 vssd1 vccd1 vccd1 _21346_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_163_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_351_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_340_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21277_ _21605_/A _21199_/B _21276_/Y _21270_/X vssd1 vssd1 vccd1 vccd1 _23907_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_351_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23016_ _23526_/CLK _23016_/D vssd1 vssd1 vccd1 vccd1 _23016_/Q sky130_fd_sc_hd__dfxtp_1
X_20228_ _21517_/A _20279_/B vssd1 vssd1 vccd1 vccd1 _20228_/Y sky130_fd_sc_hd__nand2_1
XFILLER_231_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_292_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20159_ _21285_/A _14133_/X _20139_/Y _20140_/X vssd1 vssd1 vccd1 vccd1 _21084_/B
+ sky130_fd_sc_hd__o31a_4
XFILLER_77_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _13084_/A _12976_/X _12980_/X _11133_/A vssd1 vssd1 vccd1 vccd1 _12981_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14720_ _22497_/Q _13691_/A _14238_/X _14719_/X _14242_/X vssd1 vssd1 vccd1 vccd1
+ _14720_/Y sky130_fd_sc_hd__o221ai_4
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23918_ _23918_/CLK _23918_/D vssd1 vssd1 vccd1 vccd1 _23918_/Q sky130_fd_sc_hd__dfxtp_4
X_11932_ _11914_/A _11929_/X _11931_/X _11348_/A vssd1 vssd1 vccd1 vccd1 _11932_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_273_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ _14651_/A _14651_/B vssd1 vssd1 vccd1 vccd1 _14651_/Y sky130_fd_sc_hd__nor2_1
X_11863_ _11863_/A _11863_/B vssd1 vssd1 vccd1 vccd1 _11863_/Y sky130_fd_sc_hd__nor2_1
X_23849_ _23851_/CLK _23849_/D vssd1 vssd1 vccd1 vccd1 _23849_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _23933_/Q _13884_/A _13601_/Y _14198_/B vssd1 vssd1 vccd1 vccd1 _13975_/A
+ sky130_fd_sc_hd__a22o_4
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _17370_/A vssd1 vssd1 vccd1 vccd1 _22605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_300_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ _22504_/Q _13691_/A _13888_/B _14581_/X vssd1 vssd1 vccd1 vccd1 _15244_/A
+ sky130_fd_sc_hd__o211ai_2
X_11794_ _14175_/A _12087_/A _11884_/B vssd1 vssd1 vccd1 vccd1 _11794_/X sky130_fd_sc_hd__a21o_1
XFILLER_158_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_300_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16321_ _16321_/A vssd1 vssd1 vccd1 vccd1 _22328_/D sky130_fd_sc_hd__clkbuf_1
X_13533_ _13619_/A _13531_/X _13532_/X _12005_/Y vssd1 vssd1 vccd1 vccd1 _13632_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_347_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19040_ _16844_/X _23214_/Q _19040_/S vssd1 vssd1 vccd1 vccd1 _19041_/A sky130_fd_sc_hd__mux2_1
X_16252_ _18817_/A vssd1 vssd1 vccd1 vccd1 _16252_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13464_ _14687_/A _13464_/B vssd1 vssd1 vccd1 vccd1 _13476_/A sky130_fd_sc_hd__xor2_4
XFILLER_335_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12415_ _23913_/Q _21340_/A _12415_/S vssd1 vssd1 vccd1 vccd1 _14791_/A sky130_fd_sc_hd__mux2_4
X_15203_ _13372_/Y _15580_/B _15202_/Y vssd1 vssd1 vccd1 vccd1 _15203_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_316_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13395_ _15718_/A _13395_/B _13395_/C _13395_/D vssd1 vssd1 vccd1 vccd1 _13400_/B
+ sky130_fd_sc_hd__or4_1
X_16183_ _11394_/A _14259_/A _16182_/X _14287_/Y _14836_/A vssd1 vssd1 vccd1 vccd1
+ _16183_/X sky130_fd_sc_hd__a221o_1
XFILLER_315_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15134_ _14854_/S _14845_/X _15249_/S vssd1 vssd1 vccd1 vccd1 _15134_/X sky130_fd_sc_hd__a21o_1
X_12346_ _14176_/A _13775_/B _20148_/A _13775_/D vssd1 vssd1 vccd1 vccd1 _13763_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_299_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_187_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23910_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_303_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_315_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19942_ _23596_/Q _19935_/C _19941_/Y vssd1 vssd1 vccd1 vccd1 _23596_/D sky130_fd_sc_hd__o21a_1
X_15065_ _23595_/Q _14450_/A _14455_/A _23627_/Q vssd1 vssd1 vccd1 vccd1 _15065_/X
+ sky130_fd_sc_hd__o22a_4
Xclkbuf_leaf_116_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23599_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_302_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12277_ _22783_/Q _22751_/Q _22652_/Q _22719_/Q _11305_/A _11869_/X vssd1 vssd1 vccd1
+ vccd1 _12278_/B sky130_fd_sc_hd__mux4_1
XFILLER_141_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14016_ input240/X _14004_/X _14015_/X vssd1 vssd1 vccd1 vccd1 _14016_/X sky130_fd_sc_hd__a21o_4
XFILLER_330_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11228_ _11705_/A vssd1 vssd1 vccd1 vccd1 _11229_/A sky130_fd_sc_hd__buf_4
X_19873_ _19873_/A vssd1 vssd1 vccd1 vccd1 _23569_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18824_ _18824_/A vssd1 vssd1 vccd1 vccd1 _18824_/X sky130_fd_sc_hd__buf_2
XFILLER_96_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_295_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11159_ _11189_/A vssd1 vssd1 vccd1 vccd1 _12538_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_283_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18755_ _16895_/X _23102_/Q _18763_/S vssd1 vssd1 vccd1 vccd1 _18756_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15967_ _15923_/A _15941_/X _15966_/X _15162_/A vssd1 vssd1 vccd1 vccd1 _15967_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput280 versionID[0] vssd1 vssd1 vccd1 vccd1 input280/X sky130_fd_sc_hd__clkbuf_2
XFILLER_341_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17706_ _17717_/A vssd1 vssd1 vccd1 vccd1 _17715_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_76_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14918_ _14918_/A vssd1 vssd1 vccd1 vccd1 _14919_/A sky130_fd_sc_hd__clkbuf_2
X_18686_ _18686_/A vssd1 vssd1 vccd1 vccd1 _23071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15898_ _19239_/A vssd1 vssd1 vccd1 vccd1 _15898_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17637_ _22706_/Q _17636_/X _17640_/S vssd1 vssd1 vccd1 vccd1 _17638_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14849_ _15538_/A _14847_/X _15011_/A vssd1 vssd1 vccd1 vccd1 _14849_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_251_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17568_ _17568_/A vssd1 vssd1 vccd1 vccd1 _22684_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19307_ _19220_/X _23318_/Q _19311_/S vssd1 vssd1 vccd1 vccd1 _19308_/A sky130_fd_sc_hd__mux2_1
X_16519_ _16519_/A vssd1 vssd1 vccd1 vccd1 _22415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_338_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17499_ _22657_/Q _16243_/X _17505_/S vssd1 vssd1 vccd1 vccd1 _17500_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19238_ _19238_/A vssd1 vssd1 vccd1 vccd1 _23291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_286_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19169_ _19169_/A vssd1 vssd1 vccd1 vccd1 _19169_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_293_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_306_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21200_ _11069_/D _21196_/X _21199_/Y _21186_/X vssd1 vssd1 vccd1 vccd1 _23879_/D
+ sky130_fd_sc_hd__o211a_1
X_22180_ _22205_/A _22181_/B vssd1 vssd1 vccd1 vccd1 _22182_/A sky130_fd_sc_hd__nand2_1
XFILLER_118_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_306_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21131_ _23860_/Q _21123_/X _21124_/X _20655_/A vssd1 vssd1 vccd1 vccd1 _21132_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_172_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21062_ _23839_/Q _20996_/B _21060_/Y _21061_/X vssd1 vssd1 vccd1 vccd1 _23839_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20013_ _20016_/B _20021_/C _23616_/Q vssd1 vssd1 vccd1 vccd1 _20015_/B sky130_fd_sc_hd__a21oi_1
XFILLER_302_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21964_ _22038_/A _21940_/B _21932_/A vssd1 vssd1 vccd1 vccd1 _21965_/B sky130_fd_sc_hd__a21oi_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20915_ _13923_/B _20908_/X _20608_/B _20912_/X vssd1 vssd1 vccd1 vccd1 _20915_/X
+ sky130_fd_sc_hd__a211o_1
X_23703_ _23704_/CLK _23703_/D vssd1 vssd1 vccd1 vccd1 _23703_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21895_ _21081_/A _21880_/X _21886_/X _22215_/A _21894_/Y vssd1 vssd1 vccd1 vccd1
+ _21895_/X sky130_fd_sc_hd__a221o_1
XFILLER_14_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23634_ _23634_/CLK _23634_/D vssd1 vssd1 vccd1 vccd1 _23634_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_54_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20846_ _20864_/A vssd1 vssd1 vccd1 vccd1 _20846_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23565_ _23565_/CLK _23565_/D vssd1 vssd1 vccd1 vccd1 _23565_/Q sky130_fd_sc_hd__dfxtp_1
X_20777_ _20533_/Y _20773_/Y _20888_/C _20558_/A vssd1 vssd1 vccd1 vccd1 _20777_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_80_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_356_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22516_ _23700_/CLK _22516_/D vssd1 vssd1 vccd1 vccd1 _22516_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23496_ _23496_/CLK _23496_/D vssd1 vssd1 vccd1 vccd1 _23496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_357_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22447_ _23582_/CLK _22447_/D vssd1 vssd1 vccd1 vccd1 _22447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_309_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_346_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12200_ _22268_/Q _23084_/Q _23500_/Q _22429_/Q _11113_/A _12199_/X vssd1 vssd1 vccd1
+ vccd1 _12201_/B sky130_fd_sc_hd__mux4_2
XFILLER_325_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13180_ _13180_/A _13180_/B vssd1 vssd1 vccd1 vccd1 _13180_/X sky130_fd_sc_hd__or2_1
XFILLER_352_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_313_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22378_ _23449_/CLK _22378_/D vssd1 vssd1 vccd1 vccd1 _22378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12131_ _23473_/Q _23569_/Q _22533_/Q _22337_/Q _11151_/A _11613_/X vssd1 vssd1 vccd1
+ vccd1 _12131_/X sky130_fd_sc_hd__mux4_1
XFILLER_325_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21329_ _21922_/A vssd1 vssd1 vccd1 vccd1 _21329_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12062_ _13436_/A _12801_/A _11401_/A _12061_/Y vssd1 vssd1 vccd1 vccd1 _12168_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_145_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_321_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16870_ _19220_/A vssd1 vssd1 vccd1 vccd1 _16870_/X sky130_fd_sc_hd__buf_2
XFILLER_277_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ _14703_/X _21979_/A _15820_/X vssd1 vssd1 vccd1 vccd1 _18840_/A sky130_fd_sc_hd__a21o_4
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18540_ _18549_/A _18538_/Y _18539_/X _18203_/C vssd1 vssd1 vccd1 vccd1 _18550_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_292_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _16079_/A vssd1 vssd1 vccd1 vccd1 _15752_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_70 _13440_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _13022_/A _12964_/B vssd1 vssd1 vccd1 vccd1 _12965_/A sky130_fd_sc_hd__nor2_1
XFILLER_79_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_81 _21771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_92 _21846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14703_ _15746_/A vssd1 vssd1 vccd1 vccd1 _14703_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18471_ _22984_/Q _18478_/B vssd1 vssd1 vccd1 vccd1 _18471_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11915_ _23213_/Q _23181_/Q _23149_/Q _23117_/Q _11799_/X _11800_/X vssd1 vssd1 vccd1
+ vccd1 _11916_/B sky130_fd_sc_hd__mux4_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _15680_/Y _15682_/X _14896_/A vssd1 vssd1 vccd1 vccd1 _15683_/X sky130_fd_sc_hd__o21a_2
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _12904_/A _12895_/B vssd1 vssd1 vccd1 vccd1 _12895_/X sky130_fd_sc_hd__or2_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17422_ _17422_/A vssd1 vssd1 vccd1 vccd1 _22623_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_261_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14634_ _14301_/X _14304_/X _14651_/A vssd1 vssd1 vccd1 vccd1 _14634_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _12241_/A _11837_/Y _11839_/Y _11845_/Y vssd1 vssd1 vccd1 vccd1 _11846_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _17353_/A vssd1 vssd1 vccd1 vccd1 _22597_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _22303_/Q _23439_/Q _11777_/S vssd1 vssd1 vccd1 vccd1 _11778_/B sky130_fd_sc_hd__mux2_1
X_14565_ _15631_/A vssd1 vssd1 vccd1 vccd1 _14568_/A sky130_fd_sc_hd__buf_2
XFILLER_186_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16304_ _22323_/Q _16303_/X _16307_/S vssd1 vssd1 vccd1 vccd1 _16305_/A sky130_fd_sc_hd__mux2_1
XFILLER_348_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13516_ _12287_/B _13516_/B vssd1 vssd1 vccd1 vccd1 _13516_/X sky130_fd_sc_hd__and2b_1
X_17284_ _17245_/X _17282_/X _17262_/X _17283_/X vssd1 vssd1 vccd1 vccd1 _17284_/X
+ sky130_fd_sc_hd__a211o_1
X_14496_ _15148_/A _15148_/B vssd1 vssd1 vccd1 vccd1 _14497_/A sky130_fd_sc_hd__and2_2
XFILLER_335_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19023_ _16819_/X _23206_/Q _19029_/S vssd1 vssd1 vccd1 vccd1 _19024_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16235_ _16235_/A vssd1 vssd1 vccd1 vccd1 _22301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13447_ _14178_/A _14179_/A _23907_/Q _16016_/A vssd1 vssd1 vccd1 vccd1 _13448_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_328_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_304_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16166_ _14833_/A _15533_/Y _15942_/A vssd1 vssd1 vccd1 vccd1 _21283_/A sky130_fd_sc_hd__a21oi_4
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13378_ _13625_/A _13378_/B vssd1 vssd1 vccd1 vccd1 _13379_/C sky130_fd_sc_hd__xnor2_2
XFILLER_316_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_315_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_331_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15117_ input157/X _13652_/A _15110_/S input122/X vssd1 vssd1 vccd1 vccd1 _15117_/X
+ sky130_fd_sc_hd__a22o_4
X_12329_ _12329_/A vssd1 vssd1 vccd1 vccd1 _12329_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_336_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16097_ _16097_/A _16097_/B vssd1 vssd1 vccd1 vccd1 _16097_/X sky130_fd_sc_hd__or2_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_303_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19925_ _23592_/Q _19927_/C _18012_/X vssd1 vssd1 vccd1 vccd1 _19926_/B sky130_fd_sc_hd__o21ai_1
XFILLER_287_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15048_ _15048_/A vssd1 vssd1 vccd1 vccd1 _15048_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_142_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19856_ _19913_/S vssd1 vssd1 vccd1 vccd1 _19865_/S sky130_fd_sc_hd__buf_4
XFILLER_68_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_295_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18807_ _18807_/A vssd1 vssd1 vccd1 vccd1 _23119_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_352_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19787_ _23531_/Q _19185_/A _19793_/S vssd1 vssd1 vccd1 vccd1 _19788_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16999_ _22554_/Q _16922_/X _16973_/X _16998_/X vssd1 vssd1 vccd1 vccd1 _22554_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_37_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_84_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23576_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18738_ _18738_/A vssd1 vssd1 vccd1 vccd1 _23094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_284_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_13_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23407_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18669_ _23064_/Q _17607_/X _18669_/S vssd1 vssd1 vccd1 vccd1 _18670_/A sky130_fd_sc_hd__mux2_1
XFILLER_252_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20700_ _20700_/A _20731_/B vssd1 vssd1 vccd1 vccd1 _20705_/B sky130_fd_sc_hd__and2_2
XFILLER_252_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21680_ _21491_/X _21670_/X _21679_/Y vssd1 vssd1 vccd1 vccd1 _21680_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20631_ _20631_/A _20631_/B vssd1 vssd1 vccd1 vccd1 _20635_/B sky130_fd_sc_hd__nor2_2
XFILLER_149_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_297_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23350_ _23541_/CLK _23350_/D vssd1 vssd1 vccd1 vccd1 _23350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20562_ _20996_/A _21085_/A vssd1 vssd1 vccd1 vccd1 _20779_/B sky130_fd_sc_hd__nor2_1
XFILLER_192_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22301_ _23566_/CLK _22301_/D vssd1 vssd1 vccd1 vccd1 _22301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_354_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23281_ _23537_/CLK _23281_/D vssd1 vssd1 vccd1 vccd1 _23281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20493_ _21077_/C _20493_/B vssd1 vssd1 vccd1 vccd1 _20493_/Y sky130_fd_sc_hd__nor2_1
XFILLER_307_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22232_ _22232_/A _22232_/B vssd1 vssd1 vccd1 vccd1 _22232_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_306_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_307_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_322_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22163_ _22176_/A _22163_/B vssd1 vssd1 vccd1 vccd1 _22163_/X sky130_fd_sc_hd__xor2_4
XFILLER_322_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_322_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21114_ _23853_/Q _21110_/X _21111_/X _20605_/A vssd1 vssd1 vccd1 vccd1 _21115_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_133_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22094_ _13960_/X _22077_/X _22084_/X _22093_/Y vssd1 vssd1 vccd1 vccd1 _22094_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_6939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21045_ _23833_/Q _21048_/B vssd1 vssd1 vccd1 vccd1 _21045_/X sky130_fd_sc_hd__or2_1
XFILLER_259_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_290_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22996_ _23008_/CLK _22996_/D vssd1 vssd1 vccd1 vccd1 _22996_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_227_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21947_ _21947_/A _21947_/B vssd1 vssd1 vccd1 vccd1 _21947_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_43_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11700_/A vssd1 vssd1 vccd1 vccd1 _11700_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12680_/A vssd1 vssd1 vccd1 vccd1 _12680_/X sky130_fd_sc_hd__buf_6
XFILLER_243_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21878_ _21853_/B _21876_/X _21877_/Y vssd1 vssd1 vccd1 vccd1 _21879_/B sky130_fd_sc_hd__o21a_1
XFILLER_230_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11631_ _11631_/A vssd1 vssd1 vccd1 vccd1 _11631_/X sky130_fd_sc_hd__buf_2
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23617_ _23624_/CLK _23617_/D vssd1 vssd1 vccd1 vccd1 _23617_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20829_ _20865_/A vssd1 vssd1 vccd1 vccd1 _20829_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_357_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11562_ _23900_/Q vssd1 vssd1 vccd1 vccd1 _11701_/A sky130_fd_sc_hd__clkbuf_4
X_14350_ _13508_/B _13319_/B _15171_/A vssd1 vssd1 vccd1 vccd1 _14350_/X sky130_fd_sc_hd__mux2_1
XFILLER_356_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23548_ _23548_/CLK _23548_/D vssd1 vssd1 vccd1 vccd1 _23548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_357_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_345_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13301_ _13301_/A _16054_/A vssd1 vssd1 vccd1 vccd1 _13565_/A sky130_fd_sc_hd__nor2_2
XFILLER_357_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14281_ _14281_/A vssd1 vssd1 vccd1 vccd1 _14317_/S sky130_fd_sc_hd__buf_2
X_23479_ _23511_/CLK _23479_/D vssd1 vssd1 vccd1 vccd1 _23479_/Q sky130_fd_sc_hd__dfxtp_4
X_11493_ _22483_/Q _22643_/Q _11493_/S vssd1 vssd1 vccd1 vccd1 _11493_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16020_ _23616_/Q _14732_/X _14734_/X _23648_/Q vssd1 vssd1 vccd1 vccd1 _16020_/X
+ sky130_fd_sc_hd__o22a_2
X_13232_ _13225_/X _13227_/X _13229_/X _13231_/X _11379_/A vssd1 vssd1 vccd1 vccd1
+ _13232_/X sky130_fd_sc_hd__a221o_1
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_298_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13163_ _13212_/A _13163_/B vssd1 vssd1 vccd1 vccd1 _13163_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12114_ _22369_/Q _22401_/Q _22690_/Q _23057_/Q _11151_/A _11953_/A vssd1 vssd1 vccd1
+ vccd1 _12115_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_298_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17971_ _17971_/A vssd1 vssd1 vccd1 vccd1 _18052_/A sky130_fd_sc_hd__buf_4
X_13094_ _23231_/Q _23199_/Q _23167_/Q _23135_/Q _13088_/S _11207_/A vssd1 vssd1 vccd1
+ vccd1 _13095_/B sky130_fd_sc_hd__mux4_1
XFILLER_301_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_297_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_306_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19710_ _19178_/X _23497_/Q _19710_/S vssd1 vssd1 vccd1 vccd1 _19711_/A sky130_fd_sc_hd__mux2_1
X_12045_ _12041_/X _12042_/X _12044_/X vssd1 vssd1 vccd1 vccd1 _12045_/Y sky130_fd_sc_hd__a21oi_1
X_16922_ _17091_/A vssd1 vssd1 vccd1 vccd1 _16922_/X sky130_fd_sc_hd__buf_2
XFILLER_312_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19641_ _19181_/X _23466_/Q _19649_/S vssd1 vssd1 vccd1 vccd1 _19642_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16853_ _16853_/A vssd1 vssd1 vccd1 vccd1 _22532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15804_ _23610_/Q _14450_/A _14455_/A _23642_/Q vssd1 vssd1 vccd1 vccd1 _15804_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_93_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19572_ _19572_/A vssd1 vssd1 vccd1 vccd1 _23435_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16784_ _16784_/A vssd1 vssd1 vccd1 vccd1 _16784_/X sky130_fd_sc_hd__clkbuf_2
X_13996_ _14000_/A _14091_/A vssd1 vssd1 vccd1 vccd1 _13996_/Y sky130_fd_sc_hd__nor2_4
XFILLER_322_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18523_ _18520_/X _18522_/Y _18516_/X vssd1 vssd1 vccd1 vccd1 _23003_/D sky130_fd_sc_hd__a21oi_1
XFILLER_322_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15735_ _15735_/A _15735_/B vssd1 vssd1 vccd1 vccd1 _15735_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ _22797_/Q _22765_/Q _22666_/Q _22733_/Q _12733_/X _12734_/X vssd1 vssd1 vccd1
+ vccd1 _12947_/X sky130_fd_sc_hd__mux4_2
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _18534_/B vssd1 vssd1 vccd1 vccd1 _18465_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15666_ _14703_/X _21861_/A _15665_/X vssd1 vssd1 vccd1 vccd1 _18827_/A sky130_fd_sc_hd__a21o_4
X_12878_ _22378_/Q _22410_/Q _22699_/Q _23066_/Q _12692_/X _11594_/A vssd1 vssd1 vccd1
+ vccd1 _12878_/X sky130_fd_sc_hd__mux4_2
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _17405_/A vssd1 vssd1 vccd1 vccd1 _22615_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ _22915_/Q vssd1 vssd1 vccd1 vccd1 _18263_/B sky130_fd_sc_hd__buf_2
XFILLER_33_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18385_ _18401_/A _18385_/B _18386_/B vssd1 vssd1 vccd1 vccd1 _22955_/D sky130_fd_sc_hd__nor3_1
X_11829_ _11763_/B _21616_/A _11828_/X vssd1 vssd1 vccd1 vccd1 _11939_/B sky130_fd_sc_hd__o21a_4
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15597_ _16171_/S vssd1 vssd1 vccd1 vccd1 _16103_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ _17336_/A vssd1 vssd1 vccd1 vccd1 _22590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14548_ _23886_/Q vssd1 vssd1 vccd1 vccd1 _14548_/X sky130_fd_sc_hd__buf_8
XFILLER_267_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_308_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_131_wb_clk_i _22899_/CLK vssd1 vssd1 vccd1 vccd1 _22923_/CLK sky130_fd_sc_hd__clkbuf_16
X_17267_ _17267_/A vssd1 vssd1 vccd1 vccd1 _22114_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_336_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14479_ _20770_/A _14595_/B vssd1 vssd1 vccd1 vccd1 _14910_/A sky130_fd_sc_hd__nor2_2
XFILLER_347_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19006_ _16899_/X _23199_/Q _19012_/S vssd1 vssd1 vccd1 vccd1 _19007_/A sky130_fd_sc_hd__mux2_1
X_16218_ _22296_/Q _16217_/X _16221_/S vssd1 vssd1 vccd1 vccd1 _16219_/A sky130_fd_sc_hd__mux2_1
XFILLER_351_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_350_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17198_ _22572_/Q _17141_/X _17190_/X _17197_/X vssd1 vssd1 vccd1 vccd1 _22572_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_127_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_344_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_304_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16149_ _23941_/Q vssd1 vssd1 vccd1 vccd1 _22216_/A sky130_fd_sc_hd__buf_2
XFILLER_114_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_303_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19908_ _19908_/A vssd1 vssd1 vccd1 vccd1 _23585_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19839_ _23555_/Q _19261_/A _19841_/S vssd1 vssd1 vccd1 vccd1 _19840_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22850_ _23426_/CLK _22850_/D vssd1 vssd1 vccd1 vccd1 _22850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21801_ _21801_/A _21801_/B _21801_/C _21801_/D vssd1 vssd1 vccd1 vccd1 _21803_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_271_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22781_ _23561_/CLK _22781_/D vssd1 vssd1 vccd1 vccd1 _22781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21732_ _23826_/Q _23760_/Q vssd1 vssd1 vccd1 vccd1 _21733_/B sky130_fd_sc_hd__nor2_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_358_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21663_ _21663_/A vssd1 vssd1 vccd1 vccd1 _22234_/A sky130_fd_sc_hd__buf_2
XFILLER_339_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20614_ _23724_/Q _20593_/X _20613_/X _20602_/X vssd1 vssd1 vccd1 vccd1 _23724_/D
+ sky130_fd_sc_hd__o211a_1
X_23402_ _23466_/CLK _23402_/D vssd1 vssd1 vccd1 vccd1 _23402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21594_ _21594_/A _21594_/B vssd1 vssd1 vccd1 vccd1 _21594_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23333_ _23525_/CLK _23333_/D vssd1 vssd1 vccd1 vccd1 _23333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20545_ _20774_/A vssd1 vssd1 vccd1 vccd1 _20891_/A sky130_fd_sc_hd__buf_4
XFILLER_124_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_354_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_353_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23264_ _23264_/CLK _23264_/D vssd1 vssd1 vccd1 vccd1 _23264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20476_ _23709_/Q _20487_/B vssd1 vssd1 vccd1 vccd1 _20476_/X sky130_fd_sc_hd__or2_1
XFILLER_119_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_335_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_307_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22215_ _22215_/A _22215_/B vssd1 vssd1 vccd1 vccd1 _22215_/Y sky130_fd_sc_hd__nand2_1
XFILLER_335_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23195_ _23419_/CLK _23195_/D vssd1 vssd1 vccd1 vccd1 _23195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22146_ _22146_/A _22146_/B _22146_/C _21410_/A vssd1 vssd1 vccd1 vccd1 _22146_/X
+ sky130_fd_sc_hd__or4b_1
XTAP_6714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput370 _13679_/Y vssd1 vssd1 vccd1 vccd1 csb0[0] sky130_fd_sc_hd__buf_2
XFILLER_294_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput381 _14042_/X vssd1 vssd1 vccd1 vccd1 din0[16] sky130_fd_sc_hd__buf_2
XTAP_6747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput392 _14062_/X vssd1 vssd1 vccd1 vccd1 din0[26] sky130_fd_sc_hd__buf_2
XTAP_6758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22077_ _21613_/X _22076_/Y _21560_/X _23806_/Q vssd1 vssd1 vccd1 vccd1 _22077_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_6769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_294_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21028_ _23826_/Q _21028_/B vssd1 vssd1 vccd1 vccd1 _21028_/X sky130_fd_sc_hd__or2_1
XFILLER_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13850_ _13861_/A _14061_/C vssd1 vssd1 vccd1 vccd1 _13850_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12801_ _12801_/A _21871_/A vssd1 vssd1 vccd1 vccd1 _12801_/X sky130_fd_sc_hd__or2_2
XFILLER_56_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13781_ _13781_/A vssd1 vssd1 vccd1 vccd1 _13781_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22979_ _23424_/CLK _22979_/D vssd1 vssd1 vccd1 vccd1 _22979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_409 _14007_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_308_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15520_ _13775_/A _15478_/X _15479_/Y _15518_/Y _16195_/S vssd1 vssd1 vccd1 vccd1
+ _15520_/X sky130_fd_sc_hd__a221o_1
X_12732_ _12995_/A _12732_/B vssd1 vssd1 vccd1 vccd1 _12732_/X sky130_fd_sc_hd__or2_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15451_ _22927_/Q _15903_/B _15439_/X _15450_/Y _14897_/A vssd1 vssd1 vccd1 vccd1
+ _15451_/X sky130_fd_sc_hd__a221o_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12663_ _12636_/X _12664_/A vssd1 vssd1 vccd1 vccd1 _12665_/A sky130_fd_sc_hd__and2b_2
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _22898_/Q _14160_/X _16929_/A _22591_/Q vssd1 vssd1 vccd1 vccd1 _16936_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18170_ _18165_/X _18179_/A _18168_/X _18169_/X vssd1 vssd1 vccd1 vccd1 _18170_/X
+ sky130_fd_sc_hd__a31o_1
X_11614_ _22278_/Q _23094_/Q _23510_/Q _22439_/Q _12043_/S _11613_/X vssd1 vssd1 vccd1
+ vccd1 _11615_/B sky130_fd_sc_hd__mux4_1
X_15382_ _13833_/A _15380_/Y _15381_/Y _13737_/A vssd1 vssd1 vccd1 vccd1 _15382_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_129_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_357_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12594_ _12594_/A _12594_/B _12594_/C vssd1 vssd1 vccd1 vccd1 _21422_/A sky130_fd_sc_hd__and3_4
XFILLER_11_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17121_ input82/X input47/X _17132_/S vssd1 vssd1 vccd1 vccd1 _17121_/X sky130_fd_sc_hd__mux2_8
XFILLER_184_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14333_ _14333_/A vssd1 vssd1 vccd1 vccd1 _14333_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11545_ _22386_/Q _22418_/Q _22707_/Q _23074_/Q _11543_/X _13276_/A vssd1 vssd1 vccd1
+ vccd1 _11545_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17052_ _17052_/A vssd1 vssd1 vccd1 vccd1 _17052_/Y sky130_fd_sc_hd__inv_2
XFILLER_333_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11476_ _15630_/A _11476_/B vssd1 vssd1 vccd1 vccd1 _11476_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14264_ _16097_/A vssd1 vssd1 vccd1 vccd1 _14264_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16003_ _16003_/A _16039_/C vssd1 vssd1 vccd1 vccd1 _16004_/B sky130_fd_sc_hd__xnor2_4
X_13215_ _22381_/Q _22413_/Q _22702_/Q _23069_/Q _11526_/A _11519_/A vssd1 vssd1 vccd1
+ vccd1 _13216_/B sky130_fd_sc_hd__mux4_1
X_14195_ _14195_/A vssd1 vssd1 vccd1 vccd1 _14195_/X sky130_fd_sc_hd__buf_4
XFILLER_325_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13146_ _11195_/A _13145_/X _13206_/A vssd1 vssd1 vccd1 vccd1 _13146_/X sky130_fd_sc_hd__a21o_1
XFILLER_98_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_301_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17954_ _22828_/Q _17938_/X _17939_/X input274/X _17951_/X vssd1 vssd1 vccd1 vccd1
+ _17954_/X sky130_fd_sc_hd__a221o_1
X_13077_ _11278_/A _13067_/X _13076_/X _13295_/A vssd1 vssd1 vccd1 vccd1 _20374_/A
+ sky130_fd_sc_hd__a211o_4
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12028_ _12028_/A vssd1 vssd1 vccd1 vccd1 _12708_/A sky130_fd_sc_hd__buf_2
X_16905_ _19255_/A vssd1 vssd1 vccd1 vccd1 _16905_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_238_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17885_ _22893_/Q _22892_/Q vssd1 vssd1 vccd1 vccd1 _18172_/A sky130_fd_sc_hd__or2_1
XFILLER_239_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19624_ _19624_/A vssd1 vssd1 vccd1 vccd1 _23459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16836_ _16835_/X _22527_/Q _16845_/S vssd1 vssd1 vccd1 vccd1 _16837_/A sky130_fd_sc_hd__mux2_1
XFILLER_254_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19555_ _19555_/A _19555_/B vssd1 vssd1 vccd1 vccd1 _19612_/A sky130_fd_sc_hd__nor2_8
X_16767_ _22507_/Q _16765_/X _16766_/X input22/X vssd1 vssd1 vccd1 vccd1 _16768_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13979_ _13979_/A _13979_/B vssd1 vssd1 vccd1 vccd1 _13980_/A sky130_fd_sc_hd__and2_1
XFILLER_202_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18506_ _18494_/X _18505_/Y _18503_/X vssd1 vssd1 vccd1 vccd1 _22997_/D sky130_fd_sc_hd__a21oi_1
XFILLER_234_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15718_ _15718_/A _15718_/B vssd1 vssd1 vccd1 vccd1 _15718_/Y sky130_fd_sc_hd__nor2_1
XFILLER_179_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19486_ _19163_/X _23397_/Q _19494_/S vssd1 vssd1 vccd1 vccd1 _19487_/A sky130_fd_sc_hd__mux2_1
X_16698_ _16704_/A _16698_/B vssd1 vssd1 vccd1 vccd1 _16699_/A sky130_fd_sc_hd__or2_1
X_18437_ _22974_/Q _18440_/C vssd1 vssd1 vccd1 vccd1 _18438_/B sky130_fd_sc_hd__and2_1
XFILLER_222_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15649_ _23766_/Q _14911_/X _14913_/X _15647_/X _15648_/X vssd1 vssd1 vccd1 vccd1
+ _15649_/X sky130_fd_sc_hd__a221o_1
XFILLER_221_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_349_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18368_ _19962_/A vssd1 vssd1 vccd1 vccd1 _18403_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_336_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17319_ _17245_/A _17318_/X _16996_/A _17283_/X vssd1 vssd1 vccd1 vccd1 _17319_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18299_ _18307_/D vssd1 vssd1 vccd1 vccd1 _18305_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20330_ _20302_/X _20328_/X _20329_/Y _21954_/A _20307_/X vssd1 vssd1 vccd1 vccd1
+ _20700_/A sky130_fd_sc_hd__a32o_4
XFILLER_335_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_350_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20261_ _20295_/A vssd1 vssd1 vccd1 vccd1 _20261_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22000_ _22000_/A _22000_/B vssd1 vssd1 vccd1 vccd1 _22002_/A sky130_fd_sc_hd__nand2_1
XFILLER_350_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20192_ _20307_/A vssd1 vssd1 vccd1 vccd1 _20192_/X sky130_fd_sc_hd__buf_2
XFILLER_103_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput109 dout1[11] vssd1 vssd1 vccd1 vccd1 input109/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23951_ _23951_/A vssd1 vssd1 vccd1 vccd1 _23951_/X sky130_fd_sc_hd__buf_2
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22902_ _22908_/CLK _22902_/D vssd1 vssd1 vccd1 vccd1 _22902_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23882_ _23926_/CLK _23882_/D vssd1 vssd1 vccd1 vccd1 _23882_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_256_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22833_ _22893_/CLK _22833_/D vssd1 vssd1 vccd1 vccd1 _22833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22764_ _23450_/CLK _22764_/D vssd1 vssd1 vccd1 vccd1 _22764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21715_ _15377_/X _21479_/X _21699_/Y _21714_/Y _21681_/X vssd1 vssd1 vccd1 vccd1
+ _23923_/D sky130_fd_sc_hd__o221a_1
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22695_ _22695_/CLK _22695_/D vssd1 vssd1 vccd1 vccd1 _22695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21646_ _14548_/X _21518_/X _21336_/B _21868_/A _21925_/A vssd1 vssd1 vccd1 vccd1
+ _21646_/X sky130_fd_sc_hd__a32o_1
XFILLER_185_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_327_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_355_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21577_ _21767_/A vssd1 vssd1 vccd1 vccd1 _21577_/X sky130_fd_sc_hd__buf_2
XFILLER_126_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11330_ _11330_/A vssd1 vssd1 vccd1 vccd1 _11863_/A sky130_fd_sc_hd__clkbuf_8
X_23316_ _23542_/CLK _23316_/D vssd1 vssd1 vccd1 vccd1 _23316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20528_ _14713_/C _21289_/A _21313_/B _21605_/B _21357_/C vssd1 vssd1 vccd1 vccd1
+ _20528_/X sky130_fd_sc_hd__a41o_2
XFILLER_338_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_326_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11261_ _23909_/Q _11080_/A _14180_/D _23908_/Q _23910_/Q vssd1 vssd1 vccd1 vccd1
+ _14371_/B sky130_fd_sc_hd__a2111o_4
X_23247_ _23535_/CLK _23247_/D vssd1 vssd1 vccd1 vccd1 _23247_/Q sky130_fd_sc_hd__dfxtp_1
X_20459_ _20602_/A vssd1 vssd1 vccd1 vccd1 _20459_/X sky130_fd_sc_hd__buf_2
XFILLER_354_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_7212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13000_ _12745_/A _12993_/X _12995_/X _12999_/X _11379_/A vssd1 vssd1 vccd1 vccd1
+ _13010_/B sky130_fd_sc_hd__a311o_2
XTAP_7234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_341_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11192_ _11837_/A vssd1 vssd1 vccd1 vccd1 _12071_/A sky130_fd_sc_hd__buf_4
X_23178_ _23370_/CLK _23178_/D vssd1 vssd1 vccd1 vccd1 _23178_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_7245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22129_ _22129_/A _22128_/Y vssd1 vssd1 vccd1 vccd1 _22129_/X sky130_fd_sc_hd__or2b_1
XTAP_7289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_294_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14951_ _14951_/A vssd1 vssd1 vccd1 vccd1 _14951_/Y sky130_fd_sc_hd__inv_2
XTAP_6599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13902_ _14794_/A _13902_/B vssd1 vssd1 vccd1 vccd1 _13903_/B sky130_fd_sc_hd__nand2_1
XTAP_5887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17670_ _17670_/A vssd1 vssd1 vccd1 vccd1 _22716_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14882_ _14882_/A vssd1 vssd1 vccd1 vccd1 _14882_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_291_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16621_ _22459_/Q _16223_/X _16629_/S vssd1 vssd1 vccd1 vccd1 _16622_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13833_ _13833_/A vssd1 vssd1 vccd1 vccd1 _13834_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_303_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_206 _14393_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_217 _14827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19340_ _19396_/A vssd1 vssd1 vccd1 vccd1 _19409_/S sky130_fd_sc_hd__buf_6
XFILLER_16_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16552_ _16552_/A vssd1 vssd1 vccd1 vccd1 _22428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_228 _15107_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13764_ _13764_/A _14074_/A vssd1 vssd1 vccd1 vccd1 _13815_/B sky130_fd_sc_hd__or2_1
XINSDIODE2_239 _15223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15503_ _23603_/Q vssd1 vssd1 vccd1 vccd1 _19976_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12715_ _12995_/A _12715_/B vssd1 vssd1 vccd1 vccd1 _12715_/X sky130_fd_sc_hd__or2_1
X_19271_ _19271_/A vssd1 vssd1 vccd1 vccd1 _23301_/D sky130_fd_sc_hd__clkbuf_1
X_16483_ _15324_/X _22399_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _16484_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13695_ _13779_/A _13695_/B _19969_/D vssd1 vssd1 vccd1 vccd1 _14006_/C sky130_fd_sc_hd__and3_2
XFILLER_31_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18222_ _22852_/Q _18216_/X _18221_/X _18219_/X vssd1 vssd1 vccd1 vccd1 _22900_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_188_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15434_ _13833_/A _15432_/Y _15433_/Y _13738_/A vssd1 vssd1 vccd1 vccd1 _15434_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12646_ _12656_/A vssd1 vssd1 vccd1 vccd1 _12759_/A sky130_fd_sc_hd__clkbuf_4
XPHY_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_321_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_318_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_321_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_317_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18153_ _18476_/A _18153_/B vssd1 vssd1 vccd1 vccd1 _18154_/A sky130_fd_sc_hd__or2_1
XFILLER_200_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15365_ _15775_/A vssd1 vssd1 vccd1 vccd1 _15365_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12577_ _12586_/A _12577_/B vssd1 vssd1 vccd1 vccd1 _12577_/X sky130_fd_sc_hd__or2_1
XFILLER_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17104_ _23472_/Q _17061_/X _17062_/X _17094_/X _17103_/Y vssd1 vssd1 vccd1 vccd1
+ _17104_/X sky130_fd_sc_hd__a32o_1
XFILLER_117_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14316_ _13028_/A _13340_/B _14317_/S vssd1 vssd1 vccd1 vccd1 _14316_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18084_ _18099_/A vssd1 vssd1 vccd1 vccd1 _18084_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_318_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11528_ _23490_/Q _23586_/Q _22550_/Q _22354_/Q _13275_/A _11527_/X vssd1 vssd1 vccd1
+ vccd1 _11529_/B sky130_fd_sc_hd__mux4_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15296_ _14839_/A _15801_/B _15798_/B _15801_/A _15295_/Y vssd1 vssd1 vccd1 vccd1
+ _15296_/X sky130_fd_sc_hd__o221a_2
XFILLER_116_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_305_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17035_ _16940_/X _17648_/B _16947_/X _17024_/X _17034_/X vssd1 vssd1 vccd1 vccd1
+ _17035_/X sky130_fd_sc_hd__a311o_1
XFILLER_7_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14247_ _14247_/A vssd1 vssd1 vccd1 vccd1 _14247_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_332_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11459_ _12634_/A vssd1 vssd1 vccd1 vccd1 _13295_/A sky130_fd_sc_hd__buf_12
XFILLER_264_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14178_ _14178_/A vssd1 vssd1 vccd1 vccd1 _21925_/A sky130_fd_sc_hd__buf_6
XFILLER_112_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13129_ _13117_/A _13128_/X _12745_/X vssd1 vssd1 vccd1 vccd1 _13129_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_301_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18986_ _16870_/X _23190_/Q _18990_/S vssd1 vssd1 vccd1 vccd1 _18987_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_301_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17937_ _22824_/Q _17932_/X _17936_/X _17930_/X vssd1 vssd1 vccd1 vccd1 _22824_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17868_ _22805_/Q _17636_/X _17870_/S vssd1 vssd1 vccd1 vccd1 _17869_/A sky130_fd_sc_hd__mux2_1
XFILLER_253_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19607_ _19607_/A vssd1 vssd1 vccd1 vccd1 _23451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16819_ _19169_/A vssd1 vssd1 vccd1 vccd1 _16819_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17799_ _17799_/A vssd1 vssd1 vccd1 vccd1 _22774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19538_ _19242_/X _23421_/Q _19538_/S vssd1 vssd1 vccd1 vccd1 _19539_/A sky130_fd_sc_hd__mux2_1
XFILLER_253_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19469_ _23390_/Q _18852_/X _19477_/S vssd1 vssd1 vccd1 vccd1 _19470_/A sky130_fd_sc_hd__mux2_1
XFILLER_250_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21500_ _21500_/A _21500_/B vssd1 vssd1 vccd1 vccd1 _21501_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22480_ _23583_/CLK _22480_/D vssd1 vssd1 vccd1 vccd1 _22480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_309_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21431_ _21431_/A _21437_/A vssd1 vssd1 vccd1 vccd1 _21472_/A sky130_fd_sc_hd__nor2_1
XFILLER_337_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21362_ _21465_/A vssd1 vssd1 vccd1 vccd1 _22093_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_3_1_1_wb_clk_i clkbuf_3_1_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_308_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23101_ _23547_/CLK _23101_/D vssd1 vssd1 vccd1 vccd1 _23101_/Q sky130_fd_sc_hd__dfxtp_1
X_20313_ _20376_/A _20313_/B vssd1 vssd1 vccd1 vccd1 _20313_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput80 dout0[43] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__clkbuf_1
X_21293_ _21293_/A _21320_/B vssd1 vssd1 vccd1 vccd1 _21293_/Y sky130_fd_sc_hd__nor2_1
Xinput91 dout0[53] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23032_ _23354_/CLK _23032_/D vssd1 vssd1 vccd1 vccd1 _23032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_323_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20244_ _20187_/X _20242_/X _20243_/Y _21594_/A _20200_/X vssd1 vssd1 vccd1 vccd1
+ _20622_/A sky130_fd_sc_hd__a32o_4
XFILLER_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20175_ _20355_/A _20171_/X _20174_/X vssd1 vssd1 vccd1 vccd1 _20175_/X sky130_fd_sc_hd__a21o_1
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23934_ _23934_/CLK _23934_/D vssd1 vssd1 vccd1 vccd1 _23934_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_229_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23865_ _23918_/CLK _23865_/D vssd1 vssd1 vccd1 vccd1 _23865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22816_ _22830_/CLK _22816_/D vssd1 vssd1 vccd1 vccd1 _22816_/Q sky130_fd_sc_hd__dfxtp_1
X_23796_ _23942_/CLK _23796_/D vssd1 vssd1 vccd1 vccd1 _23796_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_344_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22747_ _22779_/CLK _22747_/D vssd1 vssd1 vccd1 vccd1 _22747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12500_ _12506_/A _12500_/B vssd1 vssd1 vccd1 vccd1 _12500_/X sky130_fd_sc_hd__or2_1
XFILLER_347_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13480_ _13890_/A _13882_/A _13479_/X vssd1 vssd1 vccd1 vccd1 _13481_/B sky130_fd_sc_hd__o21a_2
XFILLER_232_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22678_ _23555_/CLK _22678_/D vssd1 vssd1 vccd1 vccd1 _22678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12431_ _12570_/A _12431_/B vssd1 vssd1 vccd1 vccd1 _12431_/Y sky130_fd_sc_hd__nor2_1
XFILLER_200_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21629_ _21627_/Y _21629_/B vssd1 vssd1 vccd1 vccd1 _21632_/A sky130_fd_sc_hd__and2b_1
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15150_ _15150_/A vssd1 vssd1 vccd1 vccd1 _15150_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12362_ _23464_/Q _23560_/Q _22524_/Q _22328_/Q _11112_/A _11702_/A vssd1 vssd1 vccd1
+ vccd1 _12362_/X sky130_fd_sc_hd__mux4_1
XFILLER_343_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14101_ _22890_/Q vssd1 vssd1 vccd1 vccd1 _18178_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_299_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11313_ _23895_/Q vssd1 vssd1 vccd1 vccd1 _12476_/A sky130_fd_sc_hd__buf_2
X_12293_ _22362_/Q _22394_/Q _22683_/Q _23050_/Q _12349_/S _12292_/X vssd1 vssd1 vccd1
+ vccd1 _12293_/X sky130_fd_sc_hd__mux4_1
X_15081_ _15081_/A _15081_/B vssd1 vssd1 vccd1 vccd1 _15583_/A sky130_fd_sc_hd__or2_4
XFILLER_180_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_299_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_302_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11244_ _11244_/A vssd1 vssd1 vccd1 vccd1 _11559_/A sky130_fd_sc_hd__clkbuf_4
X_14032_ _14046_/A _14052_/B _14032_/C vssd1 vssd1 vccd1 vccd1 _14032_/X sky130_fd_sc_hd__or3_1
XFILLER_351_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18840_ _18840_/A vssd1 vssd1 vccd1 vccd1 _18840_/X sky130_fd_sc_hd__clkbuf_2
X_11175_ _12532_/A vssd1 vssd1 vccd1 vccd1 _12307_/A sky130_fd_sc_hd__clkbuf_4
XTAP_7075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_7097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18771_ _19555_/B _19018_/B vssd1 vssd1 vccd1 vccd1 _18853_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15983_ _23615_/Q vssd1 vssd1 vccd1 vccd1 _20016_/B sky130_fd_sc_hd__buf_2
XTAP_5640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_310_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17722_ _22740_/Q _17633_/X _17726_/S vssd1 vssd1 vccd1 vccd1 _17723_/A sky130_fd_sc_hd__mux2_1
XTAP_5662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14934_ _15001_/A vssd1 vssd1 vccd1 vccd1 _14934_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17653_ _17653_/A _17653_/B vssd1 vssd1 vccd1 vccd1 _17653_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14865_ _14865_/A _15335_/B vssd1 vssd1 vccd1 vccd1 _14865_/Y sky130_fd_sc_hd__nor2_1
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16604_ _16604_/A vssd1 vssd1 vccd1 vccd1 _22452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_250_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13816_ _13790_/X _13864_/A _13814_/Y _13863_/A vssd1 vssd1 vccd1 vccd1 _13817_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_223_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17584_ _17584_/A vssd1 vssd1 vccd1 vccd1 _22689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14796_ _14794_/B _14676_/B _14942_/A _14794_/Y _15636_/A vssd1 vssd1 vccd1 vccd1
+ _14796_/X sky130_fd_sc_hd__o221a_1
XFILLER_90_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19323_ _19323_/A vssd1 vssd1 vccd1 vccd1 _23325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_251_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16535_ _19699_/A _19771_/A vssd1 vssd1 vccd1 vccd1 _16592_/A sky130_fd_sc_hd__or2_4
XFILLER_16_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_330_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13747_ _13793_/B _13739_/X _13842_/A _13746_/X vssd1 vssd1 vccd1 vccd1 _13748_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_188_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19254_ _19254_/A vssd1 vssd1 vccd1 vccd1 _23296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16466_ _16466_/A vssd1 vssd1 vccd1 vccd1 _22391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13678_ _13678_/A vssd1 vssd1 vccd1 vccd1 _13678_/X sky130_fd_sc_hd__clkbuf_1
X_18205_ _22894_/Q _18214_/B vssd1 vssd1 vccd1 vccd1 _18205_/X sky130_fd_sc_hd__or2_1
XFILLER_339_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15417_ _15417_/A vssd1 vssd1 vccd1 vccd1 _15621_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12629_ _22793_/Q _22761_/Q _22662_/Q _22729_/Q _12024_/X _12025_/X vssd1 vssd1 vccd1
+ vccd1 _12630_/B sky130_fd_sc_hd__mux4_1
XPHY_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19185_ _19185_/A vssd1 vssd1 vccd1 vccd1 _19185_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_192_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16397_ _16397_/A vssd1 vssd1 vccd1 vccd1 _22361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_319_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18136_ _18198_/A _18138_/A _22884_/Q vssd1 vssd1 vccd1 vccd1 _18136_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_38_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23571_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_200_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15348_ _22957_/Q vssd1 vssd1 vccd1 vccd1 _15351_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_191_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_334_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18067_ _18097_/A vssd1 vssd1 vccd1 vccd1 _18067_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15279_ _22987_/Q _15416_/A _15417_/A input246/X vssd1 vssd1 vccd1 vccd1 _15280_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_144_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17018_ _23464_/Q _17016_/X _17017_/X _17042_/A _14879_/X vssd1 vssd1 vccd1 vccd1
+ _17018_/X sky130_fd_sc_hd__a32o_1
XFILLER_99_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_302_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18969_ _18969_/A vssd1 vssd1 vccd1 vccd1 _23182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_287_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21980_ _21569_/X _21978_/X _21979_/Y _21577_/X vssd1 vssd1 vccd1 vccd1 _21981_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_273_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20931_ _15377_/X _20922_/X _20652_/B _20926_/X vssd1 vssd1 vccd1 vccd1 _20931_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_270_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23650_ _23651_/CLK _23650_/D vssd1 vssd1 vccd1 vccd1 _23650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20862_ _20862_/A vssd1 vssd1 vccd1 vccd1 _23772_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22601_ _23649_/CLK _22601_/D vssd1 vssd1 vccd1 vccd1 _22601_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_23581_ _23581_/CLK _23581_/D vssd1 vssd1 vccd1 vccd1 _23581_/Q sky130_fd_sc_hd__dfxtp_2
X_20793_ _20591_/B _20791_/X _20792_/X _23753_/Q vssd1 vssd1 vccd1 vccd1 _20794_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22532_ _23504_/CLK _22532_/D vssd1 vssd1 vccd1 vccd1 _22532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_329_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22463_ _23566_/CLK _22463_/D vssd1 vssd1 vccd1 vccd1 _22463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_325_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21414_ _23817_/Q _23751_/Q vssd1 vssd1 vccd1 vccd1 _21416_/A sky130_fd_sc_hd__nor2_1
X_22394_ _23564_/CLK _22394_/D vssd1 vssd1 vccd1 vccd1 _22394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_324_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21345_ _21345_/A _21345_/B vssd1 vssd1 vccd1 vccd1 _21345_/X sky130_fd_sc_hd__or2_1
XFILLER_351_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_324_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_352_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_324_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21276_ _21276_/A _21283_/B vssd1 vssd1 vccd1 vccd1 _21276_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_340_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20227_ _20305_/A vssd1 vssd1 vccd1 vccd1 _20227_/X sky130_fd_sc_hd__clkbuf_2
X_23015_ _23555_/CLK _23015_/D vssd1 vssd1 vccd1 vccd1 _23015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_270_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_289_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20158_ _20147_/X _17655_/A _20157_/X vssd1 vssd1 vccd1 vccd1 _20543_/A sky130_fd_sc_hd__o21ai_4
XFILLER_351_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_311_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20089_ _23638_/Q vssd1 vssd1 vccd1 vccd1 _20098_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_292_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12980_ _13195_/A _12977_/X _12979_/X vssd1 vssd1 vccd1 vccd1 _12980_/X sky130_fd_sc_hd__a21o_1
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23917_ _23917_/CLK _23917_/D vssd1 vssd1 vccd1 vccd1 _23917_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_100_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11931_ _12318_/A _11931_/B vssd1 vssd1 vccd1 vccd1 _11931_/X sky130_fd_sc_hd__or2_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14650_ _14642_/X _14649_/X _15339_/S vssd1 vssd1 vccd1 vccd1 _15488_/A sky130_fd_sc_hd__mux2_2
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23848_ _23851_/CLK _23848_/D vssd1 vssd1 vccd1 vccd1 _23848_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _23470_/Q _23566_/Q _22530_/Q _22334_/Q _11821_/X _11317_/A vssd1 vssd1 vccd1
+ vccd1 _11863_/B sky130_fd_sc_hd__mux4_1
XFILLER_260_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13601_ _13601_/A _13601_/B vssd1 vssd1 vccd1 vccd1 _13601_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_150_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ input150/X _13651_/B _14719_/S input115/X _14235_/X vssd1 vssd1 vccd1 vccd1
+ _14581_/X sky130_fd_sc_hd__a221o_4
XFILLER_214_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11793_ _12134_/A _11793_/B _11793_/C vssd1 vssd1 vccd1 vccd1 _13752_/A sky130_fd_sc_hd__or3_4
X_23779_ _23866_/CLK _23779_/D vssd1 vssd1 vccd1 vccd1 _23779_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16320_ _14893_/X _22328_/Q _16322_/S vssd1 vssd1 vccd1 vccd1 _16321_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13532_ _13532_/A _13611_/A _13532_/C _13532_/D vssd1 vssd1 vccd1 vccd1 _13532_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_198_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16251_ _16251_/A vssd1 vssd1 vccd1 vccd1 _22306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13463_ _13474_/A vssd1 vssd1 vccd1 vccd1 _13587_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_159_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15202_ _13936_/X _15580_/B _14866_/A vssd1 vssd1 vccd1 vccd1 _15202_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_334_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12414_ _12414_/A _12414_/B _12414_/C vssd1 vssd1 vccd1 vccd1 _21340_/A sky130_fd_sc_hd__nor3_4
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16182_ _11394_/A _14251_/A _14760_/A vssd1 vssd1 vccd1 vccd1 _16182_/X sky130_fd_sc_hd__a21o_1
XFILLER_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_327_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13394_ _13323_/A _13023_/X _13389_/X _15635_/A _13393_/Y vssd1 vssd1 vccd1 vccd1
+ _13395_/D sky130_fd_sc_hd__a311o_2
XFILLER_182_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15133_ _15133_/A _15133_/B vssd1 vssd1 vccd1 vccd1 _15133_/Y sky130_fd_sc_hd__nor2_1
XFILLER_299_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12345_ _14132_/A _12345_/B _14172_/B vssd1 vssd1 vccd1 vccd1 _13775_/D sky130_fd_sc_hd__or3b_1
XFILLER_153_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_299_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19941_ _19950_/A _19971_/B vssd1 vssd1 vccd1 vccd1 _19941_/Y sky130_fd_sc_hd__nor2_1
X_15064_ _22920_/Q _15000_/X _15001_/X _22952_/Q vssd1 vssd1 vccd1 vccd1 _15064_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_114_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12276_ _12401_/A _12275_/X _11819_/X vssd1 vssd1 vccd1 vccd1 _12276_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_142_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14015_ _14015_/A _14036_/B _14015_/C vssd1 vssd1 vccd1 vccd1 _14015_/X sky130_fd_sc_hd__and3_1
XFILLER_268_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11227_ _23902_/Q vssd1 vssd1 vccd1 vccd1 _11705_/A sky130_fd_sc_hd__inv_2
XFILLER_311_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19872_ _16246_/X _23569_/Q _19876_/S vssd1 vssd1 vccd1 vccd1 _19873_/A sky130_fd_sc_hd__mux2_1
XFILLER_268_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18823_ _18823_/A vssd1 vssd1 vccd1 vccd1 _23124_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_311_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_156_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23818_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_122_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11158_ _23900_/Q vssd1 vssd1 vccd1 vccd1 _11189_/A sky130_fd_sc_hd__clkbuf_8
XTAP_6171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_295_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18754_ _18754_/A vssd1 vssd1 vccd1 vccd1 _18763_/S sky130_fd_sc_hd__buf_6
X_15966_ _14215_/A _21269_/A _15965_/Y _16154_/A vssd1 vssd1 vccd1 vccd1 _15966_/X
+ sky130_fd_sc_hd__o211a_1
X_11089_ _23893_/Q _23885_/Q _12345_/B _23884_/Q vssd1 vssd1 vccd1 vccd1 _11090_/C
+ sky130_fd_sc_hd__or4b_1
XTAP_5470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput270 partID[15] vssd1 vssd1 vccd1 vccd1 input270/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput281 versionID[1] vssd1 vssd1 vccd1 vccd1 input281/X sky130_fd_sc_hd__clkbuf_2
XTAP_5492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17705_ _17705_/A vssd1 vssd1 vccd1 vccd1 _22732_/D sky130_fd_sc_hd__clkbuf_1
X_14917_ _14917_/A vssd1 vssd1 vccd1 vccd1 _14917_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18685_ _23071_/Q _17630_/X _18691_/S vssd1 vssd1 vccd1 vccd1 _18686_/A sky130_fd_sc_hd__mux2_1
X_15897_ _18846_/A vssd1 vssd1 vccd1 vccd1 _19239_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17636_ _18862_/A vssd1 vssd1 vccd1 vccd1 _17636_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_223_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14848_ _14848_/A vssd1 vssd1 vccd1 vccd1 _15011_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_263_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17567_ _22684_/Q _17566_/X _17576_/S vssd1 vssd1 vccd1 vccd1 _17568_/A sky130_fd_sc_hd__mux2_1
X_14779_ _15018_/S _14776_/X _14778_/X vssd1 vssd1 vccd1 vccd1 _14779_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_17_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16518_ _16013_/X _22415_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _16519_/A sky130_fd_sc_hd__mux2_1
X_19306_ _19306_/A vssd1 vssd1 vccd1 vccd1 _23317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17498_ _17498_/A vssd1 vssd1 vccd1 vccd1 _22656_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19237_ _19236_/X _23291_/Q _19243_/S vssd1 vssd1 vccd1 vccd1 _19238_/A sky130_fd_sc_hd__mux2_1
X_16449_ _16089_/X _22385_/Q _16451_/S vssd1 vssd1 vccd1 vccd1 _16450_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19168_ _19168_/A vssd1 vssd1 vccd1 vccd1 _23269_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18119_ _18118_/X _14107_/X _22878_/Q vssd1 vssd1 vccd1 vccd1 _18119_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19099_ _19099_/A vssd1 vssd1 vccd1 vccd1 _23239_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_333_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21130_ _21134_/A _21130_/B vssd1 vssd1 vccd1 vccd1 _23859_/D sky130_fd_sc_hd__nor2_1
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21061_ _21163_/A vssd1 vssd1 vccd1 vccd1 _21061_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20012_ _20121_/A vssd1 vssd1 vccd1 vccd1 _20041_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_286_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21963_ _21961_/Y _21963_/B vssd1 vssd1 vccd1 vccd1 _22038_/B sky130_fd_sc_hd__and2b_1
XFILLER_261_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23702_ _23706_/CLK _23702_/D vssd1 vssd1 vccd1 vccd1 _23702_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_254_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20914_ _23786_/Q _20911_/X _20913_/X _20906_/X vssd1 vssd1 vccd1 vccd1 _23786_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_242_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21894_ _21767_/X _21893_/X _21410_/A vssd1 vssd1 vccd1 vccd1 _21894_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_199_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23633_ _23634_/CLK _23633_/D vssd1 vssd1 vccd1 vccd1 _23633_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_243_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20845_ _20881_/A vssd1 vssd1 vccd1 vccd1 _20861_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_154_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23564_ _23564_/CLK _23564_/D vssd1 vssd1 vccd1 vccd1 _23564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20776_ _20811_/A vssd1 vssd1 vccd1 vccd1 _20888_/C sky130_fd_sc_hd__buf_2
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22515_ _23693_/CLK _22515_/D vssd1 vssd1 vccd1 vccd1 _22515_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_356_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23495_ _23896_/CLK _23495_/D vssd1 vssd1 vccd1 vccd1 _23495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22446_ _23515_/CLK _22446_/D vssd1 vssd1 vccd1 vccd1 _22446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22377_ _23451_/CLK _22377_/D vssd1 vssd1 vccd1 vccd1 _22377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_324_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12130_ _12130_/A _12130_/B vssd1 vssd1 vccd1 vccd1 _12130_/Y sky130_fd_sc_hd__nor2_1
XFILLER_163_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21328_ _21328_/A vssd1 vssd1 vccd1 vccd1 _21922_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_352_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_340_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12061_ _12661_/A _13768_/A vssd1 vssd1 vccd1 vccd1 _12061_/Y sky130_fd_sc_hd__nand2_1
X_21259_ _21259_/A vssd1 vssd1 vccd1 vccd1 _23899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_277_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15820_ _14393_/X _15574_/X _15818_/X _15819_/Y _15618_/A vssd1 vssd1 vccd1 vccd1
+ _15820_/X sky130_fd_sc_hd__o221a_1
XFILLER_292_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _15751_/A vssd1 vssd1 vccd1 vccd1 _22280_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ _13022_/A _12964_/B vssd1 vssd1 vccd1 vccd1 _13328_/A sky130_fd_sc_hd__and2_1
XFILLER_46_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_60 _21186_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_71 _13440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14702_ _15519_/A vssd1 vssd1 vccd1 vccd1 _15746_/A sky130_fd_sc_hd__buf_4
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_82 _15616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18470_ _18467_/X _18469_/Y _18463_/X vssd1 vssd1 vccd1 vccd1 _22983_/D sky130_fd_sc_hd__a21oi_1
XINSDIODE2_93 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _11914_/A _11914_/B vssd1 vssd1 vccd1 vccd1 _11914_/X sky130_fd_sc_hd__or2_1
XFILLER_46_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15682_ _14264_/X _15459_/X _15681_/X _14837_/X vssd1 vssd1 vccd1 vccd1 _15682_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12894_ _22378_/Q _22410_/Q _22699_/Q _23066_/Q _12792_/X _12793_/X vssd1 vssd1 vccd1
+ vccd1 _12895_/B sky130_fd_sc_hd__mux4_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _22623_/Q _16236_/X _17421_/S vssd1 vssd1 vccd1 vccd1 _17422_/A sky130_fd_sc_hd__mux2_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14633_ _14298_/X _14300_/X _14651_/A vssd1 vssd1 vccd1 vccd1 _14633_/X sky130_fd_sc_hd__mux2_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11845_ _12291_/A _11841_/X _11844_/X vssd1 vssd1 vccd1 vccd1 _11845_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17352_ _22597_/Q input191/X _17358_/S vssd1 vssd1 vccd1 vccd1 _17353_/A sky130_fd_sc_hd__mux2_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14564_/A vssd1 vssd1 vccd1 vccd1 _15631_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11776_ _11837_/A _11776_/B vssd1 vssd1 vccd1 vccd1 _11776_/Y sky130_fd_sc_hd__nand2_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16303_ _18868_/A vssd1 vssd1 vccd1 vccd1 _16303_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13515_ _13513_/X _12600_/A _13514_/X vssd1 vssd1 vccd1 vccd1 _13516_/B sky130_fd_sc_hd__o21a_1
X_17283_ _17283_/A vssd1 vssd1 vccd1 vccd1 _17283_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14495_ _14500_/A _20770_/A vssd1 vssd1 vccd1 vccd1 _15148_/B sky130_fd_sc_hd__nor2_1
XFILLER_201_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19022_ _19022_/A vssd1 vssd1 vccd1 vccd1 _23205_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16234_ _22301_/Q _16233_/X _16237_/S vssd1 vssd1 vccd1 vccd1 _16235_/A sky130_fd_sc_hd__mux2_1
XFILLER_335_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13446_ _23906_/Q vssd1 vssd1 vccd1 vccd1 _16016_/A sky130_fd_sc_hd__buf_8
XFILLER_357_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16165_ _23942_/Q _16165_/B vssd1 vssd1 vccd1 vccd1 _16165_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_318_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13377_ _13375_/A _13341_/X _13344_/X vssd1 vssd1 vccd1 vccd1 _13378_/B sky130_fd_sc_hd__o21a_1
XFILLER_170_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_336_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15116_ _14247_/A _15114_/X _15115_/X vssd1 vssd1 vccd1 vccd1 _15116_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12328_ _12334_/A vssd1 vssd1 vccd1 vccd1 _12590_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_315_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16096_ _15176_/A _13548_/A _15583_/X _11558_/A _16095_/Y vssd1 vssd1 vccd1 vccd1
+ _16096_/X sky130_fd_sc_hd__o221a_1
XFILLER_181_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19924_ _23592_/Q _19927_/C vssd1 vssd1 vccd1 vccd1 _19926_/A sky130_fd_sc_hd__and2_1
X_15047_ _15047_/A vssd1 vssd1 vccd1 vccd1 _22266_/D sky130_fd_sc_hd__clkbuf_1
X_12259_ _12252_/Y _12254_/Y _12256_/Y _12258_/Y _11242_/A vssd1 vssd1 vccd1 vccd1
+ _12260_/C sky130_fd_sc_hd__o221a_1
XFILLER_272_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19855_ _19855_/A vssd1 vssd1 vccd1 vccd1 _23561_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_268_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18806_ _23119_/Q _18804_/X _18818_/S vssd1 vssd1 vccd1 vccd1 _18807_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19786_ _19786_/A vssd1 vssd1 vccd1 vccd1 _23530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16998_ _17000_/A _16975_/X _16995_/X _16996_/X _16997_/X vssd1 vssd1 vccd1 vccd1
+ _16998_/X sky130_fd_sc_hd__o221a_2
XFILLER_49_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18737_ _16870_/X _23094_/Q _18741_/S vssd1 vssd1 vccd1 vccd1 _18738_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15949_ _15946_/Y _15948_/X _14690_/X vssd1 vssd1 vccd1 vccd1 _15949_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_237_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18668_ _18668_/A vssd1 vssd1 vccd1 vccd1 _23063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17619_ _17619_/A vssd1 vssd1 vccd1 vccd1 _22700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18599_ _18610_/A vssd1 vssd1 vccd1 vccd1 _18608_/S sky130_fd_sc_hd__buf_4
XFILLER_251_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_53_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23444_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20630_ _20630_/A vssd1 vssd1 vccd1 vccd1 _20631_/A sky130_fd_sc_hd__inv_2
XFILLER_211_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20561_ _20891_/A vssd1 vssd1 vccd1 vccd1 _21085_/A sky130_fd_sc_hd__buf_6
XFILLER_220_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22300_ _23144_/CLK _22300_/D vssd1 vssd1 vccd1 vccd1 _22300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_307_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23280_ _23409_/CLK _23280_/D vssd1 vssd1 vccd1 vccd1 _23280_/Q sky130_fd_sc_hd__dfxtp_1
X_20492_ _20765_/A _20428_/A _20491_/X _20483_/X vssd1 vssd1 vccd1 vccd1 _23716_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_354_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22231_ _22231_/A _22231_/B vssd1 vssd1 vccd1 vccd1 _22232_/B sky130_fd_sc_hd__xnor2_1
XFILLER_334_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22162_ _22177_/A _22162_/B vssd1 vssd1 vccd1 vccd1 _22163_/B sky130_fd_sc_hd__and2_1
XFILLER_279_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21113_ _21121_/A _21113_/B vssd1 vssd1 vccd1 vccd1 _23852_/D sky130_fd_sc_hd__nor2_1
XTAP_6907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22093_ _22093_/A _22093_/B vssd1 vssd1 vccd1 vccd1 _22093_/Y sky130_fd_sc_hd__nand2_1
XTAP_6929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21044_ _23832_/Q _20996_/B _21043_/Y _21037_/X vssd1 vssd1 vccd1 vccd1 _23832_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_286_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22995_ _23008_/CLK _22995_/D vssd1 vssd1 vccd1 vccd1 _22995_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_28_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_264_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21946_ _21911_/A _21913_/B _21910_/Y vssd1 vssd1 vccd1 vccd1 _21947_/B sky130_fd_sc_hd__o21ai_1
XFILLER_216_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21877_ _21877_/A vssd1 vssd1 vccd1 vccd1 _21877_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23616_ _23637_/CLK _23616_/D vssd1 vssd1 vccd1 vccd1 _23616_/Q sky130_fd_sc_hd__dfxtp_2
X_11630_ _11630_/A vssd1 vssd1 vccd1 vccd1 _11631_/A sky130_fd_sc_hd__buf_4
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20828_ _20864_/A vssd1 vssd1 vccd1 vccd1 _20828_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23547_ _23547_/CLK _23547_/D vssd1 vssd1 vccd1 vccd1 _23547_/Q sky130_fd_sc_hd__dfxtp_1
X_11561_ _11561_/A vssd1 vssd1 vccd1 vccd1 _12820_/S sky130_fd_sc_hd__buf_6
XFILLER_24_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_357_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_345_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20759_ _20759_/A _20759_/B vssd1 vssd1 vccd1 vccd1 _20762_/B sky130_fd_sc_hd__and2_1
XFILLER_156_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13300_ _13319_/A _13300_/B vssd1 vssd1 vccd1 vccd1 _16054_/A sky130_fd_sc_hd__and2_2
XFILLER_287_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14280_ _14272_/X _14278_/X _14639_/A vssd1 vssd1 vccd1 vccd1 _14280_/X sky130_fd_sc_hd__mux2_1
XFILLER_312_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23478_ _23510_/CLK _23478_/D vssd1 vssd1 vccd1 vccd1 _23478_/Q sky130_fd_sc_hd__dfxtp_4
X_11492_ _22322_/Q _23458_/Q _11492_/S vssd1 vssd1 vccd1 vccd1 _11492_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13231_ _13216_/A _13230_/X _12745_/A vssd1 vssd1 vccd1 vccd1 _13231_/X sky130_fd_sc_hd__o21a_1
X_22429_ _23500_/CLK _22429_/D vssd1 vssd1 vccd1 vccd1 _22429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13162_ _11219_/A _13152_/X _13161_/X _13210_/A vssd1 vssd1 vccd1 vccd1 _13163_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_237_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12113_ _15460_/A _12113_/B vssd1 vssd1 vccd1 vccd1 _13623_/A sky130_fd_sc_hd__nor2_4
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17970_ _22834_/Q _17965_/X _17969_/X _17963_/X vssd1 vssd1 vccd1 vccd1 _22834_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_340_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13093_ _11169_/A _13088_/X _13092_/X vssd1 vssd1 vccd1 vccd1 _13093_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_312_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_297_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_300_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12044_ _11584_/A _12043_/X _11961_/A vssd1 vssd1 vccd1 vccd1 _12044_/X sky130_fd_sc_hd__a21o_1
X_16921_ _17255_/A vssd1 vssd1 vccd1 vccd1 _17091_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_306_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19640_ _19697_/S vssd1 vssd1 vccd1 vccd1 _19649_/S sky130_fd_sc_hd__buf_4
X_16852_ _16851_/X _22532_/Q _16861_/S vssd1 vssd1 vccd1 vccd1 _16853_/A sky130_fd_sc_hd__mux2_1
XFILLER_266_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15803_ _22935_/Q _15903_/B vssd1 vssd1 vccd1 vccd1 _15803_/X sky130_fd_sc_hd__and2_1
X_16783_ _16783_/A vssd1 vssd1 vccd1 vccd1 _16783_/X sky130_fd_sc_hd__clkbuf_2
X_19571_ _23435_/Q _19185_/A _19577_/S vssd1 vssd1 vccd1 vccd1 _19572_/A sky130_fd_sc_hd__mux2_1
X_13995_ _14046_/A vssd1 vssd1 vccd1 vccd1 _14000_/A sky130_fd_sc_hd__buf_4
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18522_ _23003_/Q _18530_/B vssd1 vssd1 vccd1 vccd1 _18522_/Y sky130_fd_sc_hd__nand2_1
X_15734_ _14745_/A _15727_/X _15733_/Y _15652_/A vssd1 vssd1 vccd1 vccd1 _15735_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_12946_ _13006_/A _12946_/B vssd1 vssd1 vccd1 vccd1 _12946_/X sky130_fd_sc_hd__or2_1
XFILLER_34_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18453_ _18521_/A vssd1 vssd1 vccd1 vccd1 _18534_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_261_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15665_ _17172_/A _15617_/X _15662_/X _15664_/Y _15618_/X vssd1 vssd1 vccd1 vccd1
+ _15665_/X sky130_fd_sc_hd__o221a_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _12919_/A _12877_/B vssd1 vssd1 vccd1 vccd1 _12877_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_324_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14616_ _22947_/Q _14615_/X _15360_/A vssd1 vssd1 vccd1 vccd1 _14616_/X sky130_fd_sc_hd__mux2_1
X_17404_ _22615_/Q _16211_/X _17410_/S vssd1 vssd1 vccd1 vccd1 _17405_/A sky130_fd_sc_hd__mux2_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18384_ _22954_/Q _22955_/Q _18384_/C vssd1 vssd1 vccd1 vccd1 _18386_/B sky130_fd_sc_hd__and3_1
X_11828_ _23921_/Q _11828_/B vssd1 vssd1 vccd1 vccd1 _11828_/X sky130_fd_sc_hd__or2_1
XFILLER_221_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15596_ _15596_/A vssd1 vssd1 vccd1 vccd1 _15596_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17335_ _22590_/Q input207/X _17335_/S vssd1 vssd1 vccd1 vccd1 _17336_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14547_ _14546_/X _16936_/C _14557_/A vssd1 vssd1 vccd1 vccd1 _16203_/B sky130_fd_sc_hd__mux2_1
X_11759_ _12139_/A _11758_/X _11681_/A vssd1 vssd1 vccd1 vccd1 _11759_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_336_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_348_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_348_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_308_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17266_ input96/X input61/X _17266_/S vssd1 vssd1 vccd1 vccd1 _17266_/X sky130_fd_sc_hd__mux2_8
XFILLER_347_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14478_ _15216_/A vssd1 vssd1 vccd1 vccd1 _14478_/X sky130_fd_sc_hd__buf_2
XFILLER_335_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19005_ _19005_/A vssd1 vssd1 vccd1 vccd1 _23198_/D sky130_fd_sc_hd__clkbuf_1
X_16217_ _18782_/A vssd1 vssd1 vccd1 vccd1 _16217_/X sky130_fd_sc_hd__buf_2
X_13429_ _14815_/B _13410_/Y _13415_/X _13428_/X vssd1 vssd1 vccd1 vccd1 _21518_/A
+ sky130_fd_sc_hd__a211o_2
X_17197_ _17167_/X _17191_/X _17196_/X _17176_/X vssd1 vssd1 vccd1 vccd1 _17197_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_289_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16148_ _15676_/X _21280_/A _16147_/X _15365_/X vssd1 vssd1 vccd1 vccd1 _16148_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_127_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_288_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_171_wb_clk_i _23917_/CLK vssd1 vssd1 vccd1 vccd1 _22520_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_331_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_288_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_331_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_100_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23552_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16079_ _16079_/A _16079_/B vssd1 vssd1 vccd1 vccd1 _16079_/X sky130_fd_sc_hd__or2_1
XFILLER_143_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19907_ _16297_/X _23585_/Q _19909_/S vssd1 vssd1 vccd1 vccd1 _19908_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19838_ _19838_/A vssd1 vssd1 vccd1 vccd1 _23554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_256_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput1 coreIndex[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_4
XFILLER_256_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19769_ _19264_/X _23524_/Q _19769_/S vssd1 vssd1 vccd1 vccd1 _19770_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21800_ _21801_/C _21798_/X _21801_/D _21799_/Y _21778_/B vssd1 vssd1 vccd1 vccd1
+ _21800_/X sky130_fd_sc_hd__a311o_1
XFILLER_37_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22780_ _23048_/CLK _22780_/D vssd1 vssd1 vccd1 vccd1 _22780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21731_ _23826_/Q _23760_/Q vssd1 vssd1 vccd1 vccd1 _21733_/A sky130_fd_sc_hd__and2_1
XFILLER_101_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21662_ _23792_/Q _21814_/B vssd1 vssd1 vccd1 vccd1 _21662_/Y sky130_fd_sc_hd__nand2_2
XFILLER_339_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23401_ _23558_/CLK _23401_/D vssd1 vssd1 vccd1 vccd1 _23401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_339_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20613_ _20626_/A _20613_/B _20613_/C vssd1 vssd1 vccd1 vccd1 _20613_/X sky130_fd_sc_hd__or3_1
XFILLER_177_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21593_ _21593_/A _21593_/B vssd1 vssd1 vccd1 vccd1 _21593_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_338_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23332_ _23556_/CLK _23332_/D vssd1 vssd1 vccd1 vccd1 _23332_/Q sky130_fd_sc_hd__dfxtp_1
X_20544_ _20544_/A vssd1 vssd1 vccd1 vccd1 _20774_/A sky130_fd_sc_hd__buf_4
XFILLER_326_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_338_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_354_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23263_ _23423_/CLK _23263_/D vssd1 vssd1 vccd1 vccd1 _23263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20475_ _23708_/Q _20416_/B _20474_/Y _20472_/X vssd1 vssd1 vccd1 vccd1 _23708_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_307_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22214_ _23843_/Q _22213_/Y _22214_/S vssd1 vssd1 vccd1 vccd1 _22215_/B sky130_fd_sc_hd__mux2_1
XFILLER_307_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23194_ _23354_/CLK _23194_/D vssd1 vssd1 vccd1 vccd1 _23194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_279_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22145_ _21594_/B _22142_/X _22143_/Y _22144_/X vssd1 vssd1 vccd1 vccd1 _22146_/C
+ sky130_fd_sc_hd__a31oi_4
XFILLER_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_295_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput360 _13726_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[6] sky130_fd_sc_hd__buf_2
XTAP_6726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput371 _13678_/X vssd1 vssd1 vccd1 vccd1 csb0[1] sky130_fd_sc_hd__buf_2
XTAP_6737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput382 _14044_/X vssd1 vssd1 vccd1 vccd1 din0[17] sky130_fd_sc_hd__buf_2
XFILLER_117_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_294_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_288_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22076_ _22076_/A _22155_/B vssd1 vssd1 vccd1 vccd1 _22076_/Y sky130_fd_sc_hd__xnor2_1
Xoutput393 _14063_/X vssd1 vssd1 vccd1 vccd1 din0[27] sky130_fd_sc_hd__buf_2
XTAP_6759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21027_ _21047_/A vssd1 vssd1 vccd1 vccd1 _21027_/X sky130_fd_sc_hd__buf_2
XFILLER_259_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12800_ _13295_/A _12800_/B _12800_/C vssd1 vssd1 vccd1 vccd1 _12800_/Y sky130_fd_sc_hd__nor3_4
XFILLER_28_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13780_ _13808_/A vssd1 vssd1 vccd1 vccd1 _13836_/B sky130_fd_sc_hd__clkbuf_2
X_22978_ _23424_/CLK _22978_/D vssd1 vssd1 vccd1 vccd1 _22978_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_83_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12731_ _22796_/Q _22764_/Q _22665_/Q _22732_/Q _12716_/X _12717_/X vssd1 vssd1 vccd1
+ vccd1 _12732_/B sky130_fd_sc_hd__mux4_1
XFILLER_243_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_308_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21929_ _21987_/A _22041_/A vssd1 vssd1 vccd1 vccd1 _21932_/A sky130_fd_sc_hd__and2_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ _15982_/B _15450_/B vssd1 vssd1 vccd1 vccd1 _15450_/Y sky130_fd_sc_hd__nand2_1
XFILLER_204_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12662_ _11323_/A _12913_/S _11401_/A _12661_/Y vssd1 vssd1 vccd1 vccd1 _12664_/A
+ sky130_fd_sc_hd__a2bb2o_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14401_ _15864_/A _22249_/D _14421_/S vssd1 vssd1 vccd1 vccd1 _14457_/A sky130_fd_sc_hd__mux2_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11613_/A vssd1 vssd1 vccd1 vccd1 _11613_/X sky130_fd_sc_hd__buf_6
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_358_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15381_ _15381_/A _15485_/B vssd1 vssd1 vccd1 vccd1 _15381_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12593_ _12586_/X _12588_/X _12590_/X _12592_/X _11273_/A vssd1 vssd1 vccd1 vccd1
+ _12594_/C sky130_fd_sc_hd__a221o_1
XFILLER_156_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_358_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17120_ _22565_/Q _17091_/X _17083_/X _17119_/X vssd1 vssd1 vccd1 vccd1 _22565_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_357_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14332_ _14328_/X _14331_/X _14639_/A vssd1 vssd1 vccd1 vccd1 _14333_/A sky130_fd_sc_hd__mux2_1
X_11544_ _11544_/A vssd1 vssd1 vccd1 vccd1 _13276_/A sky130_fd_sc_hd__buf_4
XFILLER_344_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_317_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_344_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17051_ input74/X input103/X _17084_/S vssd1 vssd1 vccd1 vccd1 _17051_/X sky130_fd_sc_hd__mux2_8
XFILLER_144_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14263_ _15798_/A vssd1 vssd1 vccd1 vccd1 _16097_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_184_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11475_ _23235_/Q _23203_/Q _23171_/Q _23139_/Q _21771_/A _15616_/A vssd1 vssd1 vccd1
+ vccd1 _11476_/B sky130_fd_sc_hd__mux4_1
XFILLER_183_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16002_ _15676_/X _21272_/A _16001_/X _15365_/X vssd1 vssd1 vccd1 vccd1 _16002_/X
+ sky130_fd_sc_hd__o22a_1
X_13214_ _23935_/Q vssd1 vssd1 vccd1 vccd1 _13214_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_344_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_298_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14194_ _14820_/A _15440_/A _15672_/A _14199_/B _14193_/Y vssd1 vssd1 vccd1 vccd1
+ _14202_/C sky130_fd_sc_hd__a41o_1
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_341_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13145_ _22479_/Q _22639_/Q _13191_/S vssd1 vssd1 vccd1 vccd1 _13145_/X sky130_fd_sc_hd__mux2_1
XFILLER_298_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_298_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _22828_/Q _17950_/X _17952_/X _17948_/X vssd1 vssd1 vccd1 vccd1 _22828_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_340_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13076_ _13069_/Y _13071_/Y _13073_/Y _13075_/Y _11483_/A vssd1 vssd1 vccd1 vccd1
+ _13076_/X sky130_fd_sc_hd__o221a_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_300_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16904_ _16904_/A vssd1 vssd1 vccd1 vccd1 _22548_/D sky130_fd_sc_hd__clkbuf_1
X_12027_ _12998_/A _12027_/B vssd1 vssd1 vccd1 vccd1 _12027_/Y sky130_fd_sc_hd__nor2_1
XFILLER_250_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17884_ _22891_/Q _22890_/Q vssd1 vssd1 vccd1 vccd1 _18142_/A sky130_fd_sc_hd__nand2_2
XFILLER_120_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19623_ _23459_/Q _19261_/A _19625_/S vssd1 vssd1 vccd1 vccd1 _19624_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_333_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16835_ _19185_/A vssd1 vssd1 vccd1 vccd1 _16835_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19554_ _19554_/A vssd1 vssd1 vccd1 vccd1 _23428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16766_ _16784_/A vssd1 vssd1 vccd1 vccd1 _16766_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13978_ _13978_/A vssd1 vssd1 vccd1 vccd1 _13978_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_206_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18505_ _22997_/Q _18505_/B vssd1 vssd1 vccd1 vccd1 _18505_/Y sky130_fd_sc_hd__nand2_1
XFILLER_222_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12929_ _11233_/A _12919_/Y _12924_/Y _12926_/Y _12928_/Y vssd1 vssd1 vccd1 vccd1
+ _12929_/X sky130_fd_sc_hd__o32a_1
XFILLER_202_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15717_ _14833_/A _15331_/Y _15578_/A vssd1 vssd1 vccd1 vccd1 _15717_/X sky130_fd_sc_hd__a21bo_2
XFILLER_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16697_ _22488_/Q _16689_/X _16693_/X input21/X vssd1 vssd1 vccd1 vccd1 _16698_/B
+ sky130_fd_sc_hd__o22a_1
X_19485_ _19553_/S vssd1 vssd1 vccd1 vccd1 _19494_/S sky130_fd_sc_hd__buf_6
XFILLER_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18436_ _19923_/A _18436_/B _18440_/C vssd1 vssd1 vccd1 vccd1 _22973_/D sky130_fd_sc_hd__nor3_1
X_15648_ _23798_/Q _14917_/X _14919_/X vssd1 vssd1 vccd1 vccd1 _15648_/X sky130_fd_sc_hd__a21o_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18367_ _18401_/A _18367_/B _18369_/B vssd1 vssd1 vccd1 vccd1 _22949_/D sky130_fd_sc_hd__nor3_1
XFILLER_175_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15579_ _15575_/X _15186_/Y _15674_/A vssd1 vssd1 vccd1 vccd1 _15579_/X sky130_fd_sc_hd__a21bo_2
XFILLER_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_336_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17318_ _17315_/X _17317_/X _17318_/S vssd1 vssd1 vccd1 vccd1 _17318_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18298_ _22924_/Q _22925_/Q _22926_/Q _18298_/D vssd1 vssd1 vccd1 vccd1 _18307_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_174_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_336_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17249_ _15929_/X _17247_/X _17291_/S vssd1 vssd1 vccd1 vccd1 _17249_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_317_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20260_ _20213_/X _20639_/A _20259_/X _20246_/X vssd1 vssd1 vccd1 vccd1 _23664_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_350_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20191_ _20191_/A vssd1 vssd1 vccd1 vccd1 _20307_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_304_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23950_ _23950_/A vssd1 vssd1 vccd1 vccd1 _23950_/X sky130_fd_sc_hd__buf_2
XFILLER_97_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_257_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22901_ _22908_/CLK _22901_/D vssd1 vssd1 vccd1 vccd1 _22901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23881_ _23888_/CLK _23881_/D vssd1 vssd1 vccd1 vccd1 _23881_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22832_ _22893_/CLK _22832_/D vssd1 vssd1 vccd1 vccd1 _22832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22763_ _23575_/CLK _22763_/D vssd1 vssd1 vccd1 vccd1 _22763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21714_ _21714_/A _21714_/B vssd1 vssd1 vccd1 vccd1 _21714_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22694_ _23414_/CLK _22694_/D vssd1 vssd1 vccd1 vccd1 _22694_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21645_ _13951_/B _21612_/X _21644_/X _21581_/X vssd1 vssd1 vccd1 vccd1 _23921_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_339_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21576_ _21576_/A _22032_/B vssd1 vssd1 vccd1 vccd1 _21576_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23315_ _23510_/CLK _23315_/D vssd1 vssd1 vccd1 vccd1 _23315_/Q sky130_fd_sc_hd__dfxtp_1
X_20527_ _20531_/A _20531_/B vssd1 vssd1 vccd1 vccd1 _21357_/C sky130_fd_sc_hd__or2_4
XFILLER_355_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_308_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11260_ _23907_/Q _23906_/Q _23905_/Q _23904_/Q vssd1 vssd1 vccd1 vccd1 _14180_/D
+ sky130_fd_sc_hd__or4_2
X_23246_ _23534_/CLK _23246_/D vssd1 vssd1 vccd1 vccd1 _23246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20458_ _20963_/A vssd1 vssd1 vccd1 vccd1 _20602_/A sky130_fd_sc_hd__buf_6
XTAP_7202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_307_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_341_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_323_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11191_ _12423_/A vssd1 vssd1 vccd1 vccd1 _11837_/A sky130_fd_sc_hd__buf_4
X_23177_ _23561_/CLK _23177_/D vssd1 vssd1 vccd1 vccd1 _23177_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_7246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20389_ _20396_/A _20389_/B vssd1 vssd1 vccd1 vccd1 _20389_/X sky130_fd_sc_hd__or2_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22128_ _22128_/A _22155_/D vssd1 vssd1 vccd1 vccd1 _22128_/Y sky130_fd_sc_hd__xnor2_2
XTAP_7279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14950_ _14858_/X _14949_/X _15084_/S vssd1 vssd1 vccd1 vccd1 _14951_/A sky130_fd_sc_hd__mux2_1
X_22059_ _22059_/A _22059_/B vssd1 vssd1 vccd1 vccd1 _22059_/Y sky130_fd_sc_hd__xnor2_1
XTAP_6589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13901_ _13901_/A vssd1 vssd1 vccd1 vccd1 _17020_/A sky130_fd_sc_hd__buf_6
XFILLER_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14881_ _15698_/A vssd1 vssd1 vccd1 vccd1 _14882_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13832_ _13832_/A vssd1 vssd1 vccd1 vccd1 _13833_/A sky130_fd_sc_hd__clkbuf_2
X_16620_ _16677_/S vssd1 vssd1 vccd1 vccd1 _16629_/S sky130_fd_sc_hd__buf_4
XFILLER_29_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_207 _21526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16551_ _15104_/X _22428_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _16552_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_218 _14879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13763_ _13763_/A _14207_/A vssd1 vssd1 vccd1 vccd1 _14074_/A sky130_fd_sc_hd__or2_1
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_229 _15110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ _23480_/Q _23576_/Q _22540_/Q _22344_/Q _12709_/X _12710_/X vssd1 vssd1 vccd1
+ vccd1 _12715_/B sky130_fd_sc_hd__mux4_1
X_15502_ _15735_/A vssd1 vssd1 vccd1 vccd1 _16144_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_71_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16482_ _16528_/S vssd1 vssd1 vccd1 vccd1 _16491_/S sky130_fd_sc_hd__buf_4
X_19270_ _19163_/X _23301_/Q _19278_/S vssd1 vssd1 vccd1 vccd1 _19271_/A sky130_fd_sc_hd__mux2_1
X_13694_ _13969_/A vssd1 vssd1 vccd1 vccd1 _13985_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_18221_ _22900_/Q _18227_/B vssd1 vssd1 vccd1 vccd1 _18221_/X sky130_fd_sc_hd__or2_1
X_15433_ _15433_/A _15433_/B vssd1 vssd1 vccd1 vccd1 _15433_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12645_ _12698_/A _12645_/B vssd1 vssd1 vccd1 vccd1 _12645_/Y sky130_fd_sc_hd__nor2_1
XPHY_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18152_ _14119_/C _22880_/Q _18158_/S vssd1 vssd1 vccd1 vccd1 _18153_/B sky130_fd_sc_hd__mux2_1
XFILLER_169_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15364_ _15336_/X _15345_/Y _15363_/Y vssd1 vssd1 vccd1 vccd1 _15364_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_156_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12576_ _22265_/Q _23081_/Q _23497_/Q _22426_/Q _11799_/A _12329_/X vssd1 vssd1 vccd1
+ vccd1 _12577_/B sky130_fd_sc_hd__mux4_1
XFILLER_357_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17103_ _17103_/A vssd1 vssd1 vccd1 vccd1 _17103_/Y sky130_fd_sc_hd__inv_2
X_14315_ _15130_/S vssd1 vssd1 vccd1 vccd1 _15084_/S sky130_fd_sc_hd__buf_2
X_18083_ _18098_/A vssd1 vssd1 vccd1 vccd1 _18083_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11527_ _11527_/A vssd1 vssd1 vccd1 vccd1 _11527_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15295_ _11940_/A _15582_/B _14674_/X _13948_/A _15769_/A vssd1 vssd1 vccd1 vccd1
+ _15295_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_117_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_328_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17034_ _17033_/B _17032_/X _17033_/Y _16951_/X vssd1 vssd1 vccd1 vccd1 _17034_/X
+ sky130_fd_sc_hd__o211a_1
X_14246_ _14246_/A _14246_/B vssd1 vssd1 vccd1 vccd1 _14247_/A sky130_fd_sc_hd__or2_2
XFILLER_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11458_ _12414_/A vssd1 vssd1 vccd1 vccd1 _12634_/A sky130_fd_sc_hd__buf_8
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_314_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_4_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_14177_ _14177_/A _15455_/A vssd1 vssd1 vccd1 vccd1 _14177_/Y sky130_fd_sc_hd__nand2_1
X_11389_ _13234_/S vssd1 vssd1 vccd1 vccd1 _13185_/S sky130_fd_sc_hd__buf_6
XFILLER_98_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_301_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13128_ _22383_/Q _22415_/Q _22704_/Q _23071_/Q _11543_/A _13127_/X vssd1 vssd1 vccd1
+ vccd1 _13128_/X sky130_fd_sc_hd__mux4_2
XFILLER_258_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18985_ _18985_/A vssd1 vssd1 vccd1 vccd1 _23189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17936_ _22823_/Q _17922_/X _17918_/X input254/X _17933_/X vssd1 vssd1 vccd1 vccd1
+ _17936_/X sky130_fd_sc_hd__a221o_1
XFILLER_285_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13059_ _22288_/Q _23104_/Q _23520_/Q _22449_/Q _13275_/A _11527_/X vssd1 vssd1 vccd1
+ vccd1 _13060_/B sky130_fd_sc_hd__mux4_1
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17867_ _17867_/A vssd1 vssd1 vccd1 vccd1 _22804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19606_ _23451_/Q _19236_/A _19610_/S vssd1 vssd1 vccd1 vccd1 _19607_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16818_ _16818_/A vssd1 vssd1 vccd1 vccd1 _22521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_282_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17798_ _22774_/Q _17639_/X _17798_/S vssd1 vssd1 vccd1 vccd1 _17799_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19537_ _19537_/A vssd1 vssd1 vccd1 vccd1 _23420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16749_ _22502_/Q _16747_/X _16748_/X input16/X vssd1 vssd1 vccd1 vccd1 _16750_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_235_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19468_ _19468_/A vssd1 vssd1 vccd1 vccd1 _19477_/S sky130_fd_sc_hd__buf_4
XFILLER_35_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18419_ _19923_/A _18419_/B _18420_/B vssd1 vssd1 vccd1 vccd1 _22967_/D sky130_fd_sc_hd__nor3_1
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19399_ _23359_/Q _18856_/X _19405_/S vssd1 vssd1 vccd1 vccd1 _19400_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21430_ _23785_/Q _21381_/X _21428_/Y _21813_/A vssd1 vssd1 vccd1 vccd1 _21430_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_296_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_337_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21361_ _21361_/A _21361_/B _21361_/C vssd1 vssd1 vccd1 vccd1 _21361_/X sky130_fd_sc_hd__or3_2
XFILLER_296_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_352_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_308_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23100_ _23100_/CLK _23100_/D vssd1 vssd1 vccd1 vccd1 _23100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20312_ _17182_/A _20295_/X _20313_/B vssd1 vssd1 vccd1 vccd1 _20312_/X sky130_fd_sc_hd__o21a_1
Xinput70 dout0[34] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_1
XFILLER_317_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21292_ _17244_/B _21290_/X _21291_/X _14160_/X vssd1 vssd1 vccd1 vccd1 _21320_/B
+ sky130_fd_sc_hd__a22o_4
Xinput81 dout0[44] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__clkbuf_1
XFILLER_305_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput92 dout0[54] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__clkbuf_1
X_23031_ _23511_/CLK _23031_/D vssd1 vssd1 vccd1 vccd1 _23031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20243_ _20250_/A _20243_/B vssd1 vssd1 vccd1 vccd1 _20243_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20174_ _20174_/A vssd1 vssd1 vccd1 vccd1 _20174_/X sky130_fd_sc_hd__buf_2
XFILLER_130_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23933_ _23934_/CLK _23933_/D vssd1 vssd1 vccd1 vccd1 _23933_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23864_ _23871_/CLK _23864_/D vssd1 vssd1 vccd1 vccd1 _23864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23054_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22815_ _22830_/CLK _22815_/D vssd1 vssd1 vccd1 vccd1 _22815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_351_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23795_ _23861_/CLK _23795_/D vssd1 vssd1 vccd1 vccd1 _23795_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22746_ _23496_/CLK _22746_/D vssd1 vssd1 vccd1 vccd1 _22746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_349_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22677_ _23588_/CLK _22677_/D vssd1 vssd1 vccd1 vccd1 _22677_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_203_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23564_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_240_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12430_ _23303_/Q _23271_/Q _23239_/Q _23527_/Q _11699_/A _11840_/A vssd1 vssd1 vccd1
+ vccd1 _12431_/B sky130_fd_sc_hd__mux4_1
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21628_ _23823_/Q _23757_/Q vssd1 vssd1 vccd1 vccd1 _21629_/B sky130_fd_sc_hd__nand2_1
XFILLER_327_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12361_ _12196_/A _12360_/X _11780_/A vssd1 vssd1 vccd1 vccd1 _12361_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_139_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21559_ _21559_/A _21559_/B vssd1 vssd1 vccd1 vccd1 _21559_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_126_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_355_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_327_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_343_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14100_ _22597_/Q _14081_/A _14099_/Y _14012_/X vssd1 vssd1 vccd1 vccd1 _14100_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_295_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11312_ _11364_/A vssd1 vssd1 vccd1 vccd1 _11468_/A sky130_fd_sc_hd__clkbuf_4
X_15080_ _15080_/A vssd1 vssd1 vccd1 vccd1 _15081_/A sky130_fd_sc_hd__buf_6
XFILLER_4_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12292_ _12292_/A vssd1 vssd1 vccd1 vccd1 _12292_/X sky130_fd_sc_hd__buf_4
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14031_ _14069_/B vssd1 vssd1 vccd1 vccd1 _14052_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_342_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23229_ _23547_/CLK _23229_/D vssd1 vssd1 vccd1 vccd1 _23229_/Q sky130_fd_sc_hd__dfxtp_1
X_11243_ _11243_/A vssd1 vssd1 vccd1 vccd1 _11244_/A sky130_fd_sc_hd__clkbuf_8
XTAP_7021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11174_ _11603_/A vssd1 vssd1 vccd1 vccd1 _12532_/A sky130_fd_sc_hd__buf_2
XFILLER_122_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_311_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18770_ _18770_/A _18770_/B _17471_/A vssd1 vssd1 vccd1 vccd1 _19018_/B sky130_fd_sc_hd__or3b_4
XFILLER_310_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15982_ _22972_/Q _15982_/B vssd1 vssd1 vccd1 vccd1 _15982_/X sky130_fd_sc_hd__or2_1
XFILLER_121_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17721_ _17721_/A vssd1 vssd1 vccd1 vccd1 _22739_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_314_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14933_ _14933_/A vssd1 vssd1 vccd1 vccd1 _15001_/A sky130_fd_sc_hd__buf_2
XFILLER_94_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ input226/X _16085_/X _14700_/X vssd1 vssd1 vccd1 vccd1 _17653_/A sky130_fd_sc_hd__a21oi_4
XFILLER_180_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_291_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14864_ _15335_/B vssd1 vssd1 vccd1 vccd1 _14940_/B sky130_fd_sc_hd__clkbuf_2
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16603_ _16161_/X _22452_/Q _16605_/S vssd1 vssd1 vccd1 vccd1 _16604_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13815_ _14241_/A _13815_/B vssd1 vssd1 vccd1 vccd1 _13863_/A sky130_fd_sc_hd__and2_1
X_17583_ _22689_/Q _17582_/X _17592_/S vssd1 vssd1 vccd1 vccd1 _17584_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14795_ _20532_/A vssd1 vssd1 vccd1 vccd1 _15636_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19322_ _19242_/X _23325_/Q _19322_/S vssd1 vssd1 vccd1 vccd1 _19323_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16534_ _20134_/A _16534_/B vssd1 vssd1 vccd1 vccd1 _22421_/D sky130_fd_sc_hd__nor2_1
X_13746_ _13781_/A vssd1 vssd1 vccd1 vccd1 _13746_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19253_ _19252_/X _23296_/Q _19259_/S vssd1 vssd1 vccd1 vccd1 _19254_/A sky130_fd_sc_hd__mux2_1
X_16465_ _14811_/X _22391_/Q _16469_/S vssd1 vssd1 vccd1 vccd1 _16466_/A sky130_fd_sc_hd__mux2_1
X_13677_ _17029_/S _13679_/B vssd1 vssd1 vccd1 vccd1 _13678_/A sky130_fd_sc_hd__or2b_1
X_18204_ _18243_/A vssd1 vssd1 vccd1 vccd1 _18214_/B sky130_fd_sc_hd__clkbuf_1
X_12628_ _12708_/A _12627_/X _11285_/A vssd1 vssd1 vccd1 vccd1 _12628_/Y sky130_fd_sc_hd__o21ai_1
XPHY_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15416_ _15416_/A vssd1 vssd1 vccd1 vccd1 _15620_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_129_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19184_ _19184_/A vssd1 vssd1 vccd1 vccd1 _23274_/D sky130_fd_sc_hd__clkbuf_1
X_16396_ _14984_/X _22361_/Q _16396_/S vssd1 vssd1 vccd1 vccd1 _16397_/A sky130_fd_sc_hd__mux2_1
XFILLER_318_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18135_ _21681_/A vssd1 vssd1 vccd1 vccd1 _18135_/X sky130_fd_sc_hd__buf_12
X_15347_ _15832_/A vssd1 vssd1 vccd1 vccd1 _15697_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_129_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12559_ _23209_/Q _23177_/Q _23145_/Q _23113_/Q _12242_/S _11611_/A vssd1 vssd1 vccd1
+ vccd1 _12559_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_333_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18066_ _18096_/A vssd1 vssd1 vccd1 vccd1 _18066_/X sky130_fd_sc_hd__clkbuf_2
X_15278_ _15161_/A _15273_/X _15277_/Y _15162_/X vssd1 vssd1 vccd1 vccd1 _15278_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17017_ _17145_/B vssd1 vssd1 vccd1 vccd1 _17017_/X sky130_fd_sc_hd__clkbuf_2
X_14229_ _22511_/Q _14219_/X _14223_/X _14228_/X vssd1 vssd1 vccd1 vccd1 _14230_/B
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_78_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23550_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_217_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_320_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_302_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_291_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18968_ _16844_/X _23182_/Q _18968_/S vssd1 vssd1 vccd1 vccd1 _18969_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_286_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17919_ _22818_/Q _17894_/X _17918_/X input259/X _17915_/X vssd1 vssd1 vccd1 vccd1
+ _17919_/X sky130_fd_sc_hd__a221o_1
X_18899_ _23151_/Q _18804_/X _18907_/S vssd1 vssd1 vccd1 vccd1 _18900_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20930_ _23792_/Q _20925_/X _20929_/X _20920_/X vssd1 vssd1 vccd1 vccd1 _23792_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_226_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20861_ _20861_/A _20861_/B vssd1 vssd1 vccd1 vccd1 _20862_/A sky130_fd_sc_hd__and2_1
XFILLER_240_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22600_ _22600_/CLK _22600_/D vssd1 vssd1 vccd1 vccd1 _22600_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_207_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23580_ _23580_/CLK _23580_/D vssd1 vssd1 vccd1 vccd1 _23580_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20792_ _20811_/A vssd1 vssd1 vccd1 vccd1 _20792_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_560 _23881_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22531_ _23535_/CLK _22531_/D vssd1 vssd1 vccd1 vccd1 _22531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22462_ _23559_/CLK _22462_/D vssd1 vssd1 vccd1 vccd1 _22462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21413_ _21373_/A _21373_/B _21372_/A vssd1 vssd1 vccd1 vccd1 _21417_/A sky130_fd_sc_hd__o21a_1
XFILLER_185_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_336_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_309_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22393_ _22779_/CLK _22393_/D vssd1 vssd1 vccd1 vccd1 _22393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_337_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21344_ _21344_/A _21344_/B vssd1 vssd1 vccd1 vccd1 _21345_/B sky130_fd_sc_hd__nor2_1
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_324_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21275_ _21077_/A _21242_/X _21274_/Y _21270_/X vssd1 vssd1 vccd1 vccd1 _23906_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_296_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_305_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23014_ _23526_/CLK _23014_/D vssd1 vssd1 vccd1 vccd1 _23014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20226_ _20307_/A vssd1 vssd1 vccd1 vccd1 _20226_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20157_ _20236_/A _20152_/X _20155_/Y _20174_/A vssd1 vssd1 vccd1 vccd1 _20157_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_311_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20088_ _20134_/A _20088_/B vssd1 vssd1 vccd1 vccd1 _23637_/D sky130_fd_sc_hd__nor2_1
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11930_ _23405_/Q _23021_/Q _23373_/Q _23341_/Q _11814_/X _11800_/A vssd1 vssd1 vccd1
+ vccd1 _11931_/B sky130_fd_sc_hd__mux4_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23916_ _23916_/CLK _23916_/D vssd1 vssd1 vccd1 vccd1 _23916_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23847_ _23851_/CLK _23847_/D vssd1 vssd1 vccd1 vccd1 _23847_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _11926_/A _11861_/B vssd1 vssd1 vccd1 vccd1 _11861_/Y sky130_fd_sc_hd__nor2_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _20533_/C _13599_/X _13884_/A _23930_/Q vssd1 vssd1 vccd1 vccd1 _13970_/A
+ sky130_fd_sc_hd__a2bb2o_2
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14580_ _22496_/Q _14219_/X _14238_/X _14579_/X _14242_/X vssd1 vssd1 vccd1 vccd1
+ _14580_/Y sky130_fd_sc_hd__o221ai_4
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _11785_/Y _11787_/Y _11789_/Y _11791_/Y _11244_/A vssd1 vssd1 vccd1 vccd1
+ _11793_/C sky130_fd_sc_hd__o221a_1
X_23778_ _23810_/CLK _23778_/D vssd1 vssd1 vccd1 vccd1 _23778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13531_ _13531_/A _15492_/S vssd1 vssd1 vccd1 vccd1 _13531_/X sky130_fd_sc_hd__or2_1
X_22729_ _23573_/CLK _22729_/D vssd1 vssd1 vccd1 vccd1 _22729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_347_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_300_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16250_ _22306_/Q _16249_/X _16253_/S vssd1 vssd1 vccd1 vccd1 _16251_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13462_ _13471_/A _23945_/Q vssd1 vssd1 vccd1 vccd1 _13474_/A sky130_fd_sc_hd__nor2_2
XFILLER_40_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15201_ _15495_/A vssd1 vssd1 vccd1 vccd1 _15580_/B sky130_fd_sc_hd__buf_4
X_12413_ _12406_/Y _12408_/Y _12410_/Y _12412_/Y _11826_/A vssd1 vssd1 vccd1 vccd1
+ _12414_/C sky130_fd_sc_hd__o221a_1
X_16181_ _13410_/A _16180_/B _16180_/Y _15636_/A vssd1 vssd1 vccd1 vccd1 _16186_/B
+ sky130_fd_sc_hd__a211o_1
X_13393_ _13646_/A _13393_/B vssd1 vssd1 vccd1 vccd1 _13393_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_316_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_327_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_309_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15132_ _14846_/X _14850_/X _15132_/S vssd1 vssd1 vccd1 vccd1 _15132_/X sky130_fd_sc_hd__mux2_2
XFILLER_5_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12344_ _13472_/B _14385_/A vssd1 vssd1 vccd1 vccd1 _12344_/X sky130_fd_sc_hd__or2_4
XFILLER_154_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_343_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19940_ _19978_/C vssd1 vssd1 vccd1 vccd1 _19971_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15063_ _14970_/S _15053_/X _15062_/Y vssd1 vssd1 vccd1 vccd1 _21217_/A sky130_fd_sc_hd__o21ai_4
XFILLER_153_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12275_ _22363_/Q _22395_/Q _22684_/Q _23051_/Q _11647_/A _12269_/X vssd1 vssd1 vccd1
+ vccd1 _12275_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_299_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14014_ _14012_/X _13712_/B _14013_/X input237/X vssd1 vssd1 vccd1 vccd1 _14014_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_330_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11226_ _23492_/Q _23588_/Q _22552_/Q _22356_/Q _13434_/A _11170_/X vssd1 vssd1 vccd1
+ vccd1 _11226_/X sky130_fd_sc_hd__mux4_1
X_19871_ _19871_/A vssd1 vssd1 vccd1 vccd1 _23568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_295_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18822_ _23124_/Q _18820_/X _18834_/S vssd1 vssd1 vccd1 vccd1 _18823_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11157_ _11493_/S vssd1 vssd1 vccd1 vccd1 _11157_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_310_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18753_ _18753_/A vssd1 vssd1 vccd1 vccd1 _23101_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_310_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15965_ _15949_/Y _15964_/Y _16188_/A vssd1 vssd1 vccd1 vccd1 _15965_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11088_ _11095_/B vssd1 vssd1 vccd1 vccd1 _20148_/A sky130_fd_sc_hd__clkbuf_4
Xinput260 manufacturerID[6] vssd1 vssd1 vccd1 vccd1 input260/X sky130_fd_sc_hd__buf_2
XTAP_5471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput271 partID[1] vssd1 vssd1 vccd1 vccd1 input271/X sky130_fd_sc_hd__clkbuf_1
XFILLER_264_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17704_ _22732_/Q _17607_/X _17704_/S vssd1 vssd1 vccd1 vccd1 _17705_/A sky130_fd_sc_hd__mux2_1
XFILLER_209_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput282 versionID[2] vssd1 vssd1 vccd1 vccd1 input282/X sky130_fd_sc_hd__clkbuf_2
XTAP_5493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14916_ _14916_/A vssd1 vssd1 vccd1 vccd1 _14917_/A sky130_fd_sc_hd__clkbuf_4
X_18684_ _18684_/A vssd1 vssd1 vccd1 vccd1 _23070_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_286_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_196_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23529_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15896_ _15894_/X _22032_/A _16047_/S vssd1 vssd1 vccd1 vccd1 _18846_/A sky130_fd_sc_hd__mux2_8
XFILLER_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17635_ _17635_/A vssd1 vssd1 vccd1 vccd1 _22705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_125_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23646_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14847_ _14845_/X _14846_/X _14852_/S vssd1 vssd1 vccd1 vccd1 _14847_/X sky130_fd_sc_hd__mux2_2
XFILLER_291_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_327_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17566_ _18792_/A vssd1 vssd1 vccd1 vccd1 _17566_/X sky130_fd_sc_hd__clkbuf_2
X_14778_ _14778_/A _15085_/S vssd1 vssd1 vccd1 vccd1 _14778_/X sky130_fd_sc_hd__or2b_1
XFILLER_16_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19305_ _19217_/X _23317_/Q _19311_/S vssd1 vssd1 vccd1 vccd1 _19306_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16517_ _16517_/A vssd1 vssd1 vccd1 vccd1 _22414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13729_ _13729_/A vssd1 vssd1 vccd1 vccd1 _13729_/X sky130_fd_sc_hd__clkbuf_1
X_17497_ _22656_/Q _16239_/X _17505_/S vssd1 vssd1 vccd1 vccd1 _17498_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19236_ _19236_/A vssd1 vssd1 vccd1 vccd1 _19236_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_338_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16448_ _16448_/A vssd1 vssd1 vccd1 vccd1 _22384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19167_ _19163_/X _23269_/Q _19179_/S vssd1 vssd1 vccd1 vccd1 _19168_/A sky130_fd_sc_hd__mux2_1
XFILLER_318_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16379_ _16161_/X _22355_/Q _16381_/S vssd1 vssd1 vccd1 vccd1 _16380_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_319_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18118_ _18118_/A vssd1 vssd1 vccd1 vccd1 _18118_/X sky130_fd_sc_hd__buf_2
XFILLER_191_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19098_ _23239_/Q _18779_/X _19102_/S vssd1 vssd1 vccd1 vccd1 _19099_/A sky130_fd_sc_hd__mux2_1
XFILLER_306_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18049_ _22854_/Q _18036_/X _18037_/X _22987_/Q _18038_/X vssd1 vssd1 vccd1 vccd1
+ _18049_/X sky130_fd_sc_hd__a221o_1
XFILLER_160_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_321_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21060_ _21173_/A _21064_/B vssd1 vssd1 vccd1 vccd1 _21060_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20011_ _20016_/B _20016_/C _20010_/Y vssd1 vssd1 vccd1 vccd1 _23615_/D sky130_fd_sc_hd__o21a_1
XFILLER_298_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21962_ _22098_/A _22041_/B vssd1 vssd1 vccd1 vccd1 _21963_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23701_ _23706_/CLK _23701_/D vssd1 vssd1 vccd1 vccd1 _23701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20913_ _13910_/X _20908_/X _20601_/B _20912_/X vssd1 vssd1 vccd1 vccd1 _20913_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21893_ _20314_/Y _21892_/Y _22091_/B vssd1 vssd1 vccd1 vccd1 _21893_/X sky130_fd_sc_hd__mux2_1
XFILLER_254_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23632_ _23632_/CLK _23632_/D vssd1 vssd1 vccd1 vccd1 _23632_/Q sky130_fd_sc_hd__dfxtp_1
X_20844_ _20844_/A vssd1 vssd1 vccd1 vccd1 _23767_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23563_ _23563_/CLK _23563_/D vssd1 vssd1 vccd1 vccd1 _23563_/Q sky130_fd_sc_hd__dfxtp_1
X_20775_ _20865_/A vssd1 vssd1 vccd1 vccd1 _20811_/A sky130_fd_sc_hd__buf_4
XFILLER_147_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_390 _14088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22514_ _23692_/CLK _22514_/D vssd1 vssd1 vccd1 vccd1 _22514_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23494_ _23494_/CLK _23494_/D vssd1 vssd1 vccd1 vccd1 _23494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_356_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22445_ _23576_/CLK _22445_/D vssd1 vssd1 vccd1 vccd1 _22445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_324_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22376_ _23576_/CLK _22376_/D vssd1 vssd1 vccd1 vccd1 _22376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21327_ _21327_/A vssd1 vssd1 vccd1 vccd1 _21327_/X sky130_fd_sc_hd__buf_4
XFILLER_124_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12060_ _11217_/A _12050_/X _12059_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _13768_/A
+ sky130_fd_sc_hd__a211oi_4
X_21258_ _21258_/A _21258_/B vssd1 vssd1 vccd1 vccd1 _21259_/A sky130_fd_sc_hd__and2_1
XFILLER_296_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_289_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_289_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20209_ _20236_/A _20209_/B vssd1 vssd1 vccd1 vccd1 _20209_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21189_ _23878_/Q _21147_/X _21188_/X _21186_/X vssd1 vssd1 vccd1 vccd1 _23878_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_320_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_292_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15750_ _15749_/X _22280_/Q _15750_/S vssd1 vssd1 vccd1 vccd1 _15751_/A sky130_fd_sc_hd__mux2_1
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ _15753_/A _20327_/A _13500_/A vssd1 vssd1 vccd1 vccd1 _12964_/B sky130_fd_sc_hd__mux2_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_50 _20966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_61 _21209_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_72 _20148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14701_ input226/X _14980_/A _14700_/X vssd1 vssd1 vccd1 vccd1 _21348_/B sky130_fd_sc_hd__a21o_4
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_83 _11483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ _22365_/Q _22397_/Q _22686_/Q _23053_/Q _11648_/A _11653_/A vssd1 vssd1 vccd1
+ vccd1 _11914_/B sky130_fd_sc_hd__mux4_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_94 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15681_ _13387_/A _13629_/Y _15718_/B vssd1 vssd1 vccd1 vccd1 _15681_/X sky130_fd_sc_hd__mux2_1
X_12893_ _23932_/Q vssd1 vssd1 vccd1 vccd1 _12893_/Y sky130_fd_sc_hd__inv_2
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _17420_/A vssd1 vssd1 vccd1 vccd1 _22622_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_260_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _11844_/A vssd1 vssd1 vccd1 vccd1 _11844_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14632_ _14632_/A _14632_/B vssd1 vssd1 vccd1 vccd1 _14632_/Y sky130_fd_sc_hd__nor2_1
XFILLER_260_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _17351_/A vssd1 vssd1 vccd1 vccd1 _22596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _14563_/A vssd1 vssd1 vccd1 vccd1 _22261_/D sky130_fd_sc_hd__clkbuf_1
X_11775_ _22464_/Q _22624_/Q _11777_/S vssd1 vssd1 vccd1 vccd1 _11776_/B sky130_fd_sc_hd__mux2_1
XFILLER_348_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16302_/A vssd1 vssd1 vccd1 vccd1 _22322_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ _13514_/A _13514_/B vssd1 vssd1 vccd1 vccd1 _13514_/X sky130_fd_sc_hd__or2_1
X_17282_ _22139_/A _17281_/X _17292_/S vssd1 vssd1 vccd1 vccd1 _17282_/X sky130_fd_sc_hd__mux2_1
X_14494_ _23685_/Q _14488_/X _14494_/S vssd1 vssd1 vccd1 vccd1 _14494_/X sky130_fd_sc_hd__mux2_4
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_347_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19021_ _16813_/X _23205_/Q _19029_/S vssd1 vssd1 vccd1 vccd1 _19022_/A sky130_fd_sc_hd__mux2_1
X_13445_ _14180_/B vssd1 vssd1 vccd1 vccd1 _21079_/B sky130_fd_sc_hd__buf_4
X_16233_ _18798_/A vssd1 vssd1 vccd1 vccd1 _16233_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_277_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_357_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16164_ _21925_/A vssd1 vssd1 vccd1 vccd1 _21079_/A sky130_fd_sc_hd__buf_4
XFILLER_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13376_ _13382_/C _13376_/B vssd1 vssd1 vccd1 vccd1 _13379_/B sky130_fd_sc_hd__nand2_1
XFILLER_357_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_343_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15115_ _22494_/Q _13688_/A _15901_/A vssd1 vssd1 vccd1 vccd1 _15115_/X sky130_fd_sc_hd__o21a_1
X_12327_ _12586_/A _12327_/B vssd1 vssd1 vccd1 vccd1 _12327_/X sky130_fd_sc_hd__or2_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_303_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16095_ _11558_/B _15582_/B _15769_/A vssd1 vssd1 vccd1 vccd1 _16095_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_336_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_343_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19923_ _19923_/A _19923_/B _19927_/C vssd1 vssd1 vccd1 vccd1 _23591_/D sky130_fd_sc_hd__nor3_1
X_15046_ _15044_/X _22266_/Q _15284_/S vssd1 vssd1 vccd1 vccd1 _15047_/A sky130_fd_sc_hd__mux2_1
X_12258_ _12241_/A _12257_/X _11706_/A vssd1 vssd1 vccd1 vccd1 _12258_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_296_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11209_ _22808_/Q _22776_/Q _22677_/Q _22744_/Q _11206_/X _11208_/X vssd1 vssd1 vccd1
+ vccd1 _11209_/X sky130_fd_sc_hd__mux4_1
XFILLER_269_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19854_ _16220_/X _23561_/Q _19854_/S vssd1 vssd1 vccd1 vccd1 _19855_/A sky130_fd_sc_hd__mux2_1
X_12189_ _12307_/A _12189_/B vssd1 vssd1 vccd1 vccd1 _12189_/Y sky130_fd_sc_hd__nor2_1
XFILLER_311_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_295_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18805_ _18872_/S vssd1 vssd1 vccd1 vccd1 _18818_/S sky130_fd_sc_hd__buf_4
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19785_ _23530_/Q _19181_/A _19793_/S vssd1 vssd1 vccd1 vccd1 _19786_/A sky130_fd_sc_hd__mux2_1
XFILLER_256_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16997_ _17237_/A vssd1 vssd1 vccd1 vccd1 _16997_/X sky130_fd_sc_hd__buf_2
XFILLER_228_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_352_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_295_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18736_ _18736_/A vssd1 vssd1 vccd1 vccd1 _23093_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15948_ _14264_/X _15092_/X _15947_/X _15636_/X vssd1 vssd1 vccd1 vccd1 _15948_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18667_ _23063_/Q _17604_/X _18669_/S vssd1 vssd1 vccd1 vccd1 _18668_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15879_ _23740_/Q _23870_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _15879_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17618_ _22700_/Q _17617_/X _17624_/S vssd1 vssd1 vccd1 vccd1 _17619_/A sky130_fd_sc_hd__mux2_1
X_18598_ _18598_/A vssd1 vssd1 vccd1 vccd1 _23032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17549_ _17549_/A vssd1 vssd1 vccd1 vccd1 _22678_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_339_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20560_ _23717_/Q _20542_/X _20558_/X _20559_/X vssd1 vssd1 vccd1 vccd1 _23717_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_177_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19219_ _19219_/A vssd1 vssd1 vccd1 vccd1 _23285_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_93_wb_clk_i _22899_/CLK vssd1 vssd1 vccd1 vccd1 _23585_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20491_ _23716_/Q _20491_/B vssd1 vssd1 vccd1 vccd1 _20491_/X sky130_fd_sc_hd__or2_1
XFILLER_319_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_307_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_307_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22230_ _11270_/Y _22044_/X _22229_/X _22048_/X vssd1 vssd1 vccd1 vccd1 _22231_/B
+ sky130_fd_sc_hd__o22a_2
Xclkbuf_leaf_22_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23896_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_306_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22161_ _22161_/A _22161_/B vssd1 vssd1 vccd1 vccd1 _22162_/B sky130_fd_sc_hd__or2_1
XFILLER_105_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_306_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21112_ _23852_/Q _21110_/X _21111_/X _20597_/A vssd1 vssd1 vccd1 vccd1 _21113_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_172_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22092_ _21829_/B _22090_/Y _22091_/Y _21327_/A vssd1 vssd1 vccd1 vccd1 _22093_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_6919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21043_ _21153_/A _21043_/B vssd1 vssd1 vccd1 vccd1 _21043_/Y sky130_fd_sc_hd__nand2_1
XFILLER_275_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_287_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_286_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22994_ _23008_/CLK _22994_/D vssd1 vssd1 vccd1 vccd1 _22994_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_262_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21945_ _21945_/A _21944_/X vssd1 vssd1 vccd1 vccd1 _21947_/A sky130_fd_sc_hd__or2b_1
XFILLER_43_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21876_ _21876_/A _21876_/B vssd1 vssd1 vccd1 vccd1 _21876_/X sky130_fd_sc_hd__or2_1
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23615_ _23624_/CLK _23615_/D vssd1 vssd1 vccd1 vccd1 _23615_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20827_ _20881_/A vssd1 vssd1 vccd1 vccd1 _20843_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_30_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23546_ _23546_/CLK _23546_/D vssd1 vssd1 vccd1 vccd1 _23546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11560_ _11972_/A vssd1 vssd1 vccd1 vccd1 _11561_/A sky130_fd_sc_hd__buf_12
XFILLER_356_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20758_ _23746_/Q _20729_/X _20757_/X _20737_/X vssd1 vssd1 vccd1 vccd1 _23746_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_211_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_345_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23477_ _23541_/CLK _23477_/D vssd1 vssd1 vccd1 vccd1 _23477_/Q sky130_fd_sc_hd__dfxtp_4
X_11491_ _11497_/A _11491_/B vssd1 vssd1 vccd1 vccd1 _11491_/Y sky130_fd_sc_hd__nor2_1
XFILLER_210_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20689_ _20695_/A _20689_/B _20689_/C vssd1 vssd1 vccd1 vccd1 _20689_/X sky130_fd_sc_hd__or3_1
X_13230_ _22285_/Q _23101_/Q _23517_/Q _22446_/Q _11526_/A _11519_/A vssd1 vssd1 vccd1
+ vccd1 _13230_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22428_ _23466_/CLK _22428_/D vssd1 vssd1 vccd1 vccd1 _22428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ _13154_/Y _13156_/Y _13158_/Y _13160_/Y _11247_/A vssd1 vssd1 vccd1 vccd1
+ _13161_/X sky130_fd_sc_hd__o221a_1
XFILLER_298_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22359_ _23459_/CLK _22359_/D vssd1 vssd1 vccd1 vccd1 _22359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_325_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12112_ _12112_/A _12112_/B vssd1 vssd1 vccd1 vccd1 _12113_/B sky130_fd_sc_hd__and2_1
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13092_ _11196_/A _13090_/X _13206_/A vssd1 vssd1 vccd1 vccd1 _13092_/X sky130_fd_sc_hd__a21o_1
XFILLER_156_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12043_ _22468_/Q _22628_/Q _12043_/S vssd1 vssd1 vccd1 vccd1 _12043_/X sky130_fd_sc_hd__mux2_1
X_16920_ _16927_/A _16927_/B vssd1 vssd1 vccd1 vccd1 _17255_/A sky130_fd_sc_hd__or2_4
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_321_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16851_ _19201_/A vssd1 vssd1 vccd1 vccd1 _16851_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15802_ _15797_/Y _15800_/Y _15801_/X _14801_/A vssd1 vssd1 vccd1 vccd1 _15802_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19570_ _19570_/A vssd1 vssd1 vccd1 vccd1 _23434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_265_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16782_ _16782_/A vssd1 vssd1 vccd1 vccd1 _22511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13994_ _14074_/B vssd1 vssd1 vccd1 vccd1 _14046_/A sky130_fd_sc_hd__buf_2
XFILLER_19_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18521_ _18521_/A vssd1 vssd1 vccd1 vccd1 _18530_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_292_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15733_ _23704_/Q _15592_/A _15732_/X vssd1 vssd1 vccd1 vccd1 _15733_/Y sky130_fd_sc_hd__o21ai_4
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _23225_/Q _23193_/Q _23161_/Q _23129_/Q _12727_/X _12728_/X vssd1 vssd1 vccd1
+ vccd1 _12946_/B sky130_fd_sc_hd__mux4_2
XFILLER_292_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _18549_/A _18536_/A vssd1 vssd1 vccd1 vccd1 _18521_/A sky130_fd_sc_hd__or2_2
XFILLER_261_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _15564_/A _13608_/Y _15663_/X vssd1 vssd1 vccd1 vccd1 _15664_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _23226_/Q _23194_/Q _23162_/Q _23130_/Q _12750_/S _12672_/A vssd1 vssd1 vccd1
+ vccd1 _12877_/B sky130_fd_sc_hd__mux4_2
XFILLER_261_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _17403_/A vssd1 vssd1 vccd1 vccd1 _22614_/D sky130_fd_sc_hd__clkbuf_1
X_14615_ _14592_/X _14594_/X _14614_/X _14498_/X vssd1 vssd1 vccd1 vccd1 _14615_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_33_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _15207_/X _18384_/C _22955_/Q vssd1 vssd1 vccd1 vccd1 _18385_/B sky130_fd_sc_hd__a21oi_1
XFILLER_159_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11827_ _11275_/A _11811_/X _11826_/X _12594_/A vssd1 vssd1 vccd1 vccd1 _21616_/A
+ sky130_fd_sc_hd__o211a_4
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _15595_/A vssd1 vssd1 vccd1 vccd1 _15595_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17334_ _17334_/A vssd1 vssd1 vccd1 vccd1 _22589_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _22465_/Q _22625_/Q _22304_/Q _23440_/Q _11745_/X _12020_/A vssd1 vssd1 vccd1
+ vccd1 _11758_/X sky130_fd_sc_hd__mux4_1
X_14546_ _23887_/Q vssd1 vssd1 vccd1 vccd1 _14546_/X sky130_fd_sc_hd__buf_6
XFILLER_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17265_ _22578_/Q _17255_/X _17240_/X _17264_/X vssd1 vssd1 vccd1 vccd1 _22578_/D
+ sky130_fd_sc_hd__a211o_1
X_11689_ _21846_/A _20303_/A _12739_/A vssd1 vssd1 vccd1 vccd1 _13536_/B sky130_fd_sc_hd__mux2_2
X_14477_ _15596_/A vssd1 vssd1 vccd1 vccd1 _15216_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_329_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19004_ _16895_/X _23198_/Q _19012_/S vssd1 vssd1 vccd1 vccd1 _19005_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16216_ _16216_/A vssd1 vssd1 vccd1 vccd1 _22295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_335_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13428_ _13428_/A _13428_/B _13427_/X vssd1 vssd1 vccd1 vccd1 _13428_/X sky130_fd_sc_hd__or3b_1
XFILLER_127_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_351_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17196_ _17169_/X _17194_/X _17195_/X _17127_/X vssd1 vssd1 vccd1 vccd1 _17196_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_155_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_344_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16147_ _14896_/A _16133_/X _17307_/A _15436_/X vssd1 vssd1 vccd1 vccd1 _16147_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_13359_ _12546_/A _13359_/B _13361_/B vssd1 vssd1 vccd1 vccd1 _13360_/A sky130_fd_sc_hd__and3b_1
XFILLER_343_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_289_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16078_ _16151_/C _16078_/B vssd1 vssd1 vccd1 vccd1 _16079_/B sky130_fd_sc_hd__or2_1
XFILLER_303_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19906_ _19906_/A vssd1 vssd1 vccd1 vccd1 _23584_/D sky130_fd_sc_hd__clkbuf_1
X_15029_ _22508_/Q _14219_/A _13887_/A _15028_/X vssd1 vssd1 vccd1 vccd1 _15433_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_269_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_296_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19837_ _23554_/Q _19258_/A _19837_/S vssd1 vssd1 vccd1 vccd1 _19838_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_140_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _23846_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 coreIndex[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_4
X_19768_ _19768_/A vssd1 vssd1 vccd1 vccd1 _23523_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_284_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18719_ _16844_/X _23086_/Q _18719_/S vssd1 vssd1 vccd1 vccd1 _18720_/A sky130_fd_sc_hd__mux2_1
XFILLER_271_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19699_ _19699_/A _19699_/B vssd1 vssd1 vccd1 vccd1 _19756_/A sky130_fd_sc_hd__or2_4
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21730_ _21703_/B _21705_/B _21703_/A vssd1 vssd1 vccd1 vccd1 _21734_/A sky130_fd_sc_hd__o21ba_1
XFILLER_149_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21661_ _11068_/Y _15330_/A _21658_/Y _21659_/X _21660_/X vssd1 vssd1 vccd1 vccd1
+ _21661_/X sky130_fd_sc_hd__a221o_2
XFILLER_80_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23400_ _23526_/CLK _23400_/D vssd1 vssd1 vccd1 vccd1 _23400_/Q sky130_fd_sc_hd__dfxtp_1
X_20612_ _13931_/B _20563_/X _20611_/X vssd1 vssd1 vccd1 vccd1 _20613_/C sky130_fd_sc_hd__o21a_1
XFILLER_338_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21592_ _21591_/X _21574_/B _21572_/B vssd1 vssd1 vccd1 vccd1 _21593_/B sky130_fd_sc_hd__a21o_1
XFILLER_32_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23331_ _23491_/CLK _23331_/D vssd1 vssd1 vccd1 vccd1 _23331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20543_ _20543_/A vssd1 vssd1 vccd1 vccd1 _20547_/A sky130_fd_sc_hd__inv_2
XFILLER_338_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_327_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_353_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_326_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23262_ _23422_/CLK _23262_/D vssd1 vssd1 vccd1 vccd1 _23262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20474_ _21165_/A _20482_/B vssd1 vssd1 vccd1 vccd1 _20474_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22213_ _22213_/A _22213_/B vssd1 vssd1 vccd1 vccd1 _22213_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_106_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23193_ _23419_/CLK _23193_/D vssd1 vssd1 vccd1 vccd1 _23193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_307_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22144_ _22140_/B _21321_/A _21321_/B _21767_/A vssd1 vssd1 vccd1 vccd1 _22144_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_160_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput350 _13850_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[26] sky130_fd_sc_hd__buf_2
XFILLER_126_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput361 _13729_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[7] sky130_fd_sc_hd__buf_2
Xoutput372 _13653_/Y vssd1 vssd1 vccd1 vccd1 csb1[0] sky130_fd_sc_hd__buf_2
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22075_ _22100_/A _22075_/B vssd1 vssd1 vccd1 vccd1 _22155_/B sky130_fd_sc_hd__xnor2_1
Xoutput383 _14045_/X vssd1 vssd1 vccd1 vccd1 din0[18] sky130_fd_sc_hd__buf_2
XFILLER_121_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput394 _14065_/X vssd1 vssd1 vccd1 vccd1 din0[28] sky130_fd_sc_hd__buf_2
XFILLER_294_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_259_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21026_ _23825_/Q _20993_/X _21025_/Y _21023_/X vssd1 vssd1 vccd1 vccd1 _23825_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22977_ _22977_/CLK _22977_/D vssd1 vssd1 vccd1 vccd1 _22977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_308_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12730_ _12993_/A _12729_/X _12707_/A vssd1 vssd1 vccd1 vccd1 _12730_/X sky130_fd_sc_hd__o21a_1
XFILLER_27_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21928_ _21949_/A _22044_/A _21927_/X _21847_/A vssd1 vssd1 vccd1 vccd1 _22041_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _23945_/CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_271_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12661_ _12661_/A _12661_/B vssd1 vssd1 vccd1 vccd1 _12661_/Y sky130_fd_sc_hd__nand2_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21859_ _21856_/Y _21857_/X _21858_/Y vssd1 vssd1 vccd1 vccd1 _21859_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _22899_/Q _14394_/X _16929_/A _22592_/Q vssd1 vssd1 vccd1 vccd1 _22249_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _11621_/A vssd1 vssd1 vccd1 vccd1 _11613_/A sky130_fd_sc_hd__buf_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _15380_/A _15484_/B vssd1 vssd1 vccd1 vccd1 _15380_/Y sky130_fd_sc_hd__nand2_2
X_12592_ _12316_/A _12591_/X _11679_/A vssd1 vssd1 vccd1 vccd1 _12592_/X sky130_fd_sc_hd__o21a_1
XFILLER_357_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11543_ _11543_/A vssd1 vssd1 vccd1 vccd1 _11543_/X sky130_fd_sc_hd__buf_6
X_14331_ _14329_/X _14330_/X _14331_/S vssd1 vssd1 vccd1 vccd1 _14331_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23529_ _23529_/CLK _23529_/D vssd1 vssd1 vccd1 vccd1 _23529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_357_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_329_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_317_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17050_ _22558_/Q _17038_/X _17028_/X _17049_/X vssd1 vssd1 vccd1 vccd1 _22558_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_156_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14262_ _15455_/A vssd1 vssd1 vccd1 vccd1 _15798_/A sky130_fd_sc_hd__clkbuf_2
X_11474_ _11464_/Y _11467_/Y _11471_/Y _11473_/Y _21898_/A vssd1 vssd1 vccd1 vccd1
+ _11485_/B sky130_fd_sc_hd__o221a_1
XFILLER_13_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_326_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13213_ _11247_/X _11398_/A _11403_/X _13212_/Y vssd1 vssd1 vccd1 vccd1 _13242_/A
+ sky130_fd_sc_hd__a22o_4
X_16001_ _15964_/A _17269_/A _16000_/X vssd1 vssd1 vccd1 vccd1 _16001_/X sky130_fd_sc_hd__o21a_1
XFILLER_183_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14193_ _20532_/C vssd1 vssd1 vccd1 vccd1 _14193_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_326_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_298_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_317_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13144_ _22318_/Q _23454_/Q _13190_/S vssd1 vssd1 vccd1 vccd1 _13144_/X sky130_fd_sc_hd__mux2_1
XFILLER_325_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_317_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_297_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17952_ _22827_/Q _17938_/X _17939_/X input273/X _17951_/X vssd1 vssd1 vccd1 vccd1
+ _17952_/X sky130_fd_sc_hd__a221o_1
XFILLER_341_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13075_ _13121_/A _13074_/X _11537_/X vssd1 vssd1 vccd1 vccd1 _13075_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_297_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16903_ _16902_/X _22548_/Q _16909_/S vssd1 vssd1 vccd1 vccd1 _16904_/A sky130_fd_sc_hd__mux2_1
X_12026_ _23219_/Q _23187_/Q _23155_/Q _23123_/Q _12024_/X _12025_/X vssd1 vssd1 vccd1
+ vccd1 _12027_/B sky130_fd_sc_hd__mux4_1
XFILLER_250_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17883_ _17883_/A vssd1 vssd1 vccd1 vccd1 _22812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19622_ _19622_/A vssd1 vssd1 vccd1 vccd1 _23458_/D sky130_fd_sc_hd__clkbuf_1
X_16834_ _16834_/A vssd1 vssd1 vccd1 vccd1 _22526_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_333_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19553_ _19264_/X _23428_/Q _19553_/S vssd1 vssd1 vccd1 vccd1 _19554_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16765_ _16783_/A vssd1 vssd1 vccd1 vccd1 _16765_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13977_ _13977_/A _13979_/B vssd1 vssd1 vccd1 vccd1 _13978_/A sky130_fd_sc_hd__and2_1
XFILLER_20_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18504_ _18494_/X _18502_/Y _18503_/X vssd1 vssd1 vccd1 vccd1 _22996_/D sky130_fd_sc_hd__a21oi_1
XFILLER_206_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15716_ _15790_/C _15716_/B vssd1 vssd1 vccd1 vccd1 _15716_/X sky130_fd_sc_hd__or2_4
X_12928_ _12968_/A _12927_/X _12687_/X vssd1 vssd1 vccd1 vccd1 _12928_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_207_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19484_ _19540_/A vssd1 vssd1 vccd1 vccd1 _19553_/S sky130_fd_sc_hd__buf_6
XFILLER_80_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16696_ _16696_/A vssd1 vssd1 vccd1 vccd1 _22487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18435_ _18435_/A _22973_/Q _18435_/C vssd1 vssd1 vccd1 vccd1 _18440_/C sky130_fd_sc_hd__and3_1
XFILLER_221_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15647_ _23734_/Q _23864_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _15647_/X sky130_fd_sc_hd__mux2_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _22800_/Q _22768_/Q _22669_/Q _22736_/Q _12843_/X _12844_/X vssd1 vssd1 vccd1
+ vccd1 _12860_/B sky130_fd_sc_hd__mux4_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_349_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18366_ _22948_/Q _22949_/Q _18366_/C vssd1 vssd1 vccd1 vccd1 _18369_/B sky130_fd_sc_hd__and3_1
X_15578_ _15578_/A vssd1 vssd1 vccd1 vccd1 _15674_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17317_ _21079_/A _17316_/X _17317_/S vssd1 vssd1 vccd1 vccd1 _17317_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_308_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14529_ _14529_/A _15519_/A vssd1 vssd1 vccd1 vccd1 _15048_/A sky130_fd_sc_hd__nor2_2
XFILLER_336_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18297_ _18315_/A _18297_/B _18297_/C vssd1 vssd1 vccd1 vccd1 _22925_/D sky130_fd_sc_hd__nor3_1
XFILLER_147_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_335_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17248_ _17248_/A vssd1 vssd1 vccd1 vccd1 _17291_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_179_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17179_ input88/X input52/X _17200_/S vssd1 vssd1 vccd1 vccd1 _17179_/X sky130_fd_sc_hd__mux2_8
XFILLER_227_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_350_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_304_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_288_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20190_ _20250_/A _20190_/B vssd1 vssd1 vccd1 vccd1 _20190_/Y sky130_fd_sc_hd__nand2_1
XFILLER_304_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_331_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22900_ _22908_/CLK _22900_/D vssd1 vssd1 vccd1 vccd1 _22900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_300_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23880_ _23880_/CLK _23880_/D vssd1 vssd1 vccd1 vccd1 _23880_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22831_ _22893_/CLK _22831_/D vssd1 vssd1 vccd1 vccd1 _22831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22762_ _23446_/CLK _22762_/D vssd1 vssd1 vccd1 vccd1 _22762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21713_ _22061_/A _21706_/X _21712_/X _21408_/X vssd1 vssd1 vccd1 vccd1 _21714_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22693_ _23572_/CLK _22693_/D vssd1 vssd1 vccd1 vccd1 _22693_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21644_ _21081_/A _21626_/X _21633_/X _22215_/A _21643_/Y vssd1 vssd1 vccd1 vccd1
+ _21644_/X sky130_fd_sc_hd__a221o_1
XFILLER_200_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21575_ _21575_/A vssd1 vssd1 vccd1 vccd1 _22032_/B sky130_fd_sc_hd__buf_2
XFILLER_354_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23314_ _23538_/CLK _23314_/D vssd1 vssd1 vccd1 vccd1 _23314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20526_ _20526_/A _20526_/B _20526_/C vssd1 vssd1 vccd1 vccd1 _20531_/B sky130_fd_sc_hd__or3_2
XFILLER_315_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_354_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23245_ _23534_/CLK _23245_/D vssd1 vssd1 vccd1 vccd1 _23245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_342_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_1_0_wb_clk_i _23931_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_20457_ _23702_/Q _20468_/B vssd1 vssd1 vccd1 vccd1 _20457_/X sky130_fd_sc_hd__or2_1
XFILLER_137_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_7203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_7225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23176_ _23528_/CLK _23176_/D vssd1 vssd1 vccd1 vccd1 _23176_/Q sky130_fd_sc_hd__dfxtp_1
X_11190_ _12536_/A vssd1 vssd1 vccd1 vccd1 _12423_/A sky130_fd_sc_hd__buf_4
XFILLER_323_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_322_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20388_ _17298_/A _20261_/X _20389_/B vssd1 vssd1 vccd1 vccd1 _20388_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_107_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_350_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22127_ _22231_/A _22127_/B vssd1 vssd1 vccd1 vccd1 _22155_/D sky130_fd_sc_hd__xnor2_1
XFILLER_134_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_322_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_350_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_294_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22058_ _22024_/A _22024_/B _22023_/A vssd1 vssd1 vccd1 vccd1 _22059_/B sky130_fd_sc_hd__a21oi_1
XTAP_6579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21009_ _23819_/Q _21009_/B vssd1 vssd1 vccd1 vccd1 _21009_/X sky130_fd_sc_hd__or2_1
X_13900_ _13933_/A _14082_/A vssd1 vssd1 vccd1 vccd1 _13900_/Y sky130_fd_sc_hd__nor2_4
XTAP_5867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14880_ _14520_/A _14863_/X _14867_/X _14879_/X _14587_/X vssd1 vssd1 vccd1 vccd1
+ _14880_/X sky130_fd_sc_hd__a32o_1
XTAP_5889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_303_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_290_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13831_ _14216_/A _13831_/B vssd1 vssd1 vccd1 vccd1 _13832_/A sky130_fd_sc_hd__nor2_1
XFILLER_291_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16550_ _16550_/A vssd1 vssd1 vccd1 vccd1 _22427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_208 _15596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13762_ _14198_/B _20530_/B vssd1 vssd1 vccd1 vccd1 _14207_/A sky130_fd_sc_hd__nand2_2
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_219 _14879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15501_ _15501_/A _15501_/B vssd1 vssd1 vccd1 vccd1 _15501_/X sky130_fd_sc_hd__or2_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12713_ _12958_/A vssd1 vssd1 vccd1 vccd1 _12995_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16481_ _16481_/A vssd1 vssd1 vccd1 vccd1 _22398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13693_ _13934_/A vssd1 vssd1 vccd1 vccd1 _13969_/A sky130_fd_sc_hd__inv_2
XFILLER_16_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18220_ _22851_/Q _18216_/X _18218_/X _18219_/X vssd1 vssd1 vccd1 vccd1 _22899_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_231_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15432_ _15432_/A _15432_/B vssd1 vssd1 vccd1 vccd1 _15432_/Y sky130_fd_sc_hd__nand2_2
XFILLER_188_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12644_ _23221_/Q _23189_/Q _23157_/Q _23125_/Q _12751_/S _12671_/A vssd1 vssd1 vccd1
+ vccd1 _12645_/B sky130_fd_sc_hd__mux4_2
XPHY_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18151_ _18151_/A vssd1 vssd1 vccd1 vccd1 _22886_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12575_ _11216_/A _12371_/B _12574_/X _11828_/B vssd1 vssd1 vccd1 vccd1 _14368_/A
+ sky130_fd_sc_hd__o211ai_4
X_15363_ _15697_/A _17103_/A vssd1 vssd1 vccd1 vccd1 _15363_/Y sky130_fd_sc_hd__nor2_1
XPHY_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_317_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17102_ input80/X input45/X _17132_/S vssd1 vssd1 vccd1 vccd1 _17102_/X sky130_fd_sc_hd__mux2_8
XFILLER_357_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14314_ _14296_/X _14312_/X _15130_/S vssd1 vssd1 vccd1 vccd1 _15541_/A sky130_fd_sc_hd__mux2_1
XFILLER_345_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18082_ _18097_/A vssd1 vssd1 vccd1 vccd1 _18082_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11526_ _11526_/A vssd1 vssd1 vccd1 vccd1 _13275_/A sky130_fd_sc_hd__buf_4
XFILLER_172_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15294_ _14671_/S _15293_/Y _15253_/X vssd1 vssd1 vccd1 vccd1 _15798_/B sky130_fd_sc_hd__a21o_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17033_ _17033_/A _17033_/B vssd1 vssd1 vccd1 vccd1 _17033_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14245_ input132/X input107/X _15052_/S vssd1 vssd1 vccd1 vccd1 _14245_/X sky130_fd_sc_hd__mux2_8
X_11457_ _11863_/A _11457_/B _11457_/C _11457_/D vssd1 vssd1 vccd1 vccd1 _12414_/A
+ sky130_fd_sc_hd__nor4_4
XFILLER_332_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_314_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14176_ _14176_/A _20139_/A vssd1 vssd1 vccd1 vccd1 _15455_/A sky130_fd_sc_hd__nand2_4
XFILLER_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11388_ _12913_/S vssd1 vssd1 vccd1 vccd1 _13234_/S sky130_fd_sc_hd__clkbuf_4
X_13127_ _13127_/A vssd1 vssd1 vccd1 vccd1 _13127_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_314_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18984_ _16867_/X _23189_/Q _18990_/S vssd1 vssd1 vccd1 vccd1 _18985_/A sky130_fd_sc_hd__mux2_1
XFILLER_344_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_298_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17935_ _22823_/Q _17932_/X _17934_/X _17930_/X vssd1 vssd1 vccd1 vccd1 _22823_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13058_ _23938_/Q vssd1 vssd1 vccd1 vccd1 _22140_/A sky130_fd_sc_hd__inv_2
XFILLER_79_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12009_ _12009_/A vssd1 vssd1 vccd1 vccd1 _12009_/X sky130_fd_sc_hd__buf_8
XFILLER_239_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17866_ _22804_/Q _17633_/X _17870_/S vssd1 vssd1 vccd1 vccd1 _17867_/A sky130_fd_sc_hd__mux2_1
XFILLER_254_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19605_ _19605_/A vssd1 vssd1 vccd1 vccd1 _23450_/D sky130_fd_sc_hd__clkbuf_1
X_16817_ _16813_/X _22521_/Q _16829_/S vssd1 vssd1 vccd1 vccd1 _16818_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17797_ _17797_/A vssd1 vssd1 vccd1 vccd1 _22773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19536_ _19239_/X _23420_/Q _19538_/S vssd1 vssd1 vccd1 vccd1 _19537_/A sky130_fd_sc_hd__mux2_1
XFILLER_281_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16748_ _16784_/A vssd1 vssd1 vccd1 vccd1 _16748_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_289_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19467_ _19467_/A vssd1 vssd1 vccd1 vccd1 _23389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16679_ _16679_/A _16679_/B vssd1 vssd1 vccd1 vccd1 _16679_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18418_ _18418_/A _22967_/Q _18418_/C vssd1 vssd1 vccd1 vccd1 _18420_/B sky130_fd_sc_hd__and3_1
XFILLER_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19398_ _19398_/A vssd1 vssd1 vccd1 vccd1 _23358_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_349_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18349_ _22942_/Q _22943_/Q _18349_/C vssd1 vssd1 vccd1 vccd1 _18351_/B sky130_fd_sc_hd__and3_1
XFILLER_159_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_309_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_296_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21360_ _23749_/Q _21816_/A _23815_/Q vssd1 vssd1 vccd1 vccd1 _21361_/C sky130_fd_sc_hd__a21oi_1
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20311_ _21871_/A _20394_/B vssd1 vssd1 vccd1 vccd1 _20313_/B sky130_fd_sc_hd__nand2_1
XFILLER_352_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_323_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21291_ _22895_/Q _22894_/Q vssd1 vssd1 vccd1 vccd1 _21291_/X sky130_fd_sc_hd__or2_2
XFILLER_162_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput60 dout0[25] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__buf_2
Xinput71 dout0[35] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_1
Xinput82 dout0[45] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__clkbuf_1
X_23030_ _23414_/CLK _23030_/D vssd1 vssd1 vccd1 vccd1 _23030_/Q sky130_fd_sc_hd__dfxtp_1
Xinput93 dout0[55] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20242_ _15271_/X _20169_/A _20243_/B vssd1 vssd1 vccd1 vccd1 _20242_/X sky130_fd_sc_hd__a21o_1
XFILLER_116_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_305_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20173_ _20250_/A vssd1 vssd1 vccd1 vccd1 _20355_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_277_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23932_ _23942_/CLK _23932_/D vssd1 vssd1 vccd1 vccd1 _23932_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23863_ _23874_/CLK _23863_/D vssd1 vssd1 vccd1 vccd1 _23863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_272_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22814_ _22822_/CLK _22814_/D vssd1 vssd1 vccd1 vccd1 _22814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23794_ _23861_/CLK _23794_/D vssd1 vssd1 vccd1 vccd1 _23794_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_225_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_344_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22745_ _23555_/CLK _22745_/D vssd1 vssd1 vccd1 vccd1 _22745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22676_ _23893_/CLK _22676_/D vssd1 vssd1 vccd1 vccd1 _22676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_328_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21627_ _23823_/Q _23757_/Q vssd1 vssd1 vccd1 vccd1 _21627_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_327_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12360_ _23400_/Q _23016_/Q _23368_/Q _23336_/Q _11112_/A _12458_/A vssd1 vssd1 vccd1
+ vccd1 _12360_/X sky130_fd_sc_hd__mux4_1
X_21558_ _21558_/A _21605_/C vssd1 vssd1 vccd1 vccd1 _21559_/B sky130_fd_sc_hd__xor2_4
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11311_ _11311_/A vssd1 vssd1 vccd1 vccd1 _11364_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_148_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20509_ _20509_/A _20509_/B _20509_/C _20509_/D vssd1 vssd1 vccd1 vccd1 _20531_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_343_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12291_ _12291_/A _12291_/B vssd1 vssd1 vccd1 vccd1 _12291_/Y sky130_fd_sc_hd__nor2_1
XFILLER_314_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21489_ _21942_/A _21489_/B vssd1 vssd1 vccd1 vccd1 _21489_/Y sky130_fd_sc_hd__nor2_1
X_14030_ _14023_/X _13756_/B _14013_/X input217/X vssd1 vssd1 vccd1 vccd1 _14030_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_7000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23228_ _23419_/CLK _23228_/D vssd1 vssd1 vccd1 vccd1 _23228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11242_ _11242_/A vssd1 vssd1 vccd1 vccd1 _11243_/A sky130_fd_sc_hd__clkbuf_8
XTAP_7011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_351_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23159_ _23543_/CLK _23159_/D vssd1 vssd1 vccd1 vccd1 _23159_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11173_ _23901_/Q vssd1 vssd1 vccd1 vccd1 _11603_/A sky130_fd_sc_hd__inv_2
XFILLER_350_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_310_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15981_ _22940_/Q _14752_/X _14753_/X _18435_/A vssd1 vssd1 vccd1 vccd1 _15981_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_311_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17720_ _22739_/Q _17630_/X _17726_/S vssd1 vssd1 vccd1 vccd1 _17721_/A sky130_fd_sc_hd__mux2_1
XTAP_6387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14932_ _15000_/A vssd1 vssd1 vccd1 vccd1 _14932_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ _20508_/B _17653_/B _17650_/Y _17390_/X vssd1 vssd1 vccd1 vccd1 _22710_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ _20186_/A _13903_/A _14838_/X _14862_/Y vssd1 vssd1 vccd1 vccd1 _14863_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_291_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16602_ _16602_/A vssd1 vssd1 vccd1 vccd1 _22451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13814_ _12891_/B _13836_/B _13746_/X vssd1 vssd1 vccd1 vccd1 _13814_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_291_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17582_ _18808_/A vssd1 vssd1 vccd1 vccd1 _17582_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14794_ _14794_/A _14794_/B vssd1 vssd1 vccd1 vccd1 _14794_/Y sky130_fd_sc_hd__nand2_1
XFILLER_235_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19321_ _19321_/A vssd1 vssd1 vccd1 vccd1 _23324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16533_ _18476_/A vssd1 vssd1 vccd1 vccd1 _20134_/A sky130_fd_sc_hd__buf_6
XFILLER_250_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13745_ _13745_/A _13745_/B vssd1 vssd1 vccd1 vccd1 _13842_/A sky130_fd_sc_hd__nand2_2
XFILLER_17_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19252_ _19252_/A vssd1 vssd1 vccd1 vccd1 _19252_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16464_ _16464_/A vssd1 vssd1 vccd1 vccd1 _22390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13676_ _22421_/Q _16534_/B _13666_/X vssd1 vssd1 vccd1 vccd1 _13679_/B sky130_fd_sc_hd__o21ai_4
XFILLER_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18203_ _22872_/Q _18203_/B _18203_/C vssd1 vssd1 vccd1 vccd1 _18243_/A sky130_fd_sc_hd__nor3_4
X_15415_ _15081_/A _15375_/X _15412_/X _15414_/X vssd1 vssd1 vccd1 vccd1 _15415_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_129_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12627_ _22373_/Q _22405_/Q _22694_/Q _23061_/Q _12013_/X _12717_/A vssd1 vssd1 vccd1
+ vccd1 _12627_/X sky130_fd_sc_hd__mux4_2
XPHY_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19183_ _19181_/X _23274_/Q _19195_/S vssd1 vssd1 vccd1 vccd1 _19184_/A sky130_fd_sc_hd__mux2_1
XPHY_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16395_ _16395_/A vssd1 vssd1 vccd1 vccd1 _22360_/D sky130_fd_sc_hd__clkbuf_1
XPHY_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_318_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18134_ _18116_/Y _18132_/X _18133_/X _18121_/X vssd1 vssd1 vccd1 vccd1 _22882_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15346_ _15346_/A _15346_/B vssd1 vssd1 vccd1 vccd1 _15832_/A sky130_fd_sc_hd__or2_2
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12558_ _11837_/A _12554_/X _12557_/X _12567_/A vssd1 vssd1 vccd1 vccd1 _12558_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_319_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18065_ _22860_/Q _18051_/X _18064_/X _18060_/X vssd1 vssd1 vccd1 vccd1 _22860_/D
+ sky130_fd_sc_hd__o211a_1
X_11509_ _11502_/Y _11504_/Y _11506_/Y _11508_/Y _11247_/X vssd1 vssd1 vccd1 vccd1
+ _11509_/X sky130_fd_sc_hd__o221a_1
XFILLER_176_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15277_ _15318_/A _15277_/B vssd1 vssd1 vccd1 vccd1 _15277_/Y sky130_fd_sc_hd__nor2_1
XFILLER_333_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12489_ _12489_/A _12489_/B vssd1 vssd1 vccd1 vccd1 _12489_/X sky130_fd_sc_hd__or2_1
XFILLER_176_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17016_ _17145_/A vssd1 vssd1 vccd1 vccd1 _17016_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14228_ input158/X input123/X _15030_/S vssd1 vssd1 vccd1 vccd1 _14228_/X sky130_fd_sc_hd__mux2_8
XFILLER_299_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14159_ _14159_/A vssd1 vssd1 vccd1 vccd1 _14394_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18967_ _18967_/A vssd1 vssd1 vccd1 vccd1 _23181_/D sky130_fd_sc_hd__clkbuf_1
X_17918_ _17959_/A vssd1 vssd1 vccd1 vccd1 _17918_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_47_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23504_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_267_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18898_ _18944_/S vssd1 vssd1 vccd1 vccd1 _18907_/S sky130_fd_sc_hd__buf_4
XFILLER_254_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17849_ _17849_/A vssd1 vssd1 vccd1 vccd1 _22796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20860_ _20721_/B _20846_/X _20847_/X _23772_/Q vssd1 vssd1 vccd1 vccd1 _20861_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_214_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19519_ _19213_/X _23412_/Q _19527_/S vssd1 vssd1 vccd1 vccd1 _19520_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20791_ _20810_/A vssd1 vssd1 vccd1 vccd1 _20791_/X sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_550 _17385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_561 _23882_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22530_ _23502_/CLK _22530_/D vssd1 vssd1 vccd1 vccd1 _22530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22461_ _23368_/CLK _22461_/D vssd1 vssd1 vccd1 vccd1 _22461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_349_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21412_ _21400_/A _21366_/X _21378_/X _21411_/Y _21175_/X vssd1 vssd1 vccd1 vccd1
+ _23914_/D sky130_fd_sc_hd__o221a_1
X_22392_ _23496_/CLK _22392_/D vssd1 vssd1 vccd1 vccd1 _22392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_337_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21343_ _21344_/A _21344_/B vssd1 vssd1 vccd1 vccd1 _21345_/A sky130_fd_sc_hd__and2_1
XFILLER_325_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_324_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21274_ _21274_/A _21274_/B vssd1 vssd1 vccd1 vccd1 _21274_/Y sky130_fd_sc_hd__nand2_1
XFILLER_190_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23013_ _23525_/CLK _23013_/D vssd1 vssd1 vccd1 vccd1 _23013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20225_ _20404_/B vssd1 vssd1 vccd1 vccd1 _20323_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20156_ _20186_/A _20186_/B vssd1 vssd1 vccd1 vccd1 _20174_/A sky130_fd_sc_hd__or2_2
XFILLER_320_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20087_ _23637_/Q _20095_/D vssd1 vssd1 vccd1 vccd1 _20088_/B sky130_fd_sc_hd__xnor2_1
XFILLER_287_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23915_ _23915_/CLK _23915_/D vssd1 vssd1 vccd1 vccd1 _23915_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23846_ _23846_/CLK _23846_/D vssd1 vssd1 vccd1 vccd1 _23846_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _22270_/Q _23086_/Q _23502_/Q _22431_/Q _12094_/A _11754_/A vssd1 vssd1 vccd1
+ vccd1 _11861_/B sky130_fd_sc_hd__mux4_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11791_ _11774_/A _11790_/X _11706_/X vssd1 vssd1 vccd1 vccd1 _11791_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20989_ _20989_/A _20989_/B _20989_/C _21084_/B vssd1 vssd1 vccd1 vccd1 _21051_/A
+ sky130_fd_sc_hd__nor4_4
X_23777_ _23804_/CLK _23777_/D vssd1 vssd1 vccd1 vccd1 _23777_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13530_ _13618_/B _13618_/C _13618_/A vssd1 vssd1 vccd1 vccd1 _13619_/A sky130_fd_sc_hd__a21oi_4
X_22728_ _23450_/CLK _22728_/D vssd1 vssd1 vccd1 vccd1 _22728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_335_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13461_ _23946_/Q vssd1 vssd1 vccd1 vccd1 _13471_/A sky130_fd_sc_hd__inv_2
XFILLER_201_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22659_ _23567_/CLK _22659_/D vssd1 vssd1 vccd1 vccd1 _22659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_328_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15200_ _14370_/X _14371_/Y _14175_/Y vssd1 vssd1 vccd1 vccd1 _15495_/A sky130_fd_sc_hd__o21ai_2
XFILLER_159_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12412_ _12397_/A _12411_/X _11347_/A vssd1 vssd1 vccd1 vccd1 _12412_/Y sky130_fd_sc_hd__o21ai_1
X_16180_ _16191_/B _16180_/B vssd1 vssd1 vccd1 vccd1 _16180_/Y sky130_fd_sc_hd__nor2_1
X_13392_ _13392_/A _13392_/B vssd1 vssd1 vccd1 vccd1 _13393_/B sky130_fd_sc_hd__nor2_2
XFILLER_355_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15131_ _15131_/A vssd1 vssd1 vccd1 vccd1 _15131_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12343_ _14371_/B _20139_/A _14371_/A vssd1 vssd1 vccd1 vccd1 _14385_/A sky130_fd_sc_hd__a21oi_2
XFILLER_327_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15062_ _14218_/X _15484_/A _15061_/X _13706_/A vssd1 vssd1 vccd1 vccd1 _15062_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_175_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12274_ _12410_/A _12274_/B vssd1 vssd1 vccd1 vccd1 _12274_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_342_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11225_ _15826_/A _11224_/X _15864_/A vssd1 vssd1 vccd1 vccd1 _11225_/Y sky130_fd_sc_hd__o21ai_1
X_14013_ _14041_/A vssd1 vssd1 vccd1 vccd1 _14013_/X sky130_fd_sc_hd__buf_2
XFILLER_296_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19870_ _16243_/X _23568_/Q _19876_/S vssd1 vssd1 vccd1 vccd1 _19871_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18821_ _18853_/A vssd1 vssd1 vccd1 vccd1 _18834_/S sky130_fd_sc_hd__buf_2
XFILLER_295_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11156_ _13190_/S vssd1 vssd1 vccd1 vccd1 _11493_/S sky130_fd_sc_hd__buf_6
XFILLER_136_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_310_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18752_ _16892_/X _23101_/Q _18752_/S vssd1 vssd1 vccd1 vccd1 _18753_/A sky130_fd_sc_hd__mux2_1
XTAP_6184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15964_ _15964_/A _17258_/A vssd1 vssd1 vccd1 vccd1 _15964_/Y sky130_fd_sc_hd__nor2_1
X_11087_ _23892_/Q _23891_/Q vssd1 vssd1 vccd1 vccd1 _11095_/B sky130_fd_sc_hd__and2_1
XTAP_6195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput250 localMemory_wb_sel_i[3] vssd1 vssd1 vccd1 vccd1 input250/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput261 manufacturerID[7] vssd1 vssd1 vccd1 vccd1 _17926_/A sky130_fd_sc_hd__clkbuf_2
X_17703_ _17703_/A vssd1 vssd1 vccd1 vccd1 _22731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_264_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput272 partID[2] vssd1 vssd1 vccd1 vccd1 _17944_/A sky130_fd_sc_hd__clkbuf_1
XTAP_5483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14915_ _23721_/Q _23851_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _14915_/X sky130_fd_sc_hd__mux2_4
Xinput283 versionID[3] vssd1 vssd1 vccd1 vccd1 input283/X sky130_fd_sc_hd__clkbuf_2
X_18683_ _23070_/Q _17626_/X _18691_/S vssd1 vssd1 vccd1 vccd1 _18684_/A sky130_fd_sc_hd__mux2_1
XTAP_5494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15895_ _23001_/Q _15931_/A _15932_/A input230/X vssd1 vssd1 vccd1 vccd1 _22032_/A
+ sky130_fd_sc_hd__a22o_4
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17634_ _22705_/Q _17633_/X _17640_/S vssd1 vssd1 vccd1 vccd1 _17635_/A sky130_fd_sc_hd__mux2_1
XFILLER_286_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14846_ _14657_/X _14633_/X _14850_/S vssd1 vssd1 vccd1 vccd1 _14846_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17565_ _17565_/A vssd1 vssd1 vccd1 vccd1 _22683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14777_ _14310_/X _14272_/X _14850_/S vssd1 vssd1 vccd1 vccd1 _14778_/A sky130_fd_sc_hd__mux2_1
X_11989_ _12141_/A _11989_/B vssd1 vssd1 vccd1 vccd1 _11989_/X sky130_fd_sc_hd__or2_1
X_19304_ _19304_/A vssd1 vssd1 vccd1 vccd1 _23316_/D sky130_fd_sc_hd__clkbuf_1
X_16516_ _15975_/X _22414_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _16517_/A sky130_fd_sc_hd__mux2_1
X_13728_ _14015_/A _13728_/B _14021_/C vssd1 vssd1 vccd1 vccd1 _13729_/A sky130_fd_sc_hd__and3_4
X_17496_ _17542_/S vssd1 vssd1 vccd1 vccd1 _17505_/S sky130_fd_sc_hd__buf_4
XFILLER_210_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_165_wb_clk_i _23917_/CLK vssd1 vssd1 vccd1 vccd1 _23918_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19235_ _19235_/A vssd1 vssd1 vccd1 vccd1 _23290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16447_ _16049_/X _22384_/Q _16451_/S vssd1 vssd1 vccd1 vccd1 _16448_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13659_ _13669_/A _22612_/Q vssd1 vssd1 vccd1 vccd1 _14211_/A sky130_fd_sc_hd__and2_2
XFILLER_286_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19166_ _19265_/S vssd1 vssd1 vccd1 vccd1 _19179_/S sky130_fd_sc_hd__buf_6
X_16378_ _16378_/A vssd1 vssd1 vccd1 vccd1 _22354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_334_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18117_ _14121_/D _18009_/B _18126_/S vssd1 vssd1 vccd1 vccd1 _18117_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15329_ _15329_/A _15376_/C vssd1 vssd1 vccd1 vccd1 _15330_/A sky130_fd_sc_hd__xnor2_1
X_19097_ _19097_/A vssd1 vssd1 vccd1 vccd1 _23238_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_322_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18048_ _22854_/Q _18035_/X _18047_/X _18045_/X vssd1 vssd1 vccd1 vccd1 _22854_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_321_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20010_ _20016_/B _20016_/C _19962_/X vssd1 vssd1 vccd1 vccd1 _20010_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_286_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19999_ _20009_/A _20009_/B _19998_/Y vssd1 vssd1 vccd1 vccd1 _23612_/D sky130_fd_sc_hd__o21a_1
XFILLER_287_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_286_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21961_ _22098_/A _22041_/B vssd1 vssd1 vccd1 vccd1 _21961_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23700_ _23700_/CLK _23700_/D vssd1 vssd1 vccd1 vccd1 _23700_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20912_ _20926_/A vssd1 vssd1 vccd1 vccd1 _20912_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_215_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21892_ _21892_/A _21892_/B vssd1 vssd1 vccd1 vccd1 _21892_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_81_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23631_ _23634_/CLK _23631_/D vssd1 vssd1 vccd1 vccd1 _23631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_270_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20843_ _20843_/A _20843_/B vssd1 vssd1 vccd1 vccd1 _20844_/A sky130_fd_sc_hd__and2_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23562_ _23564_/CLK _23562_/D vssd1 vssd1 vccd1 vccd1 _23562_/Q sky130_fd_sc_hd__dfxtp_1
X_20774_ _20774_/A _20864_/A vssd1 vssd1 vccd1 vccd1 _20865_/A sky130_fd_sc_hd__nor2_4
XFILLER_329_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_380 _22513_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_391 _14090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22513_ _23693_/CLK _22513_/D vssd1 vssd1 vccd1 vccd1 _22513_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23493_ _23493_/CLK _23493_/D vssd1 vssd1 vccd1 vccd1 _23493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22444_ _23453_/CLK _22444_/D vssd1 vssd1 vccd1 vccd1 _22444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_337_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22375_ _23544_/CLK _22375_/D vssd1 vssd1 vccd1 vccd1 _22375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_309_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_352_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_324_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21326_ _21677_/A vssd1 vssd1 vccd1 vccd1 _21327_/A sky130_fd_sc_hd__buf_2
XFILLER_135_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_340_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21257_ _13454_/A _15754_/X _21257_/S vssd1 vssd1 vccd1 vccd1 _21258_/B sky130_fd_sc_hd__mux2_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_292_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_321_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20208_ _15005_/B _20154_/X _20209_/B vssd1 vssd1 vccd1 vccd1 _20208_/X sky130_fd_sc_hd__a21o_1
X_21188_ _20765_/A _21158_/A _21142_/A _20515_/C _21150_/A vssd1 vssd1 vccd1 vccd1
+ _21188_/X sky130_fd_sc_hd__a221o_1
XFILLER_145_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_320_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20139_ _20139_/A _20532_/B vssd1 vssd1 vccd1 vccd1 _20139_/Y sky130_fd_sc_hd__nor2_2
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12961_ _11277_/A _12951_/X _12960_/X _12864_/A vssd1 vssd1 vccd1 vccd1 _20327_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_161_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_40 _20404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_51 _20658_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _23012_/Q _22979_/Q _14700_/C vssd1 vssd1 vccd1 vccd1 _14700_/X sky130_fd_sc_hd__and3_4
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_62 _21212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_73 _21077_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11912_ _12087_/A _13778_/A _11911_/X _12110_/S vssd1 vssd1 vccd1 vccd1 _13340_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_46_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_84 _11483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15680_ _13629_/A _14942_/X _15679_/X vssd1 vssd1 vccd1 vccd1 _15680_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_79_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12892_ _11196_/A _12667_/X _11402_/A _12891_/Y vssd1 vssd1 vccd1 vccd1 _13493_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_95 _20303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _15292_/S _14629_/Y _14630_/X vssd1 vssd1 vccd1 vccd1 _14632_/B sky130_fd_sc_hd__a21o_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11843_ _11843_/A vssd1 vssd1 vccd1 vccd1 _11844_/A sky130_fd_sc_hd__buf_4
X_23829_ _23871_/CLK _23829_/D vssd1 vssd1 vccd1 vccd1 _23829_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _22596_/Q input213/X _17358_/S vssd1 vssd1 vccd1 vccd1 _17351_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _14534_/X _22261_/Q _14985_/S vssd1 vssd1 vccd1 vccd1 _14563_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11774_ _11774_/A _11774_/B vssd1 vssd1 vccd1 vccd1 _11774_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _22322_/Q _16300_/X _16301_/S vssd1 vssd1 vccd1 vccd1 _16302_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13513_ _13514_/A _13514_/B vssd1 vssd1 vccd1 vccd1 _13513_/X sky130_fd_sc_hd__and2_1
X_17281_ _21077_/A _17280_/X _17291_/S vssd1 vssd1 vccd1 vccd1 _17281_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14493_ _15210_/A vssd1 vssd1 vccd1 vccd1 _14494_/S sky130_fd_sc_hd__clkbuf_4
X_19020_ _19088_/S vssd1 vssd1 vccd1 vccd1 _19029_/S sky130_fd_sc_hd__buf_6
X_16232_ _16232_/A vssd1 vssd1 vccd1 vccd1 _22300_/D sky130_fd_sc_hd__clkbuf_1
X_13444_ _23909_/Q vssd1 vssd1 vccd1 vccd1 _14180_/B sky130_fd_sc_hd__buf_4
XFILLER_16_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_357_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_316_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16163_ _16163_/A vssd1 vssd1 vccd1 vccd1 _22291_/D sky130_fd_sc_hd__clkbuf_1
X_13375_ _13375_/A _13375_/B _13943_/A vssd1 vssd1 vccd1 vccd1 _13376_/B sky130_fd_sc_hd__or3b_1
XFILLER_155_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15114_ input139/X input168/X _15114_/S vssd1 vssd1 vccd1 vccd1 _15114_/X sky130_fd_sc_hd__mux2_8
XFILLER_318_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12326_ _22266_/Q _23082_/Q _23498_/Q _22427_/Q _12324_/X _12325_/X vssd1 vssd1 vccd1
+ vccd1 _12327_/B sky130_fd_sc_hd__mux4_1
X_16094_ _13410_/C _15079_/B _16093_/Y vssd1 vssd1 vccd1 vccd1 _16094_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_336_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_330_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19922_ _23591_/Q _19922_/B _23589_/Q _19922_/D vssd1 vssd1 vccd1 vccd1 _19927_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_303_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15045_ _16198_/S vssd1 vssd1 vccd1 vccd1 _15284_/S sky130_fd_sc_hd__buf_6
XFILLER_141_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12257_ _23467_/Q _23563_/Q _22527_/Q _22331_/Q _11414_/A _12199_/X vssd1 vssd1 vccd1
+ vccd1 _12257_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11208_ _11418_/A vssd1 vssd1 vccd1 vccd1 _11208_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_214_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12188_ _23308_/Q _23276_/Q _23244_/Q _23532_/Q _11700_/A _11565_/A vssd1 vssd1 vccd1
+ vccd1 _12189_/B sky130_fd_sc_hd__mux4_2
X_19853_ _19853_/A vssd1 vssd1 vccd1 vccd1 _23560_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_269_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_311_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18804_ _18804_/A vssd1 vssd1 vccd1 vccd1 _18804_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_352_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11139_ _11834_/A vssd1 vssd1 vccd1 vccd1 _11774_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16996_ _16996_/A vssd1 vssd1 vccd1 vccd1 _16996_/X sky130_fd_sc_hd__clkbuf_2
X_19784_ _19841_/S vssd1 vssd1 vccd1 vccd1 _19793_/S sky130_fd_sc_hd__buf_4
XFILLER_110_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18735_ _16867_/X _23093_/Q _18741_/S vssd1 vssd1 vccd1 vccd1 _18736_/A sky130_fd_sc_hd__mux2_1
XFILLER_352_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15947_ _13408_/Y _13575_/B _16053_/S vssd1 vssd1 vccd1 vccd1 _15947_/X sky130_fd_sc_hd__mux2_1
XTAP_5280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18666_ _18666_/A vssd1 vssd1 vccd1 vccd1 _23062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15878_ _23676_/Q _16021_/B vssd1 vssd1 vccd1 vccd1 _15878_/X sky130_fd_sc_hd__or2_1
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17617_ _18843_/A vssd1 vssd1 vccd1 vccd1 _17617_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14829_ _14829_/A vssd1 vssd1 vccd1 vccd1 _14829_/Y sky130_fd_sc_hd__inv_2
X_18597_ _16876_/X _23032_/Q _18597_/S vssd1 vssd1 vccd1 vccd1 _18598_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17548_ _22678_/Q _17544_/X _17560_/S vssd1 vssd1 vccd1 vccd1 _17549_/A sky130_fd_sc_hd__mux2_1
XFILLER_297_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17479_ _22648_/Q _16214_/X _17483_/S vssd1 vssd1 vccd1 vccd1 _17480_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19218_ _19217_/X _23285_/Q _19227_/S vssd1 vssd1 vccd1 vccd1 _19219_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20490_ _20759_/A _20428_/A _20489_/X _20483_/X vssd1 vssd1 vccd1 vccd1 _23715_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_319_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_301_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19149_ _23262_/Q _18852_/X _19157_/S vssd1 vssd1 vccd1 vccd1 _19150_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22160_ _22161_/A _22161_/B vssd1 vssd1 vccd1 vccd1 _22177_/A sky130_fd_sc_hd__nand2_1
XFILLER_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21111_ _21124_/A vssd1 vssd1 vccd1 vccd1 _21111_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_62_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23349_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22091_ _22116_/B _22091_/B vssd1 vssd1 vccd1 vccd1 _22091_/Y sky130_fd_sc_hd__nor2_1
XTAP_6909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_303_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21042_ _23831_/Q _20993_/X _21041_/Y _21037_/X vssd1 vssd1 vccd1 vccd1 _23831_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_287_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22993_ _23424_/CLK _22993_/D vssd1 vssd1 vccd1 vccd1 _22993_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_243_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21944_ _23833_/Q _23767_/Q vssd1 vssd1 vccd1 vccd1 _21944_/X sky130_fd_sc_hd__or2_1
XFILLER_83_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21875_ _21933_/A vssd1 vssd1 vccd1 vccd1 _21879_/A sky130_fd_sc_hd__inv_2
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23614_ _23637_/CLK _23614_/D vssd1 vssd1 vccd1 vccd1 _23614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20826_ _20826_/A vssd1 vssd1 vccd1 vccd1 _23762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23545_ _23545_/CLK _23545_/D vssd1 vssd1 vccd1 vccd1 _23545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20757_ _20757_/A _20757_/B _20757_/C vssd1 vssd1 vccd1 vccd1 _20757_/X sky130_fd_sc_hd__or3_1
XFILLER_126_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11490_ _22806_/Q _22774_/Q _22675_/Q _22742_/Q _13255_/S _11418_/A vssd1 vssd1 vccd1
+ vccd1 _11491_/B sky130_fd_sc_hd__mux4_1
XFILLER_345_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23476_ _23542_/CLK _23476_/D vssd1 vssd1 vccd1 vccd1 _23476_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20688_ _17180_/X _20632_/X _20687_/X vssd1 vssd1 vccd1 vccd1 _20689_/C sky130_fd_sc_hd__o21a_2
XFILLER_149_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22427_ _23530_/CLK _22427_/D vssd1 vssd1 vccd1 vccd1 _22427_/Q sky130_fd_sc_hd__dfxtp_1
X_23948__507 vssd1 vssd1 vccd1 vccd1 _23948__507/HI core_wb_adr_o[1] sky130_fd_sc_hd__conb_1
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_313_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13160_ _13149_/A _13159_/X _12816_/A vssd1 vssd1 vccd1 vccd1 _13160_/Y sky130_fd_sc_hd__o21ai_1
X_22358_ _23494_/CLK _22358_/D vssd1 vssd1 vccd1 vccd1 _22358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_298_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_352_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12111_ _12112_/A _12112_/B vssd1 vssd1 vccd1 vccd1 _15460_/A sky130_fd_sc_hd__nor2_1
X_13091_ _13091_/A vssd1 vssd1 vccd1 vccd1 _13206_/A sky130_fd_sc_hd__buf_2
XFILLER_269_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21309_ _21560_/A vssd1 vssd1 vccd1 vccd1 _21683_/A sky130_fd_sc_hd__clkbuf_4
X_22289_ _23489_/CLK _22289_/D vssd1 vssd1 vccd1 vccd1 _22289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_317_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12042_ _22307_/Q _23443_/Q _12042_/S vssd1 vssd1 vccd1 vccd1 _12042_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16850_ _16850_/A vssd1 vssd1 vccd1 vccd1 _22531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15801_ _15801_/A _15801_/B vssd1 vssd1 vccd1 vccd1 _15801_/X sky130_fd_sc_hd__or2_1
XFILLER_266_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16781_ _16795_/A _16781_/B vssd1 vssd1 vccd1 vccd1 _16782_/A sky130_fd_sc_hd__or2_1
XFILLER_172_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13993_ _13993_/A vssd1 vssd1 vccd1 vccd1 _14074_/B sky130_fd_sc_hd__clkbuf_2
X_18520_ _18520_/A vssd1 vssd1 vccd1 vccd1 _18520_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_219_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15732_ _23832_/Q _14906_/A _15728_/X _15731_/X _14610_/A vssd1 vssd1 vccd1 vccd1
+ _15732_/X sky130_fd_sc_hd__a221o_2
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ _12993_/A _12944_/B vssd1 vssd1 vccd1 vccd1 _12944_/X sky130_fd_sc_hd__or2_1
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _18480_/A vssd1 vssd1 vccd1 vccd1 _18451_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_234_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ _15672_/A vssd1 vssd1 vccd1 vccd1 _15663_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12875_ _13195_/A _12872_/X _12874_/X vssd1 vssd1 vccd1 vccd1 _12875_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _22614_/Q _16200_/X _17410_/S vssd1 vssd1 vccd1 vccd1 _17403_/A sky130_fd_sc_hd__mux2_1
XFILLER_261_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14614_ _23686_/Q _14494_/S _14613_/X vssd1 vssd1 vccd1 vccd1 _14614_/X sky130_fd_sc_hd__o21a_2
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _15207_/X _18384_/C _18381_/Y vssd1 vssd1 vccd1 vccd1 _22954_/D sky130_fd_sc_hd__o21a_1
X_11826_ _11826_/A _11826_/B _11826_/C vssd1 vssd1 vccd1 vccd1 _11826_/X sky130_fd_sc_hd__or3_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _23669_/Q _16102_/B vssd1 vssd1 vccd1 vccd1 _15594_/X sky130_fd_sc_hd__or2_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_324_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17333_ _22589_/Q input206/X _17335_/S vssd1 vssd1 vccd1 vccd1 _17334_/A sky130_fd_sc_hd__mux2_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _17471_/A _17471_/B _19090_/A vssd1 vssd1 vccd1 vccd1 _19699_/A sky130_fd_sc_hd__or3_1
XFILLER_14_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11757_ _11986_/A _11757_/B vssd1 vssd1 vccd1 vccd1 _11757_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_347_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17264_ _17242_/X _17256_/X _17263_/X _17237_/X vssd1 vssd1 vccd1 vccd1 _17264_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_202_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14476_ _14912_/A vssd1 vssd1 vccd1 vccd1 _15596_/A sky130_fd_sc_hd__buf_4
XFILLER_347_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11688_ _12110_/S vssd1 vssd1 vccd1 vccd1 _12739_/A sky130_fd_sc_hd__clkbuf_2
X_19003_ _19003_/A vssd1 vssd1 vccd1 vccd1 _19012_/S sky130_fd_sc_hd__buf_6
XFILLER_347_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16215_ _22295_/Q _16214_/X _16221_/S vssd1 vssd1 vccd1 vccd1 _16216_/A sky130_fd_sc_hd__mux2_1
X_13427_ _13427_/A _13427_/B _14792_/A vssd1 vssd1 vccd1 vccd1 _13427_/X sky130_fd_sc_hd__or3_1
X_17195_ _17262_/A vssd1 vssd1 vccd1 vccd1 _17195_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_350_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16146_ _14518_/A _16134_/X _16145_/X vssd1 vssd1 vccd1 vccd1 _17307_/A sky130_fd_sc_hd__o21ai_4
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ _13897_/A _13358_/B vssd1 vssd1 vccd1 vccd1 _14759_/A sky130_fd_sc_hd__xor2_1
XFILLER_304_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12309_ _12196_/X _12308_/X _11706_/A vssd1 vssd1 vccd1 vccd1 _12309_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_303_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16077_ _22165_/A _16077_/B vssd1 vssd1 vccd1 vccd1 _16078_/B sky130_fd_sc_hd__nor2_1
XFILLER_115_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13289_ _11343_/A _13288_/X _11288_/X vssd1 vssd1 vccd1 vccd1 _13289_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_216_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_331_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19905_ _16294_/X _23584_/Q _19909_/S vssd1 vssd1 vccd1 vccd1 _19906_/A sky130_fd_sc_hd__mux2_1
X_15028_ input155/X _13650_/A _14967_/S input120/X _14235_/X vssd1 vssd1 vccd1 vccd1
+ _15028_/X sky130_fd_sc_hd__a221o_4
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_300_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19836_ _19836_/A vssd1 vssd1 vccd1 vccd1 _23553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_300_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19767_ _19261_/X _23523_/Q _19769_/S vssd1 vssd1 vccd1 vccd1 _19768_/A sky130_fd_sc_hd__mux2_1
Xinput3 coreIndex[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_4
X_16979_ _21301_/B _16978_/Y _16932_/A _16947_/X vssd1 vssd1 vccd1 vccd1 _16979_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_244_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18718_ _18718_/A vssd1 vssd1 vccd1 vccd1 _23085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19698_ _19698_/A vssd1 vssd1 vccd1 vccd1 _23492_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_180_wb_clk_i _23931_/CLK vssd1 vssd1 vccd1 vccd1 _23936_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18649_ _18695_/S vssd1 vssd1 vccd1 vccd1 _18658_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_224_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_358_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21660_ _22129_/A vssd1 vssd1 vccd1 vccd1 _21660_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_40_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20611_ _14548_/X _20564_/X _20598_/X vssd1 vssd1 vccd1 vccd1 _20611_/X sky130_fd_sc_hd__a21o_1
XFILLER_221_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21591_ _23919_/Q _21591_/B vssd1 vssd1 vccd1 vccd1 _21591_/X sky130_fd_sc_hd__or2_1
XFILLER_33_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_338_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_327_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23330_ _23426_/CLK _23330_/D vssd1 vssd1 vccd1 vccd1 _23330_/Q sky130_fd_sc_hd__dfxtp_1
X_20542_ _20628_/A vssd1 vssd1 vccd1 vccd1 _20542_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23261_ _23549_/CLK _23261_/D vssd1 vssd1 vccd1 vccd1 _23261_/Q sky130_fd_sc_hd__dfxtp_1
X_20473_ _20713_/A _20467_/X _20471_/X _20472_/X vssd1 vssd1 vccd1 vccd1 _23707_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22212_ _22187_/A _22189_/B _22187_/B vssd1 vssd1 vccd1 vccd1 _22213_/B sky130_fd_sc_hd__a21bo_1
XFILLER_106_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23192_ _23354_/CLK _23192_/D vssd1 vssd1 vccd1 vccd1 _23192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_335_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_350_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22143_ _22168_/A _22142_/B _22142_/C vssd1 vssd1 vccd1 vccd1 _22143_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_156_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput340 _13795_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[17] sky130_fd_sc_hd__buf_2
XFILLER_350_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput351 _13856_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[27] sky130_fd_sc_hd__buf_2
XFILLER_105_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput362 _13742_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[8] sky130_fd_sc_hd__buf_2
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput373 _13651_/Y vssd1 vssd1 vccd1 vccd1 csb1[1] sky130_fd_sc_hd__buf_2
X_22074_ _13165_/Y _21867_/X _22073_/X _21865_/X vssd1 vssd1 vccd1 vccd1 _22075_/B
+ sky130_fd_sc_hd__a22o_2
XTAP_6739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput384 _14047_/X vssd1 vssd1 vccd1 vccd1 din0[19] sky130_fd_sc_hd__buf_2
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput395 _14067_/X vssd1 vssd1 vccd1 vccd1 din0[29] sky130_fd_sc_hd__buf_2
XFILLER_248_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21025_ _21025_/A _21043_/B vssd1 vssd1 vccd1 vccd1 _21025_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_290_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_347_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22976_ _22977_/CLK _22976_/D vssd1 vssd1 vccd1 vccd1 _22976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21927_ _13020_/Y _21841_/A _15753_/Y _21842_/X vssd1 vssd1 vccd1 vccd1 _21927_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12660_/A _12660_/B _12660_/C vssd1 vssd1 vccd1 vccd1 _12661_/B sky130_fd_sc_hd__nor3_4
XFILLER_231_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21858_ _21828_/A _21827_/A _21826_/Y vssd1 vssd1 vccd1 vccd1 _21858_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11611_/A vssd1 vssd1 vccd1 vccd1 _11621_/A sky130_fd_sc_hd__clkbuf_4
X_20809_ _20881_/A vssd1 vssd1 vccd1 vccd1 _20825_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12591_ _22458_/Q _22618_/Q _22297_/Q _23433_/Q _12314_/X _12325_/X vssd1 vssd1 vccd1
+ vccd1 _12591_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21789_ _21763_/B _21765_/B _21763_/A vssd1 vssd1 vccd1 vccd1 _21793_/A sky130_fd_sc_hd__a21bo_1
XFILLER_230_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14330_ _12171_/B _12636_/X _14330_/S vssd1 vssd1 vccd1 vccd1 _14330_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11542_ _13114_/A vssd1 vssd1 vccd1 vccd1 _11543_/A sky130_fd_sc_hd__buf_4
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23528_ _23528_/CLK _23528_/D vssd1 vssd1 vccd1 vccd1 _23528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_345_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_357_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14261_ _14835_/A _13367_/C _14254_/X _13464_/B _14260_/X vssd1 vssd1 vccd1 vccd1
+ _14261_/X sky130_fd_sc_hd__a221o_1
X_23459_ _23459_/CLK _23459_/D vssd1 vssd1 vccd1 vccd1 _23459_/Q sky130_fd_sc_hd__dfxtp_1
X_11473_ _15630_/A _11472_/X _15671_/A vssd1 vssd1 vccd1 vccd1 _11473_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_109_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16000_ _15995_/Y _15997_/X _15999_/X _14690_/A vssd1 vssd1 vccd1 vccd1 _16000_/X
+ sky130_fd_sc_hd__a31o_2
X_13212_ _13212_/A _13836_/A vssd1 vssd1 vccd1 vccd1 _13212_/Y sky130_fd_sc_hd__nand2_1
XFILLER_332_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14192_ _14800_/A _14192_/B vssd1 vssd1 vccd1 vccd1 _14199_/B sky130_fd_sc_hd__and2_1
XFILLER_325_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13143_ _13199_/A _13143_/B vssd1 vssd1 vccd1 vccd1 _13143_/Y sky130_fd_sc_hd__nor2_1
XFILLER_298_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_341_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_297_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17951_ _17983_/A vssd1 vssd1 vccd1 vccd1 _17951_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_301_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13074_ _22481_/Q _22641_/Q _22320_/Q _23456_/Q _11311_/A _11527_/X vssd1 vssd1 vccd1
+ vccd1 _13074_/X sky130_fd_sc_hd__mux4_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16902_ _19252_/A vssd1 vssd1 vccd1 vccd1 _16902_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_250_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12025_ _12025_/A vssd1 vssd1 vccd1 vccd1 _12025_/X sky130_fd_sc_hd__buf_6
X_17882_ _22812_/Q input250/X _17882_/S vssd1 vssd1 vccd1 vccd1 _17883_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_333_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19621_ _23458_/Q _19258_/A _19621_/S vssd1 vssd1 vccd1 vccd1 _19622_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_293_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16833_ _16831_/X _22526_/Q _16845_/S vssd1 vssd1 vccd1 vccd1 _16834_/A sky130_fd_sc_hd__mux2_1
XFILLER_281_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_293_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16764_ _16764_/A vssd1 vssd1 vccd1 vccd1 _22506_/D sky130_fd_sc_hd__clkbuf_1
X_19552_ _19552_/A vssd1 vssd1 vccd1 vccd1 _23427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13976_ _13976_/A vssd1 vssd1 vccd1 vccd1 _13976_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_207_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18503_ _18516_/A vssd1 vssd1 vccd1 vccd1 _18503_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15715_ _21916_/A _21868_/B vssd1 vssd1 vccd1 vccd1 _15716_/B sky130_fd_sc_hd__nor2_1
X_12927_ _22377_/Q _22409_/Q _22698_/Q _23065_/Q _12680_/X _12637_/X vssd1 vssd1 vccd1
+ vccd1 _12927_/X sky130_fd_sc_hd__mux4_1
X_19483_ _19627_/A _19483_/B vssd1 vssd1 vccd1 vccd1 _19540_/A sky130_fd_sc_hd__or2_4
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16695_ _16704_/A _16695_/B vssd1 vssd1 vccd1 vccd1 _16696_/A sky130_fd_sc_hd__or2_1
XFILLER_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18434_ _18435_/A _18435_/C _22973_/Q vssd1 vssd1 vccd1 vccd1 _18436_/B sky130_fd_sc_hd__a21oi_1
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15646_ _23670_/Q _15985_/B vssd1 vssd1 vccd1 vccd1 _15646_/X sky130_fd_sc_hd__or2_1
X_12858_ _12953_/A _12857_/X _12707_/A vssd1 vssd1 vccd1 vccd1 _12858_/X sky130_fd_sc_hd__o21a_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18365_ _14729_/X _18366_/C _22949_/Q vssd1 vssd1 vccd1 vccd1 _18367_/B sky130_fd_sc_hd__a21oi_1
X_11809_ _22464_/Q _22624_/Q _22303_/Q _23439_/Q _11745_/A _11742_/A vssd1 vssd1 vccd1
+ vccd1 _11809_/X sky130_fd_sc_hd__mux4_1
XFILLER_187_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15577_ _13737_/A _15533_/Y _15576_/Y vssd1 vssd1 vccd1 vccd1 _15578_/A sky130_fd_sc_hd__a21oi_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _12906_/A _12789_/B vssd1 vssd1 vccd1 vccd1 _12789_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _23492_/Q _17016_/X _17017_/X _17042_/A _16179_/X vssd1 vssd1 vccd1 vccd1
+ _17316_/X sky130_fd_sc_hd__a32o_1
X_14528_ _14557_/A vssd1 vssd1 vccd1 vccd1 _15519_/A sky130_fd_sc_hd__buf_4
XFILLER_187_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18296_ _18296_/A _22925_/Q _18296_/C vssd1 vssd1 vccd1 vccd1 _18297_/C sky130_fd_sc_hd__and3_1
XFILLER_174_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_358_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_348_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_308_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17247_ _23485_/Q _17230_/X _17231_/X _17181_/X _15914_/X vssd1 vssd1 vccd1 vccd1
+ _17247_/X sky130_fd_sc_hd__a32o_1
XFILLER_335_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14459_ _14506_/B _14465_/C vssd1 vssd1 vccd1 vccd1 _20989_/B sky130_fd_sc_hd__or2_2
XFILLER_294_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17178_ _22570_/Q _17141_/X _17131_/X _17177_/X vssd1 vssd1 vccd1 vccd1 _22570_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_227_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16129_ _15082_/X _16128_/X _13307_/A vssd1 vssd1 vccd1 vccd1 _16129_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_304_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_288_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_297_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_300_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19819_ _19819_/A vssd1 vssd1 vccd1 vccd1 _23545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_257_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22830_ _22830_/CLK _22830_/D vssd1 vssd1 vccd1 vccd1 _22830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22761_ _23446_/CLK _22761_/D vssd1 vssd1 vccd1 vccd1 _22761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21712_ _20268_/Y _21711_/X _21712_/S vssd1 vssd1 vccd1 vccd1 _21712_/X sky130_fd_sc_hd__mux2_2
XFILLER_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22692_ _23580_/CLK _22692_/D vssd1 vssd1 vccd1 vccd1 _22692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21643_ _21922_/A _21643_/B vssd1 vssd1 vccd1 vccd1 _21643_/Y sky130_fd_sc_hd__nand2_1
XFILLER_178_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21574_ _21574_/A _21574_/B vssd1 vssd1 vccd1 vccd1 _21574_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_193_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23313_ _23537_/CLK _23313_/D vssd1 vssd1 vccd1 vccd1 _23313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20525_ _20525_/A _20525_/B _20525_/C _20525_/D vssd1 vssd1 vccd1 vccd1 _20526_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_326_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_342_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_314_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23244_ _23950_/A _23244_/D vssd1 vssd1 vccd1 vccd1 _23244_/Q sky130_fd_sc_hd__dfxtp_1
X_20456_ _20675_/A _20447_/X _20455_/X _20445_/X vssd1 vssd1 vccd1 vccd1 _23701_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20387_ _20387_/A _20387_/B vssd1 vssd1 vccd1 vccd1 _20389_/B sky130_fd_sc_hd__or2_1
X_23175_ _23367_/CLK _23175_/D vssd1 vssd1 vccd1 vccd1 _23175_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_7226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22126_ _22139_/A _22044_/X _22125_/X _22048_/X vssd1 vssd1 vccd1 vccd1 _22127_/B
+ sky130_fd_sc_hd__o22a_2
XTAP_7259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_322_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22057_ _22057_/A _22057_/B vssd1 vssd1 vccd1 vccd1 _22059_/A sky130_fd_sc_hd__nor2_1
XFILLER_48_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21008_ _21008_/A vssd1 vssd1 vccd1 vccd1 _21008_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_290_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13830_ _13874_/A _13830_/B _13874_/C vssd1 vssd1 vccd1 vccd1 _13830_/Y sky130_fd_sc_hd__nand3_1
XFILLER_262_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13761_ _13893_/A vssd1 vssd1 vccd1 vccd1 _13807_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_290_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22959_ _22961_/CLK _22959_/D vssd1 vssd1 vccd1 vccd1 _22959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_209 _15596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15500_ _22928_/Q _14752_/A _14753_/A _15501_/A vssd1 vssd1 vccd1 vccd1 _15500_/X
+ sky130_fd_sc_hd__o22a_1
X_12712_ _12953_/A _12712_/B vssd1 vssd1 vccd1 vccd1 _12712_/X sky130_fd_sc_hd__or2_1
XFILLER_280_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16480_ _15283_/X _22398_/Q _16480_/S vssd1 vssd1 vccd1 vccd1 _16481_/A sky130_fd_sc_hd__mux2_1
X_13692_ _13692_/A vssd1 vssd1 vccd1 vccd1 _13934_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_243_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15431_ _15529_/C _15431_/B vssd1 vssd1 vccd1 vccd1 _15431_/X sky130_fd_sc_hd__or2_4
XFILLER_43_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12643_ _12047_/A _12642_/X _11598_/X vssd1 vssd1 vccd1 vccd1 _12643_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_30_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18150_ _18159_/A _18150_/B vssd1 vssd1 vccd1 vccd1 _18151_/A sky130_fd_sc_hd__and2_1
XPHY_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15362_ _14937_/X _15349_/X _15361_/X vssd1 vssd1 vccd1 vccd1 _17103_/A sky130_fd_sc_hd__o21ai_4
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12574_ _11404_/A _12368_/B _13718_/B _13718_/C _12573_/X vssd1 vssd1 vccd1 vccd1
+ _12574_/X sky130_fd_sc_hd__a41o_1
XFILLER_357_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_345_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17101_ _22563_/Q _17091_/X _17083_/X _17100_/X vssd1 vssd1 vccd1 vccd1 _22563_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_12_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14313_ _14313_/A vssd1 vssd1 vccd1 vccd1 _15130_/S sky130_fd_sc_hd__clkbuf_2
X_18081_ _18096_/A vssd1 vssd1 vccd1 vccd1 _18081_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_317_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11525_ _13114_/A vssd1 vssd1 vccd1 vccd1 _11526_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_184_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15293_ _15293_/A vssd1 vssd1 vccd1 vccd1 _15293_/Y sky130_fd_sc_hd__inv_2
XFILLER_346_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_317_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17032_ _13440_/C _17030_/X _17144_/A vssd1 vssd1 vccd1 vccd1 _17032_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14244_ _14218_/X _15189_/A _15186_/A _13829_/B _14243_/Y vssd1 vssd1 vccd1 vccd1
+ _14244_/X sky130_fd_sc_hd__o221a_1
XFILLER_171_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11456_ _11745_/A vssd1 vssd1 vccd1 vccd1 _11457_/C sky130_fd_sc_hd__buf_6
XFILLER_172_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14175_ _14175_/A _14175_/B vssd1 vssd1 vccd1 vccd1 _14175_/Y sky130_fd_sc_hd__nor2_4
XFILLER_341_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_298_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11387_ _12157_/S vssd1 vssd1 vccd1 vccd1 _12913_/S sky130_fd_sc_hd__buf_6
XFILLER_152_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13126_ _13180_/A _13126_/B vssd1 vssd1 vccd1 vccd1 _13126_/Y sky130_fd_sc_hd__nor2_1
XFILLER_341_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18983_ _18983_/A vssd1 vssd1 vccd1 vccd1 _23188_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_119_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23632_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17934_ _22822_/Q _17922_/X _17918_/X input263/X _17933_/X vssd1 vssd1 vccd1 vccd1
+ _17934_/X sky130_fd_sc_hd__a221o_1
X_13057_ _23906_/Q _11486_/B _11403_/X _13056_/Y vssd1 vssd1 vccd1 vccd1 _13249_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12008_ _12024_/A vssd1 vssd1 vccd1 vccd1 _12008_/X sky130_fd_sc_hd__buf_6
XFILLER_121_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17865_ _17865_/A vssd1 vssd1 vccd1 vccd1 _22803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19604_ _23450_/Q _19233_/A _19610_/S vssd1 vssd1 vccd1 vccd1 _19605_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16816_ _16915_/S vssd1 vssd1 vccd1 vccd1 _16829_/S sky130_fd_sc_hd__buf_6
XFILLER_93_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17796_ _22773_/Q _17636_/X _17798_/S vssd1 vssd1 vccd1 vccd1 _17797_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19535_ _19535_/A vssd1 vssd1 vccd1 vccd1 _23419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_282_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13959_ _21289_/A vssd1 vssd1 vccd1 vccd1 _21081_/A sky130_fd_sc_hd__buf_4
XFILLER_35_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16747_ _16783_/A vssd1 vssd1 vccd1 vccd1 _16747_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_281_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19466_ _23389_/Q _18849_/X _19466_/S vssd1 vssd1 vccd1 vccd1 _19467_/A sky130_fd_sc_hd__mux2_1
X_16678_ _16678_/A vssd1 vssd1 vccd1 vccd1 _22485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18417_ _18418_/A _18418_/C _22967_/Q vssd1 vssd1 vccd1 vccd1 _18419_/B sky130_fd_sc_hd__a21oi_1
XFILLER_34_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15629_ _21890_/B vssd1 vssd1 vccd1 vccd1 _21861_/A sky130_fd_sc_hd__buf_4
X_19397_ _23358_/Q _18852_/X _19405_/S vssd1 vssd1 vccd1 vccd1 _19398_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18348_ _16059_/X _18349_/C _22943_/Q vssd1 vssd1 vccd1 vccd1 _18350_/B sky130_fd_sc_hd__a21oi_1
XFILLER_188_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18279_ _22918_/Q _22919_/Q _22920_/Q _18279_/D vssd1 vssd1 vccd1 vccd1 _18288_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_296_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_352_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20310_ _20272_/X _20680_/A _20309_/X _20285_/X vssd1 vssd1 vccd1 vccd1 _23670_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21290_ _22587_/Q _22588_/Q vssd1 vssd1 vccd1 vccd1 _21290_/X sky130_fd_sc_hd__or2_2
XFILLER_163_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput50 dout0[16] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_2
XFILLER_351_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput61 dout0[26] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_2
XFILLER_337_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput72 dout0[36] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__clkbuf_1
XFILLER_289_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput83 dout0[46] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__clkbuf_1
X_20241_ _21596_/A _20340_/B vssd1 vssd1 vccd1 vccd1 _20243_/B sky130_fd_sc_hd__nor2_1
Xinput94 dout0[56] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__clkbuf_1
XFILLER_351_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_320_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_320_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20172_ _14619_/X _20169_/X _20171_/X vssd1 vssd1 vccd1 vccd1 _20172_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23931_ _23931_/CLK _23931_/D vssd1 vssd1 vccd1 vccd1 _23931_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_285_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23862_ _23862_/CLK _23862_/D vssd1 vssd1 vccd1 vccd1 _23862_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22813_ _23551_/CLK _22813_/D vssd1 vssd1 vccd1 vccd1 _22813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23793_ _23861_/CLK _23793_/D vssd1 vssd1 vccd1 vccd1 _23793_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_213_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22744_ _23588_/CLK _22744_/D vssd1 vssd1 vccd1 vccd1 _22744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_305_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22675_ _23586_/CLK _22675_/D vssd1 vssd1 vccd1 vccd1 _22675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_279_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21626_ _21613_/X _21625_/Y _21560_/X _23791_/Q vssd1 vssd1 vccd1 vccd1 _21626_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_139_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_327_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21557_ _21570_/A _21867_/A _21554_/Y _21556_/X vssd1 vssd1 vccd1 vccd1 _21605_/C
+ sky130_fd_sc_hd__a22o_2
XFILLER_328_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11310_ _11517_/A vssd1 vssd1 vccd1 vccd1 _11311_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_354_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20508_ _23705_/Q _20508_/B _20508_/C vssd1 vssd1 vccd1 vccd1 _20509_/D sky130_fd_sc_hd__and3_1
XFILLER_315_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12290_ _23210_/Q _23178_/Q _23146_/Q _23114_/Q _11700_/A _11840_/X vssd1 vssd1 vccd1
+ vccd1 _12291_/B sky130_fd_sc_hd__mux4_1
XFILLER_193_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21488_ _23787_/Q _21814_/B _21487_/Y _21346_/X vssd1 vssd1 vccd1 vccd1 _21489_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_308_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23227_ _23419_/CLK _23227_/D vssd1 vssd1 vccd1 vccd1 _23227_/Q sky130_fd_sc_hd__dfxtp_1
X_11241_ _11241_/A vssd1 vssd1 vccd1 vccd1 _11242_/A sky130_fd_sc_hd__buf_4
XTAP_7001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20439_ _20622_/A _20428_/X _20438_/X _20433_/X vssd1 vssd1 vccd1 vccd1 _23694_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_7012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23158_ _23543_/CLK _23158_/D vssd1 vssd1 vccd1 vccd1 _23158_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11172_ _13259_/A _11172_/B vssd1 vssd1 vccd1 vccd1 _11172_/Y sky130_fd_sc_hd__nor2_1
XFILLER_162_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22109_ _22109_/A _22108_/Y vssd1 vssd1 vccd1 vccd1 _22110_/B sky130_fd_sc_hd__or2b_1
XTAP_7089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15980_ _22972_/Q vssd1 vssd1 vccd1 vccd1 _18435_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_6355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23089_ _23409_/CLK _23089_/D vssd1 vssd1 vccd1 vccd1 _23089_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14931_ _14931_/A vssd1 vssd1 vccd1 vccd1 _15000_/A sky130_fd_sc_hd__buf_2
XFILLER_94_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17650_ _21351_/B _17653_/B vssd1 vssd1 vccd1 vccd1 _17650_/Y sky130_fd_sc_hd__nand2_1
X_14862_ _14839_/X _16057_/B _14861_/X _14632_/A vssd1 vssd1 vccd1 vccd1 _14862_/Y
+ sky130_fd_sc_hd__o22ai_4
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ _16124_/X _22451_/Q _16601_/S vssd1 vssd1 vccd1 vccd1 _16602_/A sky130_fd_sc_hd__mux2_1
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13813_ _13813_/A vssd1 vssd1 vccd1 vccd1 _13813_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17581_ _17581_/A vssd1 vssd1 vccd1 vccd1 _22688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_251_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14793_ _14793_/A vssd1 vssd1 vccd1 vccd1 _14942_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_291_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19320_ _19239_/X _23324_/Q _19322_/S vssd1 vssd1 vccd1 vccd1 _19321_/A sky130_fd_sc_hd__mux2_1
X_16532_ _18277_/A vssd1 vssd1 vccd1 vccd1 _18476_/A sky130_fd_sc_hd__buf_2
XFILLER_244_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13744_ _13893_/A vssd1 vssd1 vccd1 vccd1 _13974_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_204_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19251_ _19251_/A vssd1 vssd1 vccd1 vccd1 _23295_/D sky130_fd_sc_hd__clkbuf_1
X_16463_ _14706_/X _22390_/Q _16469_/S vssd1 vssd1 vccd1 vccd1 _16464_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13675_ _17219_/S vssd1 vssd1 vccd1 vccd1 _17029_/S sky130_fd_sc_hd__buf_8
X_18202_ _18242_/A vssd1 vssd1 vccd1 vccd1 _18202_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15414_ _14807_/A _15391_/A _15574_/A vssd1 vssd1 vccd1 vccd1 _15414_/X sky130_fd_sc_hd__o21a_1
X_12626_ _12958_/A _12626_/B vssd1 vssd1 vccd1 vccd1 _12626_/Y sky130_fd_sc_hd__nor2_1
XPHY_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19182_ _19265_/S vssd1 vssd1 vccd1 vccd1 _19195_/S sky130_fd_sc_hd__buf_4
XPHY_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16394_ _14893_/X _22360_/Q _16396_/S vssd1 vssd1 vccd1 vccd1 _16395_/A sky130_fd_sc_hd__mux2_1
XPHY_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18133_ _18116_/A _18166_/B _22882_/Q vssd1 vssd1 vccd1 vccd1 _18133_/X sky130_fd_sc_hd__a21o_1
XPHY_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15345_ _15345_/A _15345_/B vssd1 vssd1 vccd1 vccd1 _15345_/Y sky130_fd_sc_hd__nor2_1
XFILLER_318_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12557_ _13455_/A _23433_/Q _12556_/X _11703_/A vssd1 vssd1 vccd1 vccd1 _12557_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18064_ hold7/A _18052_/X _18053_/X _22992_/Q _18054_/X vssd1 vssd1 vccd1 vccd1 _18064_/X
+ sky130_fd_sc_hd__a221o_1
X_11508_ _11497_/A _11507_/X _11236_/A vssd1 vssd1 vccd1 vccd1 _11508_/Y sky130_fd_sc_hd__o21ai_1
X_15276_ _15316_/B _15276_/B vssd1 vssd1 vccd1 vccd1 _15277_/B sky130_fd_sc_hd__or2_2
XFILLER_334_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12488_ _22778_/Q _22746_/Q _22647_/Q _22714_/Q _11919_/A _12476_/X vssd1 vssd1 vccd1
+ vccd1 _12489_/B sky130_fd_sc_hd__mux4_2
XFILLER_355_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17015_ input71/X input76/X _17029_/S vssd1 vssd1 vccd1 vccd1 _17015_/X sky130_fd_sc_hd__mux2_8
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14227_ _15057_/S vssd1 vssd1 vccd1 vccd1 _15030_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_172_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11439_ _13032_/S vssd1 vssd1 vccd1 vccd1 _13255_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_125_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_314_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14158_ _14421_/S _21294_/A vssd1 vssd1 vccd1 vccd1 _16962_/A sky130_fd_sc_hd__nand2_2
XFILLER_99_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_298_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13109_ _11219_/A _13099_/X _13108_/X _13210_/A vssd1 vssd1 vccd1 vccd1 _13110_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_98_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14089_ _14089_/A _14089_/B vssd1 vssd1 vccd1 vccd1 _14089_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18966_ _16841_/X _23181_/Q _18968_/S vssd1 vssd1 vccd1 vccd1 _18967_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17917_ _22818_/Q _17914_/X _17916_/X _17912_/X vssd1 vssd1 vccd1 vccd1 _22818_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_255_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18897_ _18897_/A vssd1 vssd1 vccd1 vccd1 _23150_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_254_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17848_ _22796_/Q _17607_/X _17848_/S vssd1 vssd1 vccd1 vccd1 _17849_/A sky130_fd_sc_hd__mux2_1
XFILLER_254_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_87_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23451_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17779_ _22765_/Q _17610_/X _17787_/S vssd1 vssd1 vccd1 vccd1 _17780_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19518_ _19540_/A vssd1 vssd1 vccd1 vccd1 _19527_/S sky130_fd_sc_hd__buf_4
XFILLER_281_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20790_ _20790_/A vssd1 vssd1 vccd1 vccd1 _20806_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_16_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23567_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_223_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_540 _23917_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_551 _14224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19449_ _23381_/Q _18824_/X _19455_/S vssd1 vssd1 vccd1 vccd1 _19450_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_562 _23911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22460_ _23563_/CLK _22460_/D vssd1 vssd1 vccd1 vccd1 _22460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_249_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21411_ _21379_/X _21396_/X _21409_/X _21410_/X vssd1 vssd1 vccd1 vccd1 _21411_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_309_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22391_ _23047_/CLK _22391_/D vssd1 vssd1 vccd1 vccd1 _22391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21342_ _21342_/A _21342_/B vssd1 vssd1 vccd1 vccd1 _21344_/B sky130_fd_sc_hd__xor2_1
XFILLER_190_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_352_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21273_ _21078_/A _21242_/X _21272_/Y _21270_/X vssd1 vssd1 vccd1 vccd1 _23905_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_352_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23012_ _23599_/CLK _23012_/D vssd1 vssd1 vccd1 vccd1 _23012_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20224_ _20213_/X _20604_/A _20223_/X _20203_/X vssd1 vssd1 vccd1 vccd1 _23659_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_320_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20155_ _14520_/B _20154_/X _20152_/X vssd1 vssd1 vccd1 vccd1 _20155_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_277_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_320_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_311_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20086_ _20086_/A _20086_/B _20095_/D vssd1 vssd1 vccd1 vccd1 _23636_/D sky130_fd_sc_hd__nor3_1
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23914_ _23915_/CLK _23914_/D vssd1 vssd1 vccd1 vccd1 _23914_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23845_ _23846_/CLK _23845_/D vssd1 vssd1 vccd1 vccd1 _23845_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _23471_/Q _23567_/Q _22531_/Q _22335_/Q _11708_/S _11613_/A vssd1 vssd1 vccd1
+ vccd1 _11790_/X sky130_fd_sc_hd__mux4_1
X_23776_ _23776_/CLK _23776_/D vssd1 vssd1 vccd1 vccd1 _23776_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20988_ _21008_/A vssd1 vssd1 vccd1 vccd1 _20988_/X sky130_fd_sc_hd__buf_2
XFILLER_300_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22727_ _23580_/CLK _22727_/D vssd1 vssd1 vccd1 vccd1 _22727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_347_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13460_ _23912_/Q vssd1 vssd1 vccd1 vccd1 _16980_/A sky130_fd_sc_hd__buf_4
XFILLER_230_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22658_ _23568_/CLK _22658_/D vssd1 vssd1 vccd1 vccd1 _22658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12411_ _22456_/Q _22616_/Q _22295_/Q _23431_/Q _11647_/A _12269_/X vssd1 vssd1 vccd1
+ vccd1 _12411_/X sky130_fd_sc_hd__mux4_2
X_21609_ _21663_/A _21608_/X _21922_/A vssd1 vssd1 vccd1 vccd1 _21609_/Y sky130_fd_sc_hd__o21ai_1
X_13391_ _13608_/A _13391_/B vssd1 vssd1 vccd1 vccd1 _15635_/A sky130_fd_sc_hd__xnor2_4
XFILLER_138_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_316_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22589_ _22968_/CLK _22589_/D vssd1 vssd1 vccd1 vccd1 _22589_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_159_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_355_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15130_ _14377_/X _15538_/B _15130_/S vssd1 vssd1 vccd1 vccd1 _15131_/A sky130_fd_sc_hd__mux2_1
XFILLER_355_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12342_ _13421_/A _23891_/Q vssd1 vssd1 vccd1 vccd1 _20139_/A sky130_fd_sc_hd__nor2b_4
XFILLER_309_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_342_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15061_ _13738_/A _15483_/A _15485_/A _13789_/A vssd1 vssd1 vccd1 vccd1 _15061_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_142_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12273_ _23211_/Q _23179_/Q _23147_/Q _23115_/Q _11305_/A _11869_/X vssd1 vssd1 vccd1
+ vccd1 _12274_/B sky130_fd_sc_hd__mux4_2
XFILLER_181_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14012_ _14049_/A vssd1 vssd1 vccd1 vccd1 _14012_/X sky130_fd_sc_hd__clkbuf_4
X_11224_ _23428_/Q _23044_/Q _23396_/Q _23364_/Q _11157_/X _11170_/X vssd1 vssd1 vccd1
+ vccd1 _11224_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18820_ _18820_/A vssd1 vssd1 vccd1 vccd1 _18820_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11155_ _13191_/S vssd1 vssd1 vccd1 vccd1 _13190_/S sky130_fd_sc_hd__buf_4
XTAP_6141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18751_ _18751_/A vssd1 vssd1 vccd1 vccd1 _23100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15963_ _14518_/A _15951_/X _15962_/X vssd1 vssd1 vccd1 vccd1 _17258_/A sky130_fd_sc_hd__o21ai_4
XFILLER_237_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11086_ _23882_/Q _23881_/Q _23880_/Q _23879_/Q vssd1 vssd1 vccd1 vccd1 _13775_/B
+ sky130_fd_sc_hd__or4bb_2
XTAP_6196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput240 localMemory_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input240/X sky130_fd_sc_hd__buf_4
XTAP_5462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput251 localMemory_wb_stb_i vssd1 vssd1 vccd1 vccd1 _17326_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_48_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17702_ _22731_/Q _17604_/X _17704_/S vssd1 vssd1 vccd1 vccd1 _17703_/A sky130_fd_sc_hd__mux2_1
XTAP_5473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput262 manufacturerID[8] vssd1 vssd1 vccd1 vccd1 input262/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14914_ _15806_/S vssd1 vssd1 vccd1 vccd1 _15879_/S sky130_fd_sc_hd__buf_4
Xinput273 partID[3] vssd1 vssd1 vccd1 vccd1 input273/X sky130_fd_sc_hd__clkbuf_1
XTAP_5484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18682_ _18682_/A vssd1 vssd1 vccd1 vccd1 _18691_/S sky130_fd_sc_hd__buf_6
XFILLER_208_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15894_ _15864_/X _15672_/X _15892_/X _15893_/X vssd1 vssd1 vccd1 vccd1 _15894_/X
+ sky130_fd_sc_hd__o22a_4
XTAP_5495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput284 wb_rst_i vssd1 vssd1 vccd1 vccd1 _16530_/A sky130_fd_sc_hd__buf_12
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_0_1_wb_clk_i clkbuf_3_0_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_341_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17633_ _18859_/A vssd1 vssd1 vccd1 vccd1 _17633_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_291_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14845_ _14654_/X _14656_/X _14845_/S vssd1 vssd1 vccd1 vccd1 _14845_/X sky130_fd_sc_hd__mux2_2
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_327_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17564_ _22683_/Q _17562_/X _17576_/S vssd1 vssd1 vccd1 vccd1 _17565_/A sky130_fd_sc_hd__mux2_1
X_14776_ _14302_/X _14306_/X _14841_/S vssd1 vssd1 vccd1 vccd1 _14776_/X sky130_fd_sc_hd__mux2_1
X_11988_ _23412_/Q _23028_/Q _23380_/Q _23348_/Q _12029_/A _11676_/A vssd1 vssd1 vccd1
+ vccd1 _11989_/B sky130_fd_sc_hd__mux4_2
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19303_ _19213_/X _23316_/Q _19311_/S vssd1 vssd1 vccd1 vccd1 _19304_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16515_ _16515_/A vssd1 vssd1 vccd1 vccd1 _16524_/S sky130_fd_sc_hd__buf_6
XFILLER_220_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13727_ _13727_/A _13765_/C vssd1 vssd1 vccd1 vccd1 _14021_/C sky130_fd_sc_hd__nor2_4
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17495_ _17495_/A vssd1 vssd1 vccd1 vccd1 _22655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19234_ _19233_/X _23290_/Q _19243_/S vssd1 vssd1 vccd1 vccd1 _19235_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16446_ _16446_/A vssd1 vssd1 vccd1 vccd1 _22383_/D sky130_fd_sc_hd__clkbuf_1
X_13658_ _22613_/Q vssd1 vssd1 vccd1 vccd1 _13669_/A sky130_fd_sc_hd__inv_2
XFILLER_220_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _12110_/S _20234_/A _11935_/X vssd1 vssd1 vccd1 vccd1 _12611_/B sky130_fd_sc_hd__a21boi_4
X_16377_ _16124_/X _22354_/Q _16377_/S vssd1 vssd1 vccd1 vccd1 _16378_/A sky130_fd_sc_hd__mux2_1
X_19165_ _19246_/A vssd1 vssd1 vccd1 vccd1 _19265_/S sky130_fd_sc_hd__buf_8
X_13589_ _13632_/B _13632_/C _13632_/A vssd1 vssd1 vccd1 vccd1 _13633_/A sky130_fd_sc_hd__o21a_2
XFILLER_319_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_334_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18116_ _18116_/A _18166_/B vssd1 vssd1 vccd1 vccd1 _18116_/Y sky130_fd_sc_hd__nand2_2
XFILLER_200_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15328_ _21673_/A vssd1 vssd1 vccd1 vccd1 _15329_/A sky130_fd_sc_hd__buf_8
XFILLER_219_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_346_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19096_ _23238_/Q _18776_/X _19102_/S vssd1 vssd1 vccd1 vccd1 _19097_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_134_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _22600_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_333_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15259_ _22923_/Q _15259_/B vssd1 vssd1 vccd1 vccd1 _15259_/X sky130_fd_sc_hd__and2_1
X_18047_ _22853_/Q _18036_/X _18037_/X _22986_/Q _18038_/X vssd1 vssd1 vccd1 vccd1
+ _18047_/X sky130_fd_sc_hd__a221o_1
XFILLER_322_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_287_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_302_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19998_ _20027_/A _19998_/B vssd1 vssd1 vccd1 vccd1 _19998_/Y sky130_fd_sc_hd__nor2_1
XFILLER_301_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18949_ _16813_/X _23173_/Q _18957_/S vssd1 vssd1 vccd1 vccd1 _18950_/A sky130_fd_sc_hd__mux2_1
XFILLER_301_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21960_ _21975_/A _22044_/A _21959_/Y _22048_/A vssd1 vssd1 vccd1 vccd1 _22041_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_239_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20911_ _20925_/A vssd1 vssd1 vccd1 vccd1 _20911_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_215_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21891_ _21890_/X _21858_/Y _21857_/X vssd1 vssd1 vccd1 vccd1 _21892_/B sky130_fd_sc_hd__a21oi_1
XFILLER_243_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23630_ _23634_/CLK _23630_/D vssd1 vssd1 vccd1 vccd1 _23630_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20842_ _20689_/B _20828_/X _20829_/X _23767_/Q vssd1 vssd1 vccd1 vccd1 _20843_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23561_ _23561_/CLK _23561_/D vssd1 vssd1 vccd1 vccd1 _23561_/Q sky130_fd_sc_hd__dfxtp_1
X_20773_ _20773_/A _20781_/A vssd1 vssd1 vccd1 vccd1 _20773_/Y sky130_fd_sc_hd__nor2_1
XINSDIODE2_370 _23483_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_381 _22517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22512_ _23692_/CLK _22512_/D vssd1 vssd1 vccd1 vccd1 _22512_/Q sky130_fd_sc_hd__dfxtp_4
XINSDIODE2_392 _14090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23492_ _23556_/CLK _23492_/D vssd1 vssd1 vccd1 vccd1 _23492_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_309_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22443_ _23546_/CLK _22443_/D vssd1 vssd1 vccd1 vccd1 _22443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22374_ _23574_/CLK _22374_/D vssd1 vssd1 vccd1 vccd1 _22374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21325_ _17653_/A _21319_/Y _21594_/B vssd1 vssd1 vccd1 vccd1 _21325_/X sky130_fd_sc_hd__mux2_1
XFILLER_324_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_312_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_306_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21256_ _21256_/A vssd1 vssd1 vccd1 vccd1 _23898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20207_ _21444_/A _20340_/B vssd1 vssd1 vccd1 vccd1 _20209_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21187_ _23877_/Q _21168_/X _21184_/X _21186_/X vssd1 vssd1 vccd1 vccd1 _23877_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_278_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20138_ _20191_/A _20138_/B _20214_/B vssd1 vssd1 vccd1 vccd1 _20186_/B sky130_fd_sc_hd__or3_2
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_292_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20069_ _21122_/A _20069_/B vssd1 vssd1 vccd1 vccd1 _20069_/Y sky130_fd_sc_hd__nor2_1
XINSDIODE2_30 _18135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12960_ _12707_/X _12953_/X _12955_/X _12959_/X _11378_/A vssd1 vssd1 vccd1 vccd1
+ _12960_/X sky130_fd_sc_hd__a311o_2
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_41 _20713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_52 _20678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ _23907_/Q _11911_/B vssd1 vssd1 vccd1 vccd1 _11911_/X sky130_fd_sc_hd__or2_1
XFILLER_18_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_63 _21215_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_74 _21077_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12891_ _12891_/A _12891_/B vssd1 vssd1 vccd1 vccd1 _12891_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_85 _14179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_96 _20303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14630_ _15253_/A vssd1 vssd1 vccd1 vccd1 _14630_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _23902_/Q vssd1 vssd1 vccd1 vccd1 _11843_/A sky130_fd_sc_hd__buf_2
X_23828_ _23832_/CLK _23828_/D vssd1 vssd1 vccd1 vccd1 _23828_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _16198_/S vssd1 vssd1 vccd1 vccd1 _14985_/S sky130_fd_sc_hd__buf_6
XFILLER_242_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11773_ _23215_/Q _23183_/Q _23151_/Q _23119_/Q _11708_/S _11613_/A vssd1 vssd1 vccd1
+ vccd1 _11774_/B sky130_fd_sc_hd__mux4_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23759_ _23862_/CLK _23759_/D vssd1 vssd1 vccd1 vccd1 _23759_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_348_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _18865_/A vssd1 vssd1 vccd1 vccd1 _16300_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _11935_/B _21444_/A _12338_/Y vssd1 vssd1 vccd1 vccd1 _13514_/B sky130_fd_sc_hd__a21oi_4
X_17280_ _23488_/Q _17230_/X _17231_/X _17268_/X _17279_/Y vssd1 vssd1 vccd1 vccd1
+ _17280_/X sky130_fd_sc_hd__a32o_1
XFILLER_207_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _15592_/A vssd1 vssd1 vccd1 vccd1 _15210_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_347_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16231_ _22300_/Q _16230_/X _16237_/S vssd1 vssd1 vccd1 vccd1 _16232_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13443_ _14866_/A _20532_/B _20214_/B _20532_/C vssd1 vssd1 vccd1 vccd1 _13455_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_13_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16162_ _16161_/X _22291_/Q _16198_/S vssd1 vssd1 vccd1 vccd1 _16163_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13374_ _13375_/A _13375_/B _13943_/A vssd1 vssd1 vccd1 vccd1 _13382_/C sky130_fd_sc_hd__o21bai_1
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_315_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15113_ _15113_/A _15113_/B vssd1 vssd1 vccd1 vccd1 _15113_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12325_ _12329_/A vssd1 vssd1 vccd1 vccd1 _12325_/X sky130_fd_sc_hd__clkbuf_4
X_16093_ _13549_/B _15079_/B _14837_/X vssd1 vssd1 vccd1 vccd1 _16093_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_182_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19921_ _19922_/B _19915_/X _19916_/X _23591_/Q vssd1 vssd1 vccd1 vccd1 _19923_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15044_ _19181_/A vssd1 vssd1 vccd1 vccd1 _15044_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12256_ _12256_/A _12256_/B vssd1 vssd1 vccd1 vccd1 _12256_/Y sky130_fd_sc_hd__nor2_1
XFILLER_330_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_287_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_11207_ _11207_/A vssd1 vssd1 vccd1 vccd1 _11418_/A sky130_fd_sc_hd__buf_2
X_19852_ _16217_/X _23560_/Q _19854_/S vssd1 vssd1 vccd1 vccd1 _19853_/A sky130_fd_sc_hd__mux2_1
XFILLER_268_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12187_ _11713_/A _12174_/Y _12176_/Y _12186_/X _11214_/A vssd1 vssd1 vccd1 vccd1
+ _12203_/B sky130_fd_sc_hd__o311a_1
X_18803_ _18803_/A vssd1 vssd1 vccd1 vccd1 _23118_/D sky130_fd_sc_hd__clkbuf_1
X_11138_ _11138_/A vssd1 vssd1 vccd1 vccd1 _11834_/A sky130_fd_sc_hd__buf_2
XFILLER_122_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19783_ _19783_/A vssd1 vssd1 vccd1 vccd1 _23529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_311_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16995_ _16976_/X _16979_/X _16983_/X _16994_/X vssd1 vssd1 vccd1 vccd1 _16995_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_352_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18734_ _18734_/A vssd1 vssd1 vccd1 vccd1 _23092_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15946_ _15995_/A _15090_/B _15945_/X vssd1 vssd1 vccd1 vccd1 _15946_/Y sky130_fd_sc_hd__a21oi_1
X_11069_ _23882_/Q _23881_/Q _11069_/C _11069_/D vssd1 vssd1 vccd1 vccd1 _14132_/D
+ sky130_fd_sc_hd__and4bb_2
XFILLER_283_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18665_ _23062_/Q _17601_/X _18669_/S vssd1 vssd1 vccd1 vccd1 _18666_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15877_ _20009_/A _14732_/X _14734_/X _23644_/Q vssd1 vssd1 vccd1 vccd1 _15877_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_237_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_291_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17616_ _17616_/A vssd1 vssd1 vccd1 vccd1 _22699_/D sky130_fd_sc_hd__clkbuf_1
X_14828_ _22498_/Q _14219_/X _14223_/X _14827_/X _14242_/X vssd1 vssd1 vccd1 vccd1
+ _14829_/A sky130_fd_sc_hd__o221a_1
XFILLER_63_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18596_ _18596_/A vssd1 vssd1 vccd1 vccd1 _23031_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17547_ _17646_/S vssd1 vssd1 vccd1 vccd1 _17560_/S sky130_fd_sc_hd__buf_8
X_14759_ _14759_/A _15335_/B vssd1 vssd1 vccd1 vccd1 _14759_/Y sky130_fd_sc_hd__nand2_1
XFILLER_251_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_339_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17478_ _17478_/A vssd1 vssd1 vccd1 vccd1 _22647_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19217_ _19217_/A vssd1 vssd1 vccd1 vccd1 _19217_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16429_ _15749_/X _22376_/Q _16429_/S vssd1 vssd1 vccd1 vccd1 _16430_/A sky130_fd_sc_hd__mux2_1
XFILLER_319_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_301_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19148_ _19148_/A vssd1 vssd1 vccd1 vccd1 _19157_/S sky130_fd_sc_hd__buf_4
XFILLER_30_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19079_ _19079_/A vssd1 vssd1 vccd1 vccd1 _23231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_334_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput500 _14079_/X vssd1 vssd1 vccd1 vccd1 wmask0[3] sky130_fd_sc_hd__buf_2
XFILLER_161_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21110_ _21150_/A vssd1 vssd1 vccd1 vccd1 _21110_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22090_ _22090_/A _22090_/B vssd1 vssd1 vccd1 vccd1 _22090_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21041_ _21149_/A _21043_/B vssd1 vssd1 vccd1 vccd1 _21041_/Y sky130_fd_sc_hd__nand2_1
XFILLER_259_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22992_ _23009_/CLK _22992_/D vssd1 vssd1 vccd1 vccd1 _22992_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_31_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23556_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21943_ _23833_/Q _23767_/Q vssd1 vssd1 vccd1 vccd1 _21945_/A sky130_fd_sc_hd__and2_1
XFILLER_216_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21874_ _21936_/A _21936_/B vssd1 vssd1 vccd1 vccd1 _21933_/A sky130_fd_sc_hd__xnor2_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23613_ _23643_/CLK _23613_/D vssd1 vssd1 vccd1 vccd1 _23613_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_230_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20825_ _20825_/A _20825_/B vssd1 vssd1 vccd1 vccd1 _20826_/A sky130_fd_sc_hd__and2_1
XFILLER_23_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23544_ _23544_/CLK _23544_/D vssd1 vssd1 vccd1 vccd1 _23544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20756_ _16114_/A _20732_/X _20755_/Y vssd1 vssd1 vccd1 vccd1 _20757_/C sky130_fd_sc_hd__a21oi_2
XFILLER_196_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23475_ _23507_/CLK _23475_/D vssd1 vssd1 vccd1 vccd1 _23475_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20687_ _15671_/X _20617_/X _20662_/X vssd1 vssd1 vccd1 vccd1 _20687_/X sky130_fd_sc_hd__a21o_1
X_22426_ _23560_/CLK _22426_/D vssd1 vssd1 vccd1 vccd1 _22426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_356_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_337_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22357_ _23902_/CLK _22357_/D vssd1 vssd1 vccd1 vccd1 _22357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_276_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_313_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12110_ _21719_/A _21716_/A _12110_/S vssd1 vssd1 vccd1 vccd1 _12112_/B sky130_fd_sc_hd__mux2_1
X_21308_ _22711_/Q _21308_/B _21308_/C vssd1 vssd1 vccd1 vccd1 _21560_/A sky130_fd_sc_hd__and3_4
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13090_ _22480_/Q _22640_/Q _13090_/S vssd1 vssd1 vccd1 vccd1 _13090_/X sky130_fd_sc_hd__mux2_1
XFILLER_297_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22288_ _23584_/CLK _22288_/D vssd1 vssd1 vccd1 vccd1 _22288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12041_ _12041_/A vssd1 vssd1 vccd1 vccd1 _12041_/X sky130_fd_sc_hd__buf_4
XFILLER_172_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21239_ _21720_/A _21229_/X _21238_/Y _21236_/X vssd1 vssd1 vccd1 vccd1 _23892_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15800_ _13492_/B _14674_/X _15799_/X vssd1 vssd1 vccd1 vccd1 _15800_/Y sky130_fd_sc_hd__a21oi_2
X_16780_ _22511_/Q _16765_/X _16766_/X input26/X vssd1 vssd1 vccd1 vccd1 _16781_/B
+ sky130_fd_sc_hd__o22a_1
X_13992_ _13992_/A vssd1 vssd1 vccd1 vccd1 _13992_/X sky130_fd_sc_hd__buf_6
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12943_ _22377_/Q _22409_/Q _22698_/Q _23065_/Q _12727_/X _12728_/X vssd1 vssd1 vccd1
+ vccd1 _12944_/B sky130_fd_sc_hd__mux4_1
XFILLER_234_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15731_ _23768_/Q _14910_/A _14912_/A _15729_/X _15730_/X vssd1 vssd1 vccd1 vccd1
+ _15731_/X sky130_fd_sc_hd__a221o_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ _18520_/A vssd1 vssd1 vccd1 vccd1 _18480_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _11587_/A _12873_/X _12759_/A vssd1 vssd1 vccd1 vccd1 _12874_/X sky130_fd_sc_hd__a21o_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _15923_/A _15658_/X _15661_/Y _15480_/X vssd1 vssd1 vccd1 vccd1 _15662_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _17469_/S vssd1 vssd1 vccd1 vccd1 _17410_/S sky130_fd_sc_hd__clkbuf_8
X_14613_ _23814_/Q _14464_/X _14599_/X _14608_/X _14612_/X vssd1 vssd1 vccd1 vccd1
+ _14613_/X sky130_fd_sc_hd__a221o_1
X_11825_ _11926_/A _11822_/X _11824_/X _11680_/A vssd1 vssd1 vccd1 vccd1 _11826_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18381_ _15207_/X _18384_/C _18380_/X vssd1 vssd1 vccd1 vccd1 _18381_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_221_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15593_ _15593_/A vssd1 vssd1 vccd1 vccd1 _15593_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17332_ _17332_/A vssd1 vssd1 vccd1 vccd1 _22588_/D sky130_fd_sc_hd__clkbuf_1
X_14544_ _14541_/X _15519_/A _14543_/X vssd1 vssd1 vccd1 vccd1 _19090_/A sky130_fd_sc_hd__o21ai_2
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _22788_/Q _22756_/Q _22657_/Q _22724_/Q _11741_/X _12025_/A vssd1 vssd1 vccd1
+ vccd1 _11757_/B sky130_fd_sc_hd__mux4_1
XFILLER_159_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_347_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17263_ _17245_/X _17261_/X _17262_/X _17215_/X vssd1 vssd1 vccd1 vccd1 _17263_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14475_ _14468_/B _21097_/A _14595_/B vssd1 vssd1 vccd1 vccd1 _14912_/A sky130_fd_sc_hd__a21oi_2
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11687_ _11935_/B vssd1 vssd1 vccd1 vccd1 _12110_/S sky130_fd_sc_hd__buf_8
XFILLER_128_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_335_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19002_ _19002_/A vssd1 vssd1 vccd1 vccd1 _23197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16214_ _18779_/A vssd1 vssd1 vccd1 vccd1 _16214_/X sky130_fd_sc_hd__clkbuf_2
X_13426_ _14176_/A _14250_/A vssd1 vssd1 vccd1 vccd1 _14792_/A sky130_fd_sc_hd__nand2_2
X_17194_ _21916_/A _17193_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17194_/X sky130_fd_sc_hd__mux2_1
XFILLER_347_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16145_ _22944_/Q _14988_/B _16144_/X _14898_/A vssd1 vssd1 vccd1 vccd1 _16145_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13357_ _14687_/A vssd1 vssd1 vccd1 vccd1 _13367_/A sky130_fd_sc_hd__inv_2
XFILLER_289_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12308_ _23466_/Q _23562_/Q _22526_/Q _22330_/Q _12242_/S _11611_/A vssd1 vssd1 vccd1
+ vccd1 _12308_/X sky130_fd_sc_hd__mux4_1
XFILLER_343_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_304_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16076_ _22165_/A _16077_/B vssd1 vssd1 vccd1 vccd1 _16151_/C sky130_fd_sc_hd__and2_1
X_13288_ _22385_/Q _22417_/Q _22706_/Q _23073_/Q _13275_/X _13276_/X vssd1 vssd1 vccd1
+ vccd1 _13288_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19904_ _19904_/A vssd1 vssd1 vccd1 vccd1 _23583_/D sky130_fd_sc_hd__clkbuf_1
X_15027_ _22516_/Q _14219_/A _14238_/A _15026_/X _15056_/A vssd1 vssd1 vccd1 vccd1
+ _15432_/A sky130_fd_sc_hd__o221ai_4
X_12239_ _12256_/A _12239_/B vssd1 vssd1 vccd1 vccd1 _12239_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_297_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19835_ _23553_/Q _19255_/A _19837_/S vssd1 vssd1 vccd1 vccd1 _19836_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19766_ _19766_/A vssd1 vssd1 vccd1 vccd1 _23522_/D sky130_fd_sc_hd__clkbuf_1
X_16978_ _17244_/C vssd1 vssd1 vccd1 vccd1 _16978_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput4 coreIndex[3] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_4
XFILLER_237_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18717_ _16841_/X _23085_/Q _18719_/S vssd1 vssd1 vccd1 vccd1 _18718_/A sky130_fd_sc_hd__mux2_1
X_15929_ _15929_/A vssd1 vssd1 vccd1 vccd1 _15929_/X sky130_fd_sc_hd__buf_6
XFILLER_37_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19697_ _19264_/X _23492_/Q _19697_/S vssd1 vssd1 vccd1 vccd1 _19698_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18648_ _18648_/A vssd1 vssd1 vccd1 vccd1 _23054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18579_ _18579_/A vssd1 vssd1 vccd1 vccd1 _23023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20610_ _21013_/A _20891_/A vssd1 vssd1 vccd1 vccd1 _20613_/B sky130_fd_sc_hd__nor2_4
XFILLER_189_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21590_ _21601_/A _21594_/A vssd1 vssd1 vccd1 vccd1 _21593_/A sky130_fd_sc_hd__xnor2_1
XFILLER_193_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20541_ _20729_/A vssd1 vssd1 vccd1 vccd1 _20628_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_327_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_326_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23260_ _23420_/CLK _23260_/D vssd1 vssd1 vccd1 vccd1 _23260_/Q sky130_fd_sc_hd__dfxtp_1
X_20472_ _20602_/A vssd1 vssd1 vccd1 vccd1 _20472_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_335_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22211_ _22211_/A _22210_/X vssd1 vssd1 vccd1 vccd1 _22213_/A sky130_fd_sc_hd__or2b_1
X_23191_ _23511_/CLK _23191_/D vssd1 vssd1 vccd1 vccd1 _23191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_350_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22142_ _22168_/A _22142_/B _22142_/C vssd1 vssd1 vccd1 vccd1 _22142_/X sky130_fd_sc_hd__or3_1
XFILLER_350_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput330 _13947_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[9] sky130_fd_sc_hd__buf_2
XFILLER_105_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput341 _13802_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[18] sky130_fd_sc_hd__buf_2
XTAP_6707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput352 _13861_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[28] sky130_fd_sc_hd__buf_2
XFILLER_161_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22073_ _20362_/A _22045_/X _15941_/X _22046_/X vssd1 vssd1 vccd1 vccd1 _22073_/X
+ sky130_fd_sc_hd__a22o_1
Xoutput363 _13748_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[9] sky130_fd_sc_hd__buf_2
XTAP_6729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput374 _14007_/X vssd1 vssd1 vccd1 vccd1 din0[0] sky130_fd_sc_hd__buf_2
Xoutput385 _14010_/X vssd1 vssd1 vccd1 vccd1 din0[1] sky130_fd_sc_hd__buf_2
XFILLER_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput396 _14014_/X vssd1 vssd1 vccd1 vccd1 din0[2] sky130_fd_sc_hd__buf_2
XFILLER_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21024_ _20639_/A _21008_/X _21022_/X _21023_/X vssd1 vssd1 vccd1 vccd1 _23824_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_303_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_288_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22975_ _22977_/CLK _22975_/D vssd1 vssd1 vccd1 vccd1 _22975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21926_ _22012_/A _22012_/B vssd1 vssd1 vccd1 vccd1 _21987_/A sky130_fd_sc_hd__nor2_2
XFILLER_76_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21857_ _23928_/Q _21861_/A vssd1 vssd1 vccd1 vccd1 _21857_/X sky130_fd_sc_hd__and2_1
XFILLER_70_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_358_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11610_ _12292_/A vssd1 vssd1 vccd1 vccd1 _11611_/A sky130_fd_sc_hd__buf_6
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20808_ _20808_/A vssd1 vssd1 vccd1 vccd1 _20881_/A sky130_fd_sc_hd__buf_6
XFILLER_168_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12590_ _12590_/A _12590_/B vssd1 vssd1 vccd1 vccd1 _12590_/X sky130_fd_sc_hd__or2_1
XFILLER_298_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21788_ _23828_/Q _21787_/Y _22019_/A vssd1 vssd1 vccd1 vccd1 _21788_/X sky130_fd_sc_hd__mux2_1
XFILLER_243_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11541_ _13073_/A _11541_/B vssd1 vssd1 vccd1 vccd1 _11541_/X sky130_fd_sc_hd__or2_1
X_23527_ _23527_/CLK _23527_/D vssd1 vssd1 vccd1 vccd1 _23527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20739_ _21173_/A _20744_/B vssd1 vssd1 vccd1 vccd1 _20742_/B sky130_fd_sc_hd__nor2_2
XFILLER_204_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_329_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14260_ _14351_/S _13362_/B _14259_/X vssd1 vssd1 vccd1 vccd1 _14260_/X sky130_fd_sc_hd__o21a_2
XFILLER_310_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23458_ _23489_/CLK _23458_/D vssd1 vssd1 vccd1 vccd1 _23458_/Q sky130_fd_sc_hd__dfxtp_1
X_11472_ _23427_/Q _23043_/Q _23395_/Q _23363_/Q _11461_/X _11462_/X vssd1 vssd1 vccd1
+ vccd1 _11472_/X sky130_fd_sc_hd__mux4_1
X_13211_ _13194_/X _13200_/X _13210_/Y vssd1 vssd1 vccd1 vccd1 _13836_/A sky130_fd_sc_hd__o21a_4
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22409_ _23449_/CLK _22409_/D vssd1 vssd1 vccd1 vccd1 _22409_/Q sky130_fd_sc_hd__dfxtp_1
X_14191_ _16005_/A _14564_/A vssd1 vssd1 vccd1 vccd1 _14192_/B sky130_fd_sc_hd__nor2_1
XFILLER_354_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23389_ _23549_/CLK _23389_/D vssd1 vssd1 vccd1 vccd1 _23389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13142_ _22802_/Q _22770_/Q _22671_/Q _22738_/Q _11431_/A _13037_/A vssd1 vssd1 vccd1
+ vccd1 _13143_/B sky130_fd_sc_hd__mux4_2
XFILLER_325_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_317_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_340_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_317_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_352_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_313_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17950_ _17981_/A vssd1 vssd1 vccd1 vccd1 _17950_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_341_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13073_ _13073_/A _13073_/B vssd1 vssd1 vccd1 vccd1 _13073_/Y sky130_fd_sc_hd__nor2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_340_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16901_ _16901_/A vssd1 vssd1 vccd1 vccd1 _22547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_266_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12024_ _12024_/A vssd1 vssd1 vccd1 vccd1 _12024_/X sky130_fd_sc_hd__buf_6
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17881_ _17881_/A vssd1 vssd1 vccd1 vccd1 _22811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_265_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19620_ _19620_/A vssd1 vssd1 vccd1 vccd1 _23457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_333_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16832_ _16915_/S vssd1 vssd1 vccd1 vccd1 _16845_/S sky130_fd_sc_hd__buf_6
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_294_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19551_ _19261_/X _23427_/Q _19553_/S vssd1 vssd1 vccd1 vccd1 _19552_/A sky130_fd_sc_hd__mux2_1
XFILLER_253_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16763_ _16777_/A _16763_/B vssd1 vssd1 vccd1 vccd1 _16764_/A sky130_fd_sc_hd__or2_1
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13975_ _13975_/A _13979_/B vssd1 vssd1 vccd1 vccd1 _13976_/A sky130_fd_sc_hd__and2_1
XFILLER_265_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18502_ _22996_/Q _18505_/B vssd1 vssd1 vccd1 vccd1 _18502_/Y sky130_fd_sc_hd__nand2_1
XFILLER_207_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15714_ _23930_/Q vssd1 vssd1 vccd1 vccd1 _21916_/A sky130_fd_sc_hd__buf_12
XFILLER_62_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12926_ _12926_/A _12926_/B vssd1 vssd1 vccd1 vccd1 _12926_/Y sky130_fd_sc_hd__nor2_1
X_19482_ _19482_/A vssd1 vssd1 vccd1 vccd1 _23396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16694_ _22487_/Q _16689_/X _16693_/X input10/X vssd1 vssd1 vccd1 vccd1 _16695_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18433_ _18435_/A _18435_/C _18432_/Y vssd1 vssd1 vccd1 vccd1 _22972_/D sky130_fd_sc_hd__o21a_1
X_15645_ _23606_/Q _14732_/X _14734_/X _23638_/Q vssd1 vssd1 vccd1 vccd1 _15645_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_221_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _22380_/Q _22412_/Q _22701_/Q _23068_/Q _12709_/X _12710_/X vssd1 vssd1 vccd1
+ vccd1 _12857_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18364_ _19932_/A vssd1 vssd1 vccd1 vccd1 _18401_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_203_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ _12144_/A _11808_/B vssd1 vssd1 vccd1 vccd1 _11808_/X sky130_fd_sc_hd__or2_1
XFILLER_348_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12788_ _23223_/Q _23191_/Q _23159_/Q _23127_/Q _12776_/X _12777_/X vssd1 vssd1 vccd1
+ vccd1 _12789_/B sky130_fd_sc_hd__mux4_2
XFILLER_187_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15576_ _15576_/A _15901_/B vssd1 vssd1 vccd1 vccd1 _15576_/Y sky130_fd_sc_hd__nor2_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _23942_/Q vssd1 vssd1 vccd1 vccd1 _17315_/X sky130_fd_sc_hd__buf_8
X_11739_ _12141_/A _11738_/X _11681_/A vssd1 vssd1 vccd1 vccd1 _11739_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_202_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14527_ _14539_/S vssd1 vssd1 vccd1 vccd1 _14557_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18295_ _18296_/A _18296_/C _22925_/Q vssd1 vssd1 vccd1 vccd1 _18297_/B sky130_fd_sc_hd__a21oi_1
XFILLER_187_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_358_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17246_ _17246_/A vssd1 vssd1 vccd1 vccd1 _22064_/A sky130_fd_sc_hd__clkbuf_16
X_14458_ _14458_/A _14458_/B _14416_/B _14416_/A vssd1 vssd1 vccd1 vccd1 _14465_/C
+ sky130_fd_sc_hd__or4bb_1
XFILLER_317_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13409_ _13409_/A _13409_/B _13406_/Y _13408_/Y vssd1 vssd1 vccd1 vccd1 _13410_/D
+ sky130_fd_sc_hd__or4bb_2
X_17177_ _17167_/X _17168_/X _17175_/X _17176_/X vssd1 vssd1 vccd1 vccd1 _17177_/X
+ sky130_fd_sc_hd__o211a_4
X_14389_ _14261_/X _14389_/B _14389_/C vssd1 vssd1 vccd1 vccd1 _14389_/X sky130_fd_sc_hd__and3b_1
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16128_ _14793_/A _14676_/B _16128_/S vssd1 vssd1 vccd1 vccd1 _16128_/X sky130_fd_sc_hd__mux2_1
XFILLER_227_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_289_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_304_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16059_ _22942_/Q vssd1 vssd1 vccd1 vccd1 _16059_/X sky130_fd_sc_hd__buf_2
XFILLER_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19818_ _23545_/Q _19229_/A _19826_/S vssd1 vssd1 vccd1 vccd1 _19819_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19749_ _19749_/A vssd1 vssd1 vccd1 vccd1 _23514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_272_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22760_ _23450_/CLK _22760_/D vssd1 vssd1 vccd1 vccd1 _22760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21711_ _21711_/A _21711_/B vssd1 vssd1 vccd1 vccd1 _21711_/X sky130_fd_sc_hd__xor2_1
XFILLER_213_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22691_ _23058_/CLK _22691_/D vssd1 vssd1 vccd1 vccd1 _22691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_358_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21642_ _21829_/B _21640_/Y _21641_/Y _21327_/A vssd1 vssd1 vccd1 vccd1 _21643_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21573_ _21513_/A _21509_/Y _21513_/B _21511_/B vssd1 vssd1 vccd1 vccd1 _21574_/B
+ sky130_fd_sc_hd__o31ai_4
XFILLER_138_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23312_ _23409_/CLK _23312_/D vssd1 vssd1 vccd1 vccd1 _23312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_354_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_326_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20524_ _23703_/Q _20524_/B _20524_/C vssd1 vssd1 vccd1 vccd1 _20525_/D sky130_fd_sc_hd__and3_1
XFILLER_268_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23243_ _23467_/CLK _23243_/D vssd1 vssd1 vccd1 vccd1 _23243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20455_ _23701_/Q _20468_/B vssd1 vssd1 vccd1 vccd1 _20455_/X sky130_fd_sc_hd__or2_1
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23174_ _23496_/CLK _23174_/D vssd1 vssd1 vccd1 vccd1 _23174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20386_ _20333_/X _20749_/A _20385_/X _20360_/X vssd1 vssd1 vccd1 vccd1 _23681_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_7227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22125_ _20374_/A _22045_/X _16041_/Y _21842_/X vssd1 vssd1 vccd1 vccd1 _22125_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_7249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22056_ _23837_/Q _23771_/Q vssd1 vssd1 vccd1 vccd1 _22057_/B sky130_fd_sc_hd__nor2_1
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21007_ _20595_/A _20988_/X _21006_/X _20997_/X vssd1 vssd1 vccd1 vccd1 _23818_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_303_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13760_ _13974_/B _14032_/C vssd1 vssd1 vccd1 vccd1 _13760_/Y sky130_fd_sc_hd__nor2_1
X_22958_ _22961_/CLK _22958_/D vssd1 vssd1 vccd1 vccd1 _22958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12711_ _22280_/Q _23096_/Q _23512_/Q _22441_/Q _12709_/X _12710_/X vssd1 vssd1 vccd1
+ vccd1 _12712_/B sky130_fd_sc_hd__mux4_1
XFILLER_271_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21909_ _23832_/Q _23766_/Q vssd1 vssd1 vccd1 vccd1 _21911_/A sky130_fd_sc_hd__nor2_1
XFILLER_43_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13691_ _13691_/A vssd1 vssd1 vccd1 vccd1 _13692_/A sky130_fd_sc_hd__buf_2
XFILLER_188_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22889_ _23327_/CLK _22889_/D vssd1 vssd1 vccd1 vccd1 _22889_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_188_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12642_ _22793_/Q _22761_/Q _22662_/Q _22729_/Q _11972_/X _11973_/X vssd1 vssd1 vccd1
+ vccd1 _12642_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15430_ _21737_/A _15430_/B vssd1 vssd1 vccd1 vccd1 _15431_/B sky130_fd_sc_hd__nor2_1
XFILLER_231_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15361_ _22925_/Q _14868_/B _15351_/X _15360_/Y _14727_/X vssd1 vssd1 vccd1 vccd1
+ _15361_/X sky130_fd_sc_hd__a221o_1
XPHY_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12573_ _23890_/Q _13472_/A _12371_/B vssd1 vssd1 vccd1 vccd1 _12573_/X sky130_fd_sc_hd__a21bo_1
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_346_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17100_ _17070_/X _17093_/X _17099_/X _17057_/X vssd1 vssd1 vccd1 vccd1 _17100_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_168_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11524_ _11532_/A vssd1 vssd1 vccd1 vccd1 _13114_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_196_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14312_ _14303_/X _14311_/X _15129_/S vssd1 vssd1 vccd1 vccd1 _14312_/X sky130_fd_sc_hd__mux2_2
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18080_ _22865_/Q _18066_/X _18079_/X _18075_/X vssd1 vssd1 vccd1 vccd1 _22865_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15292_ _15012_/Y _15291_/X _15292_/S vssd1 vssd1 vccd1 vccd1 _15801_/B sky130_fd_sc_hd__mux2_1
XFILLER_317_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_317_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17031_ _17248_/A vssd1 vssd1 vccd1 vccd1 _17144_/A sky130_fd_sc_hd__buf_2
X_14243_ _22495_/Q _13692_/A _14238_/X _14240_/X _14242_/X vssd1 vssd1 vccd1 vccd1
+ _14243_/Y sky130_fd_sc_hd__o221ai_4
X_11455_ _11455_/A vssd1 vssd1 vccd1 vccd1 _11745_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_184_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_314_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_326_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14174_ _14198_/C vssd1 vssd1 vccd1 vccd1 _15672_/A sky130_fd_sc_hd__buf_2
X_11386_ _11828_/B vssd1 vssd1 vccd1 vccd1 _12157_/S sky130_fd_sc_hd__buf_2
XFILLER_139_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13125_ _23231_/Q _23199_/Q _23167_/Q _23135_/Q _13114_/X _13115_/X vssd1 vssd1 vccd1
+ vccd1 _13126_/B sky130_fd_sc_hd__mux4_1
XFILLER_298_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18982_ _16863_/X _23188_/Q _18990_/S vssd1 vssd1 vccd1 vccd1 _18983_/A sky130_fd_sc_hd__mux2_1
XFILLER_314_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17933_ _17933_/A vssd1 vssd1 vccd1 vccd1 _17933_/X sky130_fd_sc_hd__clkbuf_2
X_13056_ _13273_/A _13056_/B vssd1 vssd1 vccd1 vccd1 _13056_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_340_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12007_ _12007_/A vssd1 vssd1 vccd1 vccd1 _12949_/A sky130_fd_sc_hd__buf_2
XFILLER_289_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17864_ _22803_/Q _17630_/X _17870_/S vssd1 vssd1 vccd1 vccd1 _17865_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_159_wb_clk_i _23945_/CLK vssd1 vssd1 vccd1 vccd1 _23832_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_293_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19603_ _19603_/A vssd1 vssd1 vccd1 vccd1 _23449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16815_ _16896_/A vssd1 vssd1 vccd1 vccd1 _16915_/S sky130_fd_sc_hd__buf_6
XFILLER_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_293_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17795_ _17795_/A vssd1 vssd1 vccd1 vccd1 _22772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_253_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19534_ _19236_/X _23419_/Q _19538_/S vssd1 vssd1 vccd1 vccd1 _19535_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16746_ _16746_/A vssd1 vssd1 vccd1 vccd1 _22501_/D sky130_fd_sc_hd__clkbuf_1
X_13958_ _14198_/B vssd1 vssd1 vccd1 vccd1 _21289_/A sky130_fd_sc_hd__buf_4
XFILLER_253_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19465_ _19465_/A vssd1 vssd1 vccd1 vccd1 _23388_/D sky130_fd_sc_hd__clkbuf_1
X_12909_ _12909_/A _12909_/B vssd1 vssd1 vccd1 vccd1 _12909_/X sky130_fd_sc_hd__or2_1
XFILLER_59_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16677_ _22485_/Q _16306_/X _16677_/S vssd1 vssd1 vccd1 vccd1 _16678_/A sky130_fd_sc_hd__mux2_1
X_13889_ _13889_/A vssd1 vssd1 vccd1 vccd1 _13889_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18416_ _18418_/A _18418_/C _18415_/Y vssd1 vssd1 vccd1 vccd1 _22966_/D sky130_fd_sc_hd__o21a_1
XFILLER_179_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15628_ _22995_/Q _15780_/A _15781_/A input223/X vssd1 vssd1 vccd1 vccd1 _21890_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19396_ _19396_/A vssd1 vssd1 vccd1 vccd1 _19405_/S sky130_fd_sc_hd__buf_4
XFILLER_50_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18347_ _16059_/X _18349_/C _18346_/Y vssd1 vssd1 vccd1 vccd1 _22942_/D sky130_fd_sc_hd__o21a_1
XFILLER_309_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15559_ _22929_/Q _14728_/B _15548_/X _15557_/Y _15558_/X vssd1 vssd1 vccd1 vccd1
+ _15559_/X sky130_fd_sc_hd__a221o_1
XFILLER_349_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_337_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18278_ _19962_/A vssd1 vssd1 vccd1 vccd1 _18317_/A sky130_fd_sc_hd__buf_2
XFILLER_175_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_352_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_336_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput40 core_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_1
X_17229_ _17229_/A vssd1 vssd1 vccd1 vccd1 _22029_/A sky130_fd_sc_hd__buf_8
XFILLER_174_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput51 dout0[17] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_2
XFILLER_317_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput62 dout0[27] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__buf_2
XFILLER_305_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput73 dout0[37] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_1
XFILLER_337_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput84 dout0[47] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__clkbuf_1
X_20240_ _20213_/X _20615_/A _20239_/X _20203_/X vssd1 vssd1 vccd1 vccd1 _23661_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_351_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput95 dout0[57] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__clkbuf_1
XFILLER_337_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20171_ _17159_/A _12493_/X _20394_/B vssd1 vssd1 vccd1 vccd1 _20171_/X sky130_fd_sc_hd__mux2_1
XFILLER_331_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23930_ _23938_/CLK _23930_/D vssd1 vssd1 vccd1 vccd1 _23930_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_229_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23861_ _23861_/CLK _23861_/D vssd1 vssd1 vccd1 vccd1 _23861_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22812_ _22968_/CLK _22812_/D vssd1 vssd1 vccd1 vccd1 _22812_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23792_ _23861_/CLK _23792_/D vssd1 vssd1 vccd1 vccd1 _23792_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_232_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22743_ _23893_/CLK _22743_/D vssd1 vssd1 vccd1 vccd1 _22743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_344_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22674_ _23581_/CLK _22674_/D vssd1 vssd1 vccd1 vccd1 _22674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21625_ _21625_/A _21625_/B vssd1 vssd1 vccd1 vccd1 _21625_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21556_ _21865_/A vssd1 vssd1 vccd1 vccd1 _21556_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20507_ _23710_/Q _20508_/B _20507_/C vssd1 vssd1 vccd1 vccd1 _20509_/C sky130_fd_sc_hd__and3_1
XFILLER_194_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21487_ _21542_/A _21487_/B vssd1 vssd1 vccd1 vccd1 _21487_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_355_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23226_ _23419_/CLK _23226_/D vssd1 vssd1 vccd1 vccd1 _23226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_314_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11240_ _11240_/A vssd1 vssd1 vccd1 vccd1 _11241_/A sky130_fd_sc_hd__clkinv_4
X_20438_ _23694_/Q _20448_/B vssd1 vssd1 vccd1 vccd1 _20438_/X sky130_fd_sc_hd__or2_1
XFILLER_153_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_7013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23157_ _23349_/CLK _23157_/D vssd1 vssd1 vccd1 vccd1 _23157_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_7035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11171_ _23236_/Q _23204_/Q _23172_/Q _23140_/Q _11157_/X _11170_/X vssd1 vssd1 vccd1
+ vccd1 _11172_/B sky130_fd_sc_hd__mux4_1
XFILLER_107_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20369_ _17269_/A _20215_/X _20368_/X vssd1 vssd1 vccd1 vccd1 _20369_/Y sky130_fd_sc_hd__o21ai_1
XTAP_7046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22108_ _23839_/Q _23773_/Q vssd1 vssd1 vccd1 vccd1 _22108_/Y sky130_fd_sc_hd__nand2_1
XTAP_7079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23088_ _23504_/CLK _23088_/D vssd1 vssd1 vccd1 vccd1 _23088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14930_ _22918_/Q vssd1 vssd1 vccd1 vccd1 _18275_/A sky130_fd_sc_hd__clkbuf_2
X_22039_ _22039_/A _22040_/B vssd1 vssd1 vccd1 vccd1 _22039_/Y sky130_fd_sc_hd__nand2_1
XTAP_6389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14861_ _15292_/S _14859_/Y _14860_/X vssd1 vssd1 vccd1 vccd1 _14861_/X sky130_fd_sc_hd__a21o_1
XFILLER_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16600_ _16600_/A vssd1 vssd1 vccd1 vccd1 _22450_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ _13855_/A _13812_/B vssd1 vssd1 vccd1 vccd1 _13813_/A sky130_fd_sc_hd__and2_1
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17580_ _22688_/Q _17578_/X _17592_/S vssd1 vssd1 vccd1 vccd1 _17581_/A sky130_fd_sc_hd__mux2_1
XFILLER_290_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14792_ _14792_/A vssd1 vssd1 vccd1 vccd1 _14793_/A sky130_fd_sc_hd__buf_4
XFILLER_235_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16531_ _17382_/A vssd1 vssd1 vccd1 vccd1 _18277_/A sky130_fd_sc_hd__clkbuf_4
X_13743_ _13934_/A vssd1 vssd1 vccd1 vccd1 _13893_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19250_ _19249_/X _23295_/Q _19259_/S vssd1 vssd1 vccd1 vccd1 _19251_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16462_ _16462_/A vssd1 vssd1 vccd1 vccd1 _22389_/D sky130_fd_sc_hd__clkbuf_1
X_13674_ _17039_/A vssd1 vssd1 vccd1 vccd1 _17219_/S sky130_fd_sc_hd__buf_4
XFILLER_177_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18201_ _22872_/Q _18203_/B _18203_/C vssd1 vssd1 vccd1 vccd1 _18242_/A sky130_fd_sc_hd__or3_4
XFILLER_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15413_ _15672_/A vssd1 vssd1 vccd1 vccd1 _15574_/A sky130_fd_sc_hd__clkbuf_2
X_12625_ _23221_/Q _23189_/Q _23157_/Q _23125_/Q _12008_/X _12734_/A vssd1 vssd1 vccd1
+ vccd1 _12626_/B sky130_fd_sc_hd__mux4_2
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19181_ _19181_/A vssd1 vssd1 vccd1 vccd1 _19181_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16393_ _16393_/A vssd1 vssd1 vccd1 vccd1 _22359_/D sky130_fd_sc_hd__clkbuf_1
XPHY_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18132_ _14119_/A _22881_/Q _18187_/A vssd1 vssd1 vccd1 vccd1 _18132_/X sky130_fd_sc_hd__mux2_1
XPHY_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12556_ _12556_/A _22297_/Q vssd1 vssd1 vccd1 vccd1 _12556_/X sky130_fd_sc_hd__or2_1
XFILLER_106_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15344_ _13528_/A _15082_/X _15338_/X _15343_/X vssd1 vssd1 vccd1 vccd1 _15345_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_346_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_334_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11507_ _23490_/Q _23586_/Q _22550_/Q _22354_/Q _13255_/S _11418_/A vssd1 vssd1 vccd1
+ vccd1 _11507_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18063_ hold7/A _18051_/X _18062_/X _18060_/X vssd1 vssd1 vccd1 vccd1 _22859_/D sky130_fd_sc_hd__o211a_1
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12487_ _12489_/A _12486_/X _11818_/A vssd1 vssd1 vccd1 vccd1 _12487_/X sky130_fd_sc_hd__o21a_1
X_15275_ _21570_/A _15274_/C _13945_/B vssd1 vssd1 vccd1 vccd1 _15276_/B sky130_fd_sc_hd__a21oi_1
XFILLER_184_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17014_ _22555_/Q _16922_/X _16973_/X _17013_/X vssd1 vssd1 vccd1 vccd1 _22555_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_208_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14226_ _15114_/S vssd1 vssd1 vccd1 vccd1 _15057_/S sky130_fd_sc_hd__clkbuf_4
X_11438_ _22323_/Q _23459_/Q _13254_/S vssd1 vssd1 vccd1 vccd1 _11438_/X sky130_fd_sc_hd__mux2_1
XFILLER_355_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_342_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14157_ _16937_/A _16949_/A vssd1 vssd1 vccd1 vccd1 _21294_/A sky130_fd_sc_hd__nand2_2
XFILLER_98_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11369_ _13291_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11369_/X sky130_fd_sc_hd__or2_1
XFILLER_152_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_313_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13108_ _13101_/Y _13103_/Y _13105_/Y _13107_/Y _11247_/A vssd1 vssd1 vccd1 vccd1
+ _13108_/X sky130_fd_sc_hd__o221a_1
XFILLER_302_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_298_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14088_ _22591_/Q _14081_/X _14087_/Y _14083_/X vssd1 vssd1 vccd1 vccd1 _14088_/X
+ sky130_fd_sc_hd__a22o_4
X_18965_ _18965_/A vssd1 vssd1 vccd1 vccd1 _23180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17916_ _22817_/Q _17908_/X _17903_/X input258/X _17915_/X vssd1 vssd1 vccd1 vccd1
+ _17916_/X sky130_fd_sc_hd__a221o_1
X_13039_ _13041_/A _13039_/B vssd1 vssd1 vccd1 vccd1 _13039_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18896_ _23150_/Q _18801_/X _18896_/S vssd1 vssd1 vccd1 vccd1 _18897_/A sky130_fd_sc_hd__mux2_1
XTAP_6890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_310_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17847_ _17847_/A vssd1 vssd1 vccd1 vccd1 _22795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17778_ _17789_/A vssd1 vssd1 vccd1 vccd1 _17787_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_35_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19517_ _19517_/A vssd1 vssd1 vccd1 vccd1 _23411_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16729_ _16729_/A vssd1 vssd1 vccd1 vccd1 _16729_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_240_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_530 _14127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_541 _23919_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19448_ _19448_/A vssd1 vssd1 vccd1 vccd1 _23380_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_552 _13679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_563 _23911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19379_ _23350_/Q _18827_/X _19383_/S vssd1 vssd1 vccd1 vccd1 _19380_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_56_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23574_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_176_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21410_ _21410_/A vssd1 vssd1 vccd1 vccd1 _21410_/X sky130_fd_sc_hd__buf_2
XFILLER_336_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22390_ _23494_/CLK _22390_/D vssd1 vssd1 vccd1 vccd1 _22390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21341_ _14713_/A _21441_/A _21339_/X _20502_/A _21340_/X vssd1 vssd1 vccd1 vccd1
+ _21342_/B sky130_fd_sc_hd__a221o_1
XFILLER_336_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21272_ _21272_/A _21274_/B vssd1 vssd1 vccd1 vccd1 _21272_/Y sky130_fd_sc_hd__nand2_1
XFILLER_151_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_305_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23011_ _23599_/CLK _23011_/D vssd1 vssd1 vccd1 vccd1 _23011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_265_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20223_ _23659_/Q _20223_/B vssd1 vssd1 vccd1 vccd1 _20223_/X sky130_fd_sc_hd__or2_1
XFILLER_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_333_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_305_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_320_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_289_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20154_ _20168_/A vssd1 vssd1 vccd1 vccd1 _20154_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20085_ _23636_/Q _20090_/C _20085_/C _20085_/D vssd1 vssd1 vccd1 vccd1 _20095_/D
+ sky130_fd_sc_hd__and4_2
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23913_ _23916_/CLK _23913_/D vssd1 vssd1 vccd1 vccd1 _23913_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23844_ _23876_/CLK _23844_/D vssd1 vssd1 vccd1 vccd1 _23844_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23775_ _23804_/CLK _23775_/D vssd1 vssd1 vccd1 vccd1 _23775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20987_ _21047_/A vssd1 vssd1 vccd1 vccd1 _21008_/A sky130_fd_sc_hd__buf_4
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22726_ _23570_/CLK _22726_/D vssd1 vssd1 vccd1 vccd1 _22726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22657_ _23058_/CLK _22657_/D vssd1 vssd1 vccd1 vccd1 _22657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12410_ _12410_/A _12410_/B vssd1 vssd1 vccd1 vccd1 _12410_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21608_ _23790_/Q _22130_/B _21607_/X _21346_/A vssd1 vssd1 vccd1 vccd1 _21608_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_139_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13390_ _12664_/A _12636_/X _13350_/A vssd1 vssd1 vccd1 vccd1 _13391_/B sky130_fd_sc_hd__a21oi_2
X_22588_ _22968_/CLK _22588_/D vssd1 vssd1 vccd1 vccd1 _22588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12341_ _13334_/C vssd1 vssd1 vccd1 vccd1 _13913_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_315_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21539_ _13931_/B _21329_/X _20101_/X vssd1 vssd1 vccd1 vccd1 _21539_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_355_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_309_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_299_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15060_ _22509_/Q _14219_/A _13887_/A _15059_/X vssd1 vssd1 vccd1 vccd1 _15485_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_315_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12272_ _12264_/Y _12266_/Y _12268_/Y _12271_/Y _11273_/A vssd1 vssd1 vccd1 vccd1
+ _12282_/B sky130_fd_sc_hd__o221a_1
XFILLER_331_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14011_ _14072_/C vssd1 vssd1 vccd1 vccd1 _14049_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11223_ _13253_/A vssd1 vssd1 vccd1 vccd1 _15826_/A sky130_fd_sc_hd__buf_6
X_23209_ _23561_/CLK _23209_/D vssd1 vssd1 vccd1 vccd1 _23209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_296_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11154_ _13089_/A vssd1 vssd1 vccd1 vccd1 _13191_/S sky130_fd_sc_hd__clkbuf_4
XTAP_6120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18750_ _16889_/X _23100_/Q _18752_/S vssd1 vssd1 vccd1 vccd1 _18751_/A sky130_fd_sc_hd__mux2_1
XTAP_6175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15962_ _15950_/X _14728_/B _15952_/X _15961_/Y _15558_/X vssd1 vssd1 vccd1 vccd1
+ _15962_/X sky130_fd_sc_hd__a221o_1
XFILLER_191_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11085_ _14195_/A vssd1 vssd1 vccd1 vccd1 _13432_/A sky130_fd_sc_hd__buf_6
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput230 localMemory_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 input230/X sky130_fd_sc_hd__buf_8
XFILLER_310_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17701_ _17701_/A vssd1 vssd1 vccd1 vccd1 _22730_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput241 localMemory_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input241/X sky130_fd_sc_hd__buf_4
XTAP_5463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput252 localMemory_wb_we_i vssd1 vssd1 vccd1 vccd1 _17394_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14913_ _14913_/A vssd1 vssd1 vccd1 vccd1 _14913_/X sky130_fd_sc_hd__buf_2
Xinput263 manufacturerID[9] vssd1 vssd1 vccd1 vccd1 input263/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18681_ _18681_/A vssd1 vssd1 vccd1 vccd1 _23069_/D sky130_fd_sc_hd__clkbuf_1
Xinput274 partID[4] vssd1 vssd1 vccd1 vccd1 input274/X sky130_fd_sc_hd__clkbuf_1
XFILLER_286_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15893_ _15162_/A _13592_/Y _15478_/A vssd1 vssd1 vccd1 vccd1 _15893_/X sky130_fd_sc_hd__a21o_1
XTAP_5496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17632_ _17632_/A vssd1 vssd1 vccd1 vccd1 _22704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_264_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14844_ _14855_/A vssd1 vssd1 vccd1 vccd1 _15538_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17563_ _17646_/S vssd1 vssd1 vccd1 vccd1 _17576_/S sky130_fd_sc_hd__buf_6
X_14775_ _15085_/S vssd1 vssd1 vccd1 vccd1 _15018_/S sky130_fd_sc_hd__clkbuf_4
X_11987_ _23316_/Q _23284_/Q _23252_/Q _23540_/Q _12709_/A _11669_/X vssd1 vssd1 vccd1
+ vccd1 _11987_/X sky130_fd_sc_hd__mux4_2
XFILLER_56_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19302_ _19324_/A vssd1 vssd1 vccd1 vccd1 _19311_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16514_ _16514_/A vssd1 vssd1 vccd1 vccd1 _22413_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13726_ _13726_/A vssd1 vssd1 vccd1 vccd1 _13726_/X sky130_fd_sc_hd__clkbuf_1
X_17494_ _22655_/Q _16236_/X _17494_/S vssd1 vssd1 vccd1 vccd1 _17495_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19233_ _19233_/A vssd1 vssd1 vccd1 vccd1 _19233_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_189_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16445_ _16013_/X _22383_/Q _16451_/S vssd1 vssd1 vccd1 vccd1 _16446_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13657_ _13657_/A vssd1 vssd1 vccd1 vccd1 _14069_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_319_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19164_ _19164_/A _19771_/B vssd1 vssd1 vccd1 vccd1 _19246_/A sky130_fd_sc_hd__or2_4
X_12608_ _13518_/A vssd1 vssd1 vccd1 vccd1 _13943_/A sky130_fd_sc_hd__buf_2
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_318_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16376_ _16376_/A vssd1 vssd1 vccd1 vccd1 _22353_/D sky130_fd_sc_hd__clkbuf_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13588_ _13588_/A vssd1 vssd1 vccd1 vccd1 _13884_/A sky130_fd_sc_hd__clkbuf_4
X_18115_ _18118_/A vssd1 vssd1 vccd1 vccd1 _18116_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_185_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15327_ _15327_/A vssd1 vssd1 vccd1 vccd1 _22271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19095_ _19095_/A vssd1 vssd1 vccd1 vccd1 _23237_/D sky130_fd_sc_hd__clkbuf_1
X_12539_ _22777_/Q _22745_/Q _22646_/Q _22713_/Q _23899_/Q _11189_/A vssd1 vssd1 vccd1
+ vccd1 _12539_/X sky130_fd_sc_hd__mux4_2
XFILLER_334_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18046_ _22853_/Q _18035_/X _18043_/X _18045_/X vssd1 vssd1 vccd1 vccd1 _22853_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15258_ _15248_/Y _15255_/X _15257_/X vssd1 vssd1 vccd1 vccd1 _15258_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_334_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14209_ _14526_/A _21287_/B vssd1 vssd1 vccd1 vccd1 _15618_/A sky130_fd_sc_hd__nor2_4
XFILLER_333_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_315_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15189_ _15189_/A _15432_/B vssd1 vssd1 vccd1 vccd1 _15189_/Y sky130_fd_sc_hd__nand2_2
XFILLER_99_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_342_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_174_wb_clk_i _23917_/CLK vssd1 vssd1 vccd1 vccd1 _23768_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19997_ _20009_/A _20009_/B vssd1 vssd1 vccd1 vccd1 _19998_/B sky130_fd_sc_hd__and2_1
XFILLER_301_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_103_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23456_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18948_ _19016_/S vssd1 vssd1 vccd1 vccd1 _18957_/S sky130_fd_sc_hd__buf_6
XFILLER_230_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18879_ _23142_/Q _18776_/X _18885_/S vssd1 vssd1 vccd1 vccd1 _18880_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20910_ _23785_/Q _20893_/X _20909_/X _20906_/X vssd1 vssd1 vccd1 vccd1 _23785_/D
+ sky130_fd_sc_hd__o211a_1
X_21890_ _23928_/Q _21890_/B vssd1 vssd1 vccd1 vccd1 _21890_/X sky130_fd_sc_hd__or2_1
XFILLER_55_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20841_ _20841_/A vssd1 vssd1 vccd1 vccd1 _23766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23560_ _23560_/CLK _23560_/D vssd1 vssd1 vccd1 vccd1 _23560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20772_ _20966_/A _20810_/A vssd1 vssd1 vccd1 vccd1 _20786_/B sky130_fd_sc_hd__or2_4
XFILLER_223_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_360 _23793_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_371 _23484_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22511_ _23693_/CLK _22511_/D vssd1 vssd1 vccd1 vccd1 _22511_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_382 _22490_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_393 _14090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23491_ _23491_/CLK _23491_/D vssd1 vssd1 vccd1 vccd1 _23491_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_357_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22442_ _23100_/CLK _22442_/D vssd1 vssd1 vccd1 vccd1 _22442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22373_ _23573_/CLK _22373_/D vssd1 vssd1 vccd1 vccd1 _22373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_337_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21324_ _21712_/S vssd1 vssd1 vccd1 vccd1 _21594_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_89_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_306_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21255_ _21258_/A _21255_/B vssd1 vssd1 vccd1 vccd1 _21256_/A sky130_fd_sc_hd__and2_2
XFILLER_296_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20206_ _20262_/A vssd1 vssd1 vccd1 vccd1 _20340_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21186_ _21281_/A vssd1 vssd1 vccd1 vccd1 _21186_/X sky130_fd_sc_hd__buf_6
XFILLER_132_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_292_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_292_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20137_ _20137_/A _20137_/B _20137_/C vssd1 vssd1 vccd1 vccd1 _23652_/D sky130_fd_sc_hd__nor3_1
XFILLER_131_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_293_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20068_ _20079_/B _20071_/C vssd1 vssd1 vccd1 vccd1 _20069_/B sky130_fd_sc_hd__and2_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_20 _17575_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_31 _18135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_42 _20713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _11910_/A vssd1 vssd1 vccd1 vccd1 _11911_/B sky130_fd_sc_hd__buf_2
XFILLER_46_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_53 _20678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_64 _21607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _11218_/A _12880_/X _12889_/X _11124_/A vssd1 vssd1 vccd1 vccd1 _12891_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_75 _21077_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_86 _14179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_97 _20303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11841_ _22786_/Q _22754_/Q _22655_/Q _22722_/Q _11148_/A _11840_/X vssd1 vssd1 vccd1
+ vccd1 _11841_/X sky130_fd_sc_hd__mux4_1
X_23827_ _23877_/CLK _23827_/D vssd1 vssd1 vccd1 vccd1 _23827_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _15976_/A vssd1 vssd1 vccd1 vccd1 _16198_/S sky130_fd_sc_hd__buf_6
X_11772_ _11905_/A _11772_/B vssd1 vssd1 vccd1 vccd1 _11772_/Y sky130_fd_sc_hd__nor2_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23758_ _23862_/CLK _23758_/D vssd1 vssd1 vccd1 vccd1 _23758_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_213_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _13906_/B _13511_/B _13334_/C _13334_/D vssd1 vssd1 vccd1 vccd1 _13935_/B
+ sky130_fd_sc_hd__or4bb_2
X_22709_ _23577_/CLK _22709_/D vssd1 vssd1 vccd1 vccd1 _22709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14491_ _14491_/A vssd1 vssd1 vccd1 vccd1 _15592_/A sky130_fd_sc_hd__buf_4
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23689_ _23696_/CLK _23689_/D vssd1 vssd1 vccd1 vccd1 _23689_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _18795_/A vssd1 vssd1 vccd1 vccd1 _16230_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_347_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13442_ _23888_/Q _23886_/Q _13442_/C vssd1 vssd1 vccd1 vccd1 _20532_/C sky130_fd_sc_hd__or3_2
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_356_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16161_ _19261_/A vssd1 vssd1 vccd1 vccd1 _16161_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13373_ _15122_/A _15122_/B _13370_/X _13372_/Y vssd1 vssd1 vccd1 vccd1 _13373_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_315_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15112_ _15112_/A _15111_/X vssd1 vssd1 vccd1 vccd1 _15113_/B sky130_fd_sc_hd__or2b_1
XFILLER_154_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_355_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12324_ _12324_/A vssd1 vssd1 vccd1 vccd1 _12324_/X sky130_fd_sc_hd__buf_4
X_16092_ _15575_/X _15432_/Y _15942_/X vssd1 vssd1 vccd1 vccd1 _21278_/A sky130_fd_sc_hd__a21oi_4
Xclkbuf_leaf_1_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23466_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_127_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19920_ _19922_/B _19915_/X _19916_/X _19919_/Y _18175_/X vssd1 vssd1 vccd1 vccd1
+ _23590_/D sky130_fd_sc_hd__a311oi_1
XFILLER_315_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15043_ _18788_/A vssd1 vssd1 vccd1 vccd1 _19181_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12255_ _22267_/Q _23083_/Q _23499_/Q _22428_/Q _12554_/S _11703_/A vssd1 vssd1 vccd1
+ vccd1 _12256_/B sky130_fd_sc_hd__mux4_1
XFILLER_142_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11206_ _13032_/S vssd1 vssd1 vccd1 vccd1 _11206_/X sky130_fd_sc_hd__buf_4
XFILLER_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19851_ _19851_/A vssd1 vssd1 vccd1 vccd1 _23559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12186_ _11138_/A _12181_/Y _12183_/Y _12185_/Y vssd1 vssd1 vccd1 vccd1 _12186_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_122_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11137_ _12534_/A vssd1 vssd1 vccd1 vccd1 _11138_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18802_ _23118_/Q _18801_/X _18802_/S vssd1 vssd1 vccd1 vccd1 _18803_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19782_ _23529_/Q _19178_/A _19782_/S vssd1 vssd1 vccd1 vccd1 _19783_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16994_ _17174_/B _16993_/X _16951_/A vssd1 vssd1 vccd1 vccd1 _16994_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18733_ _16863_/X _23092_/Q _18741_/S vssd1 vssd1 vccd1 vccd1 _18734_/A sky130_fd_sc_hd__mux2_1
XFILLER_284_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15945_ _13574_/A _14674_/X _15944_/X vssd1 vssd1 vccd1 vccd1 _15945_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11068_ _14814_/C vssd1 vssd1 vccd1 vccd1 _11068_/Y sky130_fd_sc_hd__inv_8
XTAP_5271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18664_ _18664_/A vssd1 vssd1 vccd1 vccd1 _23061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_264_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15876_ _23612_/Q vssd1 vssd1 vccd1 vccd1 _20009_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_236_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17615_ _22699_/Q _17614_/X _17624_/S vssd1 vssd1 vccd1 vccd1 _17616_/A sky130_fd_sc_hd__mux2_1
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14827_ input144/X input109/X _15030_/S vssd1 vssd1 vccd1 vccd1 _14827_/X sky130_fd_sc_hd__mux2_8
XFILLER_91_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18595_ _16873_/X _23031_/Q _18597_/S vssd1 vssd1 vccd1 vccd1 _18596_/A sky130_fd_sc_hd__mux2_1
XFILLER_251_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17546_ _17627_/A vssd1 vssd1 vccd1 vccd1 _17646_/S sky130_fd_sc_hd__buf_6
X_14758_ _16131_/B vssd1 vssd1 vccd1 vccd1 _15335_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_211_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13709_ _13709_/A vssd1 vssd1 vccd1 vccd1 _13721_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_204_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17477_ _22647_/Q _16211_/X _17483_/S vssd1 vssd1 vccd1 vccd1 _17478_/A sky130_fd_sc_hd__mux2_1
X_14689_ _14800_/A vssd1 vssd1 vccd1 vccd1 _14690_/A sky130_fd_sc_hd__buf_2
XFILLER_338_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19216_ _19216_/A vssd1 vssd1 vccd1 vccd1 _23284_/D sky130_fd_sc_hd__clkbuf_1
X_16428_ _16428_/A vssd1 vssd1 vccd1 vccd1 _22375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19147_ _19147_/A vssd1 vssd1 vccd1 vccd1 _23261_/D sky130_fd_sc_hd__clkbuf_1
X_16359_ _16359_/A vssd1 vssd1 vccd1 vccd1 _22345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_319_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_307_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19078_ _16899_/X _23231_/Q _19084_/S vssd1 vssd1 vccd1 vccd1 _19079_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_334_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18029_ _18029_/A vssd1 vssd1 vccd1 vccd1 _18029_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21040_ _20680_/A _21027_/X _21039_/X _21037_/X vssd1 vssd1 vccd1 vccd1 _23830_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_303_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22991_ _23009_/CLK _22991_/D vssd1 vssd1 vccd1 vccd1 _22991_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_227_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21942_ _21942_/A _21942_/B vssd1 vssd1 vccd1 vccd1 _21942_/Y sky130_fd_sc_hd__nor2_1
XFILLER_283_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21873_ _17180_/X _21867_/X _21872_/Y vssd1 vssd1 vccd1 vccd1 _21936_/B sky130_fd_sc_hd__a21o_1
XFILLER_83_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_71_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23548_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23612_ _23643_/CLK _23612_/D vssd1 vssd1 vccd1 vccd1 _23612_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20824_ _20658_/B _20810_/X _20811_/X _23762_/Q vssd1 vssd1 vccd1 vccd1 _20825_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_230_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23543_ _23543_/CLK _23543_/D vssd1 vssd1 vccd1 vccd1 _23543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_329_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20755_ _21076_/A _20724_/X _20733_/X vssd1 vssd1 vccd1 vccd1 _20755_/Y sky130_fd_sc_hd__a21oi_4
XINSDIODE2_190 _13931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23474_ _23474_/CLK _23474_/D vssd1 vssd1 vccd1 vccd1 _23474_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_196_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20686_ _21149_/A _20744_/B vssd1 vssd1 vccd1 vccd1 _20689_/B sky130_fd_sc_hd__nor2_4
XFILLER_183_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22425_ _23528_/CLK _22425_/D vssd1 vssd1 vccd1 vccd1 _22425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_353_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22356_ _23556_/CLK _22356_/D vssd1 vssd1 vccd1 vccd1 _22356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_352_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21307_ _21663_/A vssd1 vssd1 vccd1 vccd1 _21307_/X sky130_fd_sc_hd__clkbuf_4
X_22287_ _23551_/CLK _22287_/D vssd1 vssd1 vccd1 vccd1 _22287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_313_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12040_ _12754_/A _12040_/B vssd1 vssd1 vccd1 vccd1 _12040_/Y sky130_fd_sc_hd__nor2_1
X_21238_ _21238_/A _21240_/B vssd1 vssd1 vccd1 vccd1 _21238_/Y sky130_fd_sc_hd__nand2_1
XFILLER_340_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21169_ _20723_/A _21158_/X _21142_/X _20525_/B _21161_/X vssd1 vssd1 vccd1 vccd1
+ _21169_/X sky130_fd_sc_hd__a221o_1
XFILLER_172_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13991_ _13990_/A _13991_/B vssd1 vssd1 vccd1 vccd1 _13992_/A sky130_fd_sc_hd__and2b_1
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_322_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15730_ _23800_/Q _14603_/A _14918_/A vssd1 vssd1 vccd1 vccd1 _15730_/X sky130_fd_sc_hd__a21o_1
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12942_ _23931_/Q vssd1 vssd1 vccd1 vccd1 _15753_/A sky130_fd_sc_hd__clkinv_4
XFILLER_65_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _15923_/A _15661_/B vssd1 vssd1 vccd1 vccd1 _15661_/Y sky130_fd_sc_hd__nand2_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _22475_/Q _22635_/Q _12978_/S vssd1 vssd1 vccd1 vccd1 _12873_/X sky130_fd_sc_hd__mux2_1
XFILLER_234_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _17456_/A vssd1 vssd1 vccd1 vccd1 _17469_/S sky130_fd_sc_hd__buf_6
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _15222_/A vssd1 vssd1 vccd1 vccd1 _14612_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_324_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18380_ _18423_/A vssd1 vssd1 vccd1 vccd1 _18380_/X sky130_fd_sc_hd__buf_4
X_11824_ _12318_/A _11824_/B vssd1 vssd1 vccd1 vccd1 _11824_/X sky130_fd_sc_hd__or2_1
XFILLER_27_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _15592_/A vssd1 vssd1 vccd1 vccd1 _15592_/X sky130_fd_sc_hd__buf_4
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_324_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _22588_/Q input201/X _17335_/S vssd1 vssd1 vccd1 vccd1 _17332_/A sky130_fd_sc_hd__mux2_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14543_ _15618_/A _21294_/B vssd1 vssd1 vccd1 vccd1 _14543_/X sky130_fd_sc_hd__or2_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11755_ _11755_/A vssd1 vssd1 vccd1 vccd1 _12025_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17262_ _17262_/A vssd1 vssd1 vccd1 vccd1 _17262_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_202_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_348_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14474_ _14474_/A vssd1 vssd1 vccd1 vccd1 _21097_/A sky130_fd_sc_hd__inv_4
XFILLER_159_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11686_ _12283_/B vssd1 vssd1 vccd1 vccd1 _11935_/B sky130_fd_sc_hd__clkbuf_8
X_19001_ _16892_/X _23197_/Q _19001_/S vssd1 vssd1 vccd1 vccd1 _19002_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16213_ _16213_/A vssd1 vssd1 vccd1 vccd1 _22294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13425_ _15425_/A _13470_/A vssd1 vssd1 vccd1 vccd1 _14250_/A sky130_fd_sc_hd__nor2_4
X_17193_ _11483_/X _17192_/X _17234_/S vssd1 vssd1 vccd1 vccd1 _17193_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16144_ _22976_/Q _16143_/X _16144_/S vssd1 vssd1 vccd1 vccd1 _16144_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13356_ _13356_/A _13906_/A vssd1 vssd1 vccd1 vccd1 _14940_/A sky130_fd_sc_hd__xnor2_1
XFILLER_128_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12307_ _12307_/A _12307_/B vssd1 vssd1 vccd1 vccd1 _12307_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16075_ _23939_/Q vssd1 vssd1 vccd1 vccd1 _22165_/A sky130_fd_sc_hd__clkbuf_2
X_13287_ _13287_/A _13287_/B vssd1 vssd1 vccd1 vccd1 _13287_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19903_ _16291_/X _23583_/Q _19909_/S vssd1 vssd1 vccd1 vccd1 _19904_/A sky130_fd_sc_hd__mux2_1
X_15026_ input164/X input128/X _15057_/S vssd1 vssd1 vccd1 vccd1 _15026_/X sky130_fd_sc_hd__mux2_8
XFILLER_269_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12238_ _22363_/Q _22395_/Q _22684_/Q _23051_/Q _11414_/A _12199_/X vssd1 vssd1 vccd1
+ vccd1 _12239_/B sky130_fd_sc_hd__mux4_1
XFILLER_107_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_331_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_300_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_297_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19834_ _19834_/A vssd1 vssd1 vccd1 vccd1 _23552_/D sky130_fd_sc_hd__clkbuf_1
X_12169_ _13351_/A _12167_/Y _12168_/Y vssd1 vssd1 vccd1 vccd1 _12169_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_311_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19765_ _19258_/X _23522_/Q _19765_/S vssd1 vssd1 vccd1 vccd1 _19766_/A sky130_fd_sc_hd__mux2_1
X_16977_ _22711_/Q vssd1 vssd1 vccd1 vccd1 _21301_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_56_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_300_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 coreIndex[4] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18716_ _18716_/A vssd1 vssd1 vccd1 vccd1 _23084_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15928_ _15479_/A _13581_/B _15923_/X _15927_/X _15375_/X vssd1 vssd1 vccd1 vccd1
+ _15928_/X sky130_fd_sc_hd__a221o_2
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19696_ _19696_/A vssd1 vssd1 vccd1 vccd1 _23491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18647_ _23054_/Q _17575_/X _18647_/S vssd1 vssd1 vccd1 vccd1 _18648_/A sky130_fd_sc_hd__mux2_1
X_15859_ _15857_/X _22003_/A _16047_/S vssd1 vssd1 vccd1 vccd1 _18843_/A sky130_fd_sc_hd__mux2_8
XFILLER_52_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18578_ _16847_/X _23023_/Q _18586_/S vssd1 vssd1 vccd1 vccd1 _18579_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17529_ _17529_/A vssd1 vssd1 vccd1 vccd1 _17538_/S sky130_fd_sc_hd__buf_6
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20540_ _14468_/B _20890_/B _21301_/C vssd1 vssd1 vccd1 vccd1 _20729_/A sky130_fd_sc_hd__o21ai_4
XFILLER_193_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20471_ _23707_/Q _20487_/B vssd1 vssd1 vccd1 vccd1 _20471_/X sky130_fd_sc_hd__or2_1
XFILLER_335_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22210_ _23843_/Q _23777_/Q vssd1 vssd1 vccd1 vccd1 _22210_/X sky130_fd_sc_hd__or2_1
XFILLER_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23190_ _23573_/CLK _23190_/D vssd1 vssd1 vccd1 vccd1 _23190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_307_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22141_ _22115_/A _22118_/B _22114_/Y vssd1 vssd1 vccd1 vccd1 _22142_/C sky130_fd_sc_hd__o21ai_1
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_350_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput320 _13982_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[25] sky130_fd_sc_hd__buf_2
Xoutput331 _16680_/A vssd1 vssd1 vccd1 vccd1 core_wb_cyc_o sky130_fd_sc_hd__buf_2
Xoutput342 _13807_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[19] sky130_fd_sc_hd__buf_2
XFILLER_133_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput353 _13867_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[29] sky130_fd_sc_hd__buf_2
X_22072_ _22053_/A _22155_/A _22052_/A vssd1 vssd1 vccd1 vccd1 _22076_/A sky130_fd_sc_hd__a21bo_1
XTAP_6719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_288_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput364 _13880_/Y vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[0] sky130_fd_sc_hd__buf_2
XFILLER_236_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput375 _14029_/X vssd1 vssd1 vccd1 vccd1 din0[10] sky130_fd_sc_hd__buf_2
XFILLER_87_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput386 _14048_/X vssd1 vssd1 vccd1 vccd1 din0[20] sky130_fd_sc_hd__buf_2
X_21023_ _21023_/A vssd1 vssd1 vccd1 vccd1 _21023_/X sky130_fd_sc_hd__buf_2
Xoutput397 _14068_/X vssd1 vssd1 vccd1 vccd1 din0[30] sky130_fd_sc_hd__buf_2
XFILLER_259_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_302_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22974_ _22974_/CLK _22974_/D vssd1 vssd1 vccd1 vccd1 _22974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_290_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21925_ _21925_/A vssd1 vssd1 vccd1 vccd1 _22012_/A sky130_fd_sc_hd__inv_2
XFILLER_347_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21856_ _21856_/A _21861_/A vssd1 vssd1 vccd1 vccd1 _21856_/Y sky130_fd_sc_hd__nor2_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_358_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20807_ _20807_/A vssd1 vssd1 vccd1 vccd1 _23757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21787_ _21787_/A _21787_/B vssd1 vssd1 vccd1 vccd1 _21787_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_230_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_329_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11540_ _23234_/Q _23202_/Q _23170_/Q _23138_/Q _11517_/X _11519_/X vssd1 vssd1 vccd1
+ vccd1 _11541_/B sky130_fd_sc_hd__mux4_1
X_23526_ _23526_/CLK _23526_/D vssd1 vssd1 vccd1 vccd1 _23526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20738_ _23742_/Q _20729_/X _20736_/X _20737_/X vssd1 vssd1 vccd1 vccd1 _23742_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_345_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11471_ _21848_/A _11471_/B vssd1 vssd1 vccd1 vccd1 _11471_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23457_ _23553_/CLK _23457_/D vssd1 vssd1 vccd1 vccd1 _23457_/Q sky130_fd_sc_hd__dfxtp_1
X_20669_ _21033_/A _20669_/B vssd1 vssd1 vccd1 vccd1 _20672_/B sky130_fd_sc_hd__nor2_8
XFILLER_137_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13210_ _13210_/A _13210_/B vssd1 vssd1 vccd1 vccd1 _13210_/Y sky130_fd_sc_hd__nor2_1
X_22408_ _23450_/CLK _22408_/D vssd1 vssd1 vccd1 vccd1 _22408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14190_ _21555_/A _21443_/A vssd1 vssd1 vccd1 vccd1 _14564_/A sky130_fd_sc_hd__nand2_2
X_23388_ _23420_/CLK _23388_/D vssd1 vssd1 vccd1 vccd1 _23388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_303_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13141_ _23904_/Q vssd1 vssd1 vccd1 vccd1 _21448_/B sky130_fd_sc_hd__buf_8
X_22339_ _23505_/CLK _22339_/D vssd1 vssd1 vccd1 vccd1 _22339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_325_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_297_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_340_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13072_ _22804_/Q _22772_/Q _22673_/Q _22740_/Q _11517_/X _11519_/X vssd1 vssd1 vccd1
+ vccd1 _13073_/B sky130_fd_sc_hd__mux4_1
XFILLER_124_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16900_ _16899_/X _22547_/Q _16909_/S vssd1 vssd1 vccd1 vccd1 _16901_/A sky130_fd_sc_hd__mux2_1
XFILLER_300_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12023_ _12011_/Y _12016_/Y _12019_/Y _12022_/Y _11683_/X vssd1 vssd1 vccd1 vccd1
+ _12037_/B sky130_fd_sc_hd__o221a_1
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17880_ _22811_/Q input249/X _17882_/S vssd1 vssd1 vccd1 vccd1 _17881_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16831_ _19181_/A vssd1 vssd1 vccd1 vccd1 _16831_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_266_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19550_ _19550_/A vssd1 vssd1 vccd1 vccd1 _23426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_293_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16762_ _22506_/Q _16747_/X _16748_/X input20/X vssd1 vssd1 vccd1 vccd1 _16763_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_207_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13974_ _13974_/A _13974_/B vssd1 vssd1 vccd1 vccd1 _13974_/Y sky130_fd_sc_hd__nor2_1
XFILLER_219_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18501_ _18494_/X _18500_/Y _18490_/X vssd1 vssd1 vccd1 vccd1 _22995_/D sky130_fd_sc_hd__a21oi_1
XFILLER_47_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15713_ _23930_/Q _21868_/B vssd1 vssd1 vccd1 vccd1 _15790_/C sky130_fd_sc_hd__and2_2
XFILLER_74_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12925_ _23225_/Q _23193_/Q _23161_/Q _23129_/Q _12819_/S _11166_/A vssd1 vssd1 vccd1
+ vccd1 _12926_/B sky130_fd_sc_hd__mux4_2
X_19481_ _23396_/Q _18871_/X _19481_/S vssd1 vssd1 vccd1 vccd1 _19482_/A sky130_fd_sc_hd__mux2_1
X_16693_ _16730_/A vssd1 vssd1 vccd1 vccd1 _16693_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18432_ _18435_/A _18435_/C _18423_/X vssd1 vssd1 vccd1 vccd1 _18432_/Y sky130_fd_sc_hd__a21oi_1
X_15644_ _15644_/A _15835_/B vssd1 vssd1 vccd1 vccd1 _15644_/X sky130_fd_sc_hd__or2_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _12897_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _12856_/X sky130_fd_sc_hd__or2_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _14729_/X _18366_/C _18362_/Y vssd1 vssd1 vccd1 vccd1 _22948_/D sky130_fd_sc_hd__o21a_1
XFILLER_221_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11807_ _22787_/Q _22755_/Q _22656_/Q _22723_/Q _11648_/A _11653_/A vssd1 vssd1 vccd1
+ vccd1 _11808_/B sky130_fd_sc_hd__mux4_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _15901_/A vssd1 vssd1 vccd1 vccd1 _15575_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _12779_/Y _12782_/Y _12784_/Y _12786_/Y _11276_/A vssd1 vssd1 vccd1 vccd1
+ _12800_/B sky130_fd_sc_hd__o221a_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_348_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17314_ input102/X input67/X _17314_/S vssd1 vssd1 vccd1 vccd1 _17314_/X sky130_fd_sc_hd__mux2_8
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _14526_/A _21287_/B vssd1 vssd1 vccd1 vccd1 _14539_/S sky130_fd_sc_hd__or2_4
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_309_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18294_ _18296_/A _18296_/C _18293_/Y vssd1 vssd1 vccd1 vccd1 _22924_/D sky130_fd_sc_hd__o21a_1
XFILLER_230_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11738_ _23408_/Q _23024_/Q _23376_/Q _23344_/Q _12024_/A _12014_/A vssd1 vssd1 vccd1
+ vccd1 _11738_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_348_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17245_ _17245_/A vssd1 vssd1 vccd1 vccd1 _17245_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14457_ _14457_/A _14404_/B vssd1 vssd1 vccd1 vccd1 _20989_/A sky130_fd_sc_hd__or2b_2
X_11669_ _11676_/A vssd1 vssd1 vccd1 vccd1 _11669_/X sky130_fd_sc_hd__buf_6
XFILLER_175_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13408_ _13574_/A _13408_/B vssd1 vssd1 vccd1 vccd1 _13408_/Y sky130_fd_sc_hd__xnor2_2
X_17176_ _17237_/A vssd1 vssd1 vccd1 vccd1 _17176_/X sky130_fd_sc_hd__clkbuf_2
X_14388_ _14675_/A _20305_/A _14388_/C vssd1 vssd1 vccd1 vccd1 _14389_/C sky130_fd_sc_hd__or3_1
XFILLER_127_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_317_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16127_ _15575_/X _15484_/Y _15942_/X vssd1 vssd1 vccd1 vccd1 _21280_/A sky130_fd_sc_hd__a21oi_4
XFILLER_343_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_332_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13339_ _13343_/B _13380_/A _13382_/B _13338_/Y _11945_/X vssd1 vssd1 vccd1 vccd1
+ _13344_/B sky130_fd_sc_hd__o311ai_2
XFILLER_289_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_332_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16058_ _15636_/X _16053_/X _16056_/X _16057_/X vssd1 vssd1 vccd1 vccd1 _16058_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_288_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15009_ _13370_/D _13913_/Y _15867_/S vssd1 vssd1 vccd1 vccd1 _15010_/B sky130_fd_sc_hd__mux2_1
XFILLER_124_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_312_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_300_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19817_ _19828_/A vssd1 vssd1 vccd1 vccd1 _19826_/S sky130_fd_sc_hd__buf_4
XFILLER_243_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_300_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19748_ _19233_/X _23514_/Q _19754_/S vssd1 vssd1 vccd1 vccd1 _19749_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19679_ _19679_/A vssd1 vssd1 vccd1 vccd1 _23483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21710_ _21675_/A _21675_/B _21674_/A vssd1 vssd1 vccd1 vccd1 _21711_/B sky130_fd_sc_hd__a21o_1
XFILLER_64_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22690_ _22789_/CLK _22690_/D vssd1 vssd1 vccd1 vccd1 _22690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21641_ _21641_/A _22091_/B vssd1 vssd1 vccd1 vccd1 _21641_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21572_ _21572_/A _21572_/B vssd1 vssd1 vccd1 vccd1 _21574_/A sky130_fd_sc_hd__nor2_1
XFILLER_123_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_339_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23311_ _23535_/CLK _23311_/D vssd1 vssd1 vccd1 vccd1 _23311_/Q sky130_fd_sc_hd__dfxtp_1
X_20523_ _23702_/Q _20523_/B _20523_/C vssd1 vssd1 vccd1 vccd1 _20525_/C sky130_fd_sc_hd__and3_1
XFILLER_138_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_355_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20454_ _23700_/Q _20413_/X _20453_/Y _20445_/X vssd1 vssd1 vccd1 vccd1 _23700_/D
+ sky130_fd_sc_hd__o211a_1
X_23242_ _23370_/CLK _23242_/D vssd1 vssd1 vccd1 vccd1 _23242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23173_ _23493_/CLK _23173_/D vssd1 vssd1 vccd1 vccd1 _23173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20385_ _23681_/Q _20391_/B vssd1 vssd1 vccd1 vccd1 _20385_/X sky130_fd_sc_hd__or2_1
XTAP_7206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_334_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22124_ _22155_/C _22104_/B _22101_/A vssd1 vssd1 vccd1 vccd1 _22128_/A sky130_fd_sc_hd__a21oi_1
XFILLER_350_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22055_ _23837_/Q _23771_/Q vssd1 vssd1 vccd1 vccd1 _22057_/A sky130_fd_sc_hd__and2_1
XTAP_6549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_288_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21006_ _23818_/Q _21009_/B vssd1 vssd1 vccd1 vccd1 _21006_/X sky130_fd_sc_hd__or2_1
XFILLER_287_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_303_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22957_ _22961_/CLK _22957_/D vssd1 vssd1 vccd1 vccd1 _22957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_290_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12710_ _12710_/A vssd1 vssd1 vccd1 vccd1 _12710_/X sky130_fd_sc_hd__clkbuf_4
X_21908_ _21346_/A _21907_/X _21683_/A _23800_/Q vssd1 vssd1 vccd1 vccd1 _21908_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_244_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13690_ _14219_/A vssd1 vssd1 vccd1 vccd1 _13691_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22888_ _23551_/CLK _22888_/D vssd1 vssd1 vccd1 vccd1 _22888_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_270_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_349_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12641_ _12637_/X _12638_/X _12640_/X vssd1 vssd1 vccd1 vccd1 _12641_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_203_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21839_ _23830_/Q _21418_/A _21838_/Y _21377_/X vssd1 vssd1 vccd1 vccd1 _21839_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15360_ _15360_/A _15360_/B vssd1 vssd1 vccd1 vccd1 _15360_/Y sky130_fd_sc_hd__nand2_1
XFILLER_157_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12572_ _11230_/A _12565_/X _12567_/X _12571_/X _11215_/A vssd1 vssd1 vccd1 vccd1
+ _13718_/C sky130_fd_sc_hd__a311o_4
XPHY_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14311_ _14306_/X _14310_/X _14639_/A vssd1 vssd1 vccd1 vccd1 _14311_/X sky130_fd_sc_hd__mux2_1
XFILLER_346_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23509_ _23541_/CLK _23509_/D vssd1 vssd1 vccd1 vccd1 _23509_/Q sky130_fd_sc_hd__dfxtp_1
X_11523_ _13218_/A vssd1 vssd1 vccd1 vccd1 _13073_/A sky130_fd_sc_hd__buf_2
XFILLER_184_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15291_ _14784_/Y _14779_/Y _15490_/S vssd1 vssd1 vccd1 vccd1 _15291_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17030_ _23465_/Q _16987_/X _16988_/X _16989_/X _14939_/B vssd1 vssd1 vccd1 vccd1
+ _17030_/X sky130_fd_sc_hd__a32o_1
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14242_ _15179_/A vssd1 vssd1 vccd1 vccd1 _14242_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_109_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11454_ _11821_/A vssd1 vssd1 vccd1 vccd1 _11455_/A sky130_fd_sc_hd__buf_4
XFILLER_125_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11385_ _12415_/S vssd1 vssd1 vccd1 vccd1 _11828_/B sky130_fd_sc_hd__buf_2
X_14173_ _14815_/C _14524_/B vssd1 vssd1 vccd1 vccd1 _14198_/C sky130_fd_sc_hd__nand2_1
XFILLER_313_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_314_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13124_ _11537_/X _13117_/Y _13119_/Y _13121_/Y _13123_/Y vssd1 vssd1 vccd1 vccd1
+ _13124_/X sky130_fd_sc_hd__o32a_1
XFILLER_124_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18981_ _19003_/A vssd1 vssd1 vccd1 vccd1 _18990_/S sky130_fd_sc_hd__buf_4
XFILLER_298_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17932_ _17932_/A vssd1 vssd1 vccd1 vccd1 _17932_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13055_ _11219_/A _13044_/X _13054_/X _13210_/A vssd1 vssd1 vccd1 vccd1 _13056_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_279_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12006_ _13531_/A _12005_/Y vssd1 vssd1 vccd1 vccd1 _13615_/A sky130_fd_sc_hd__nor2b_4
X_17863_ _17863_/A vssd1 vssd1 vccd1 vccd1 _22802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_294_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19602_ _23449_/Q _19229_/A _19610_/S vssd1 vssd1 vccd1 vccd1 _19603_/A sky130_fd_sc_hd__mux2_1
XFILLER_226_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16814_ _19699_/B _19843_/A vssd1 vssd1 vccd1 vccd1 _16896_/A sky130_fd_sc_hd__or2_4
XFILLER_120_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17794_ _22772_/Q _17633_/X _17798_/S vssd1 vssd1 vccd1 vccd1 _17795_/A sky130_fd_sc_hd__mux2_1
XFILLER_226_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19533_ _19533_/A vssd1 vssd1 vccd1 vccd1 _23418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16745_ _16759_/A _16745_/B vssd1 vssd1 vccd1 vccd1 _16746_/A sky130_fd_sc_hd__or2_1
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13957_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13957_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_253_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_199_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23368_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19464_ _23388_/Q _18846_/X _19466_/S vssd1 vssd1 vccd1 vccd1 _19465_/A sky130_fd_sc_hd__mux2_1
X_12908_ _23418_/Q _23034_/Q _23386_/Q _23354_/Q _12709_/A _11669_/X vssd1 vssd1 vccd1
+ vccd1 _12909_/B sky130_fd_sc_hd__mux4_2
XFILLER_234_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16676_ _16676_/A vssd1 vssd1 vccd1 vccd1 _22484_/D sky130_fd_sc_hd__clkbuf_1
X_13888_ _13967_/B _13888_/B vssd1 vssd1 vccd1 vccd1 _13889_/A sky130_fd_sc_hd__and2_4
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_128_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23651_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_234_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15627_ _15627_/A vssd1 vssd1 vccd1 vccd1 _22277_/D sky130_fd_sc_hd__clkbuf_1
X_18415_ _18418_/A _18418_/C _18380_/X vssd1 vssd1 vccd1 vccd1 _18415_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19395_ _19395_/A vssd1 vssd1 vccd1 vccd1 _23357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12839_ _12891_/A _12839_/B vssd1 vssd1 vccd1 vccd1 _12839_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18346_ _16059_/X _18349_/C _18337_/X vssd1 vssd1 vccd1 vccd1 _18346_/Y sky130_fd_sc_hd__a21oi_1
X_15558_ _15558_/A vssd1 vssd1 vccd1 vccd1 _15558_/X sky130_fd_sc_hd__buf_2
XFILLER_203_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_349_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14509_ _14509_/A vssd1 vssd1 vccd1 vccd1 _14509_/X sky130_fd_sc_hd__buf_2
XFILLER_202_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18277_ _18277_/A vssd1 vssd1 vccd1 vccd1 _19962_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_148_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15489_ _15020_/S _15488_/Y _14630_/X vssd1 vssd1 vccd1 vccd1 _15489_/X sky130_fd_sc_hd__a21o_1
XFILLER_336_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_308_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17228_ input93/X input58/X _17266_/S vssd1 vssd1 vccd1 vccd1 _17228_/X sky130_fd_sc_hd__mux2_8
XFILLER_147_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput30 core_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput41 core_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_1
XFILLER_337_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput52 dout0[18] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_2
XFILLER_174_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput63 dout0[28] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__buf_2
XFILLER_351_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17159_ _17159_/A _17172_/B vssd1 vssd1 vccd1 vccd1 _17159_/Y sky130_fd_sc_hd__nor2_1
Xinput74 dout0[38] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__clkbuf_1
XFILLER_337_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput85 dout0[48] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput96 dout0[58] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_5_0_wb_clk_i INSDIODE2_358/DIODE vssd1 vssd1 vccd1 vccd1 _23917_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_304_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20170_ _20197_/S vssd1 vssd1 vccd1 vccd1 _20394_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23860_ _23861_/CLK _23860_/D vssd1 vssd1 vccd1 vccd1 _23860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22811_ _22968_/CLK _22811_/D vssd1 vssd1 vccd1 vccd1 _22811_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23791_ _23861_/CLK _23791_/D vssd1 vssd1 vccd1 vccd1 _23791_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_344_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22742_ _23586_/CLK _22742_/D vssd1 vssd1 vccd1 vccd1 _22742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_344_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22673_ _23456_/CLK _22673_/D vssd1 vssd1 vccd1 vccd1 _22673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21624_ _21624_/A _21624_/B _21624_/C vssd1 vssd1 vccd1 vccd1 _21625_/B sky130_fd_sc_hd__or3_1
XFILLER_139_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_328_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_328_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21555_ _21555_/A vssd1 vssd1 vccd1 vccd1 _21865_/A sky130_fd_sc_hd__buf_2
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_355_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20506_ _23711_/Q _20508_/B _20506_/C vssd1 vssd1 vccd1 vccd1 _20509_/B sky130_fd_sc_hd__and3_1
XFILLER_327_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_315_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21486_ _21543_/C _21454_/B _21451_/B vssd1 vssd1 vccd1 vccd1 _21487_/B sky130_fd_sc_hd__a21oi_2
XFILLER_355_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_354_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23225_ _23419_/CLK _23225_/D vssd1 vssd1 vccd1 vccd1 _23225_/Q sky130_fd_sc_hd__dfxtp_1
X_20437_ _20615_/A _20428_/X _20436_/X _20433_/X vssd1 vssd1 vccd1 vccd1 _23693_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_307_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11170_ _11200_/A vssd1 vssd1 vccd1 vccd1 _11170_/X sky130_fd_sc_hd__buf_2
X_23156_ _23543_/CLK _23156_/D vssd1 vssd1 vccd1 vccd1 _23156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_351_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20368_ _20368_/A _20368_/B vssd1 vssd1 vccd1 vccd1 _20368_/X sky130_fd_sc_hd__or2_1
XFILLER_351_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22107_ _23839_/Q _23773_/Q vssd1 vssd1 vccd1 vccd1 _22109_/A sky130_fd_sc_hd__nor2_1
XTAP_7069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23087_ _23535_/CLK _23087_/D vssd1 vssd1 vccd1 vccd1 _23087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20299_ _20294_/X _21829_/A _20297_/Y _20298_/X vssd1 vssd1 vccd1 vccd1 _20675_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_314_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22038_ _22038_/A _22038_/B _22038_/C vssd1 vssd1 vccd1 vccd1 _22040_/B sky130_fd_sc_hd__and3_1
XTAP_6379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14860_ _15253_/A vssd1 vssd1 vccd1 vccd1 _14860_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ _13736_/B _13758_/X _13809_/X _13857_/B vssd1 vssd1 vccd1 vccd1 _13812_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_235_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14791_ _14791_/A _15018_/S vssd1 vssd1 vccd1 vccd1 _14794_/B sky130_fd_sc_hd__nand2_1
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_290_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16530_ _16530_/A vssd1 vssd1 vccd1 vccd1 _17382_/A sky130_fd_sc_hd__buf_12
XFILLER_44_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13742_ _13742_/A vssd1 vssd1 vccd1 vccd1 _13742_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16461_ _14534_/X _22389_/Q _16469_/S vssd1 vssd1 vccd1 vccd1 _16462_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13673_ _13651_/B _14001_/A _14080_/A _22598_/Q vssd1 vssd1 vccd1 vccd1 _17039_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18200_ _18549_/A _18536_/A _23010_/Q vssd1 vssd1 vccd1 vccd1 _18203_/C sky130_fd_sc_hd__or3_2
XFILLER_32_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15412_ _16191_/A _15412_/B vssd1 vssd1 vccd1 vccd1 _15412_/X sky130_fd_sc_hd__or2_1
X_12624_ _12616_/Y _12618_/Y _12621_/Y _12623_/Y _11683_/X vssd1 vssd1 vccd1 vccd1
+ _12634_/B sky130_fd_sc_hd__o221a_2
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19180_ _19180_/A vssd1 vssd1 vccd1 vccd1 _23273_/D sky130_fd_sc_hd__clkbuf_1
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16392_ _14811_/X _22359_/Q _16396_/S vssd1 vssd1 vccd1 vccd1 _16393_/A sky130_fd_sc_hd__mux2_1
XPHY_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_346_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18131_ _18116_/Y _18129_/X _18130_/X _18121_/X vssd1 vssd1 vccd1 vccd1 _22881_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15343_ _14839_/A _15341_/X _15342_/X vssd1 vssd1 vccd1 vccd1 _15343_/X sky130_fd_sc_hd__o21a_1
XPHY_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12555_ _12556_/A vssd1 vssd1 vccd1 vccd1 _13455_/A sky130_fd_sc_hd__clkinv_8
XFILLER_345_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18062_ hold8/A _18052_/X _18053_/X _22991_/Q _18054_/X vssd1 vssd1 vccd1 vccd1 _18062_/X
+ sky130_fd_sc_hd__a221o_1
X_11506_ _13268_/A _11506_/B vssd1 vssd1 vccd1 vccd1 _11506_/Y sky130_fd_sc_hd__nor2_1
X_15274_ _23920_/Q _23919_/Q _15274_/C vssd1 vssd1 vccd1 vccd1 _15316_/B sky130_fd_sc_hd__and3_1
XFILLER_184_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12486_ _23206_/Q _23174_/Q _23142_/Q _23110_/Q _12475_/X _12476_/X vssd1 vssd1 vccd1
+ vccd1 _12486_/X sky130_fd_sc_hd__mux4_2
X_17013_ _17000_/X _17001_/X _17011_/X _17012_/X vssd1 vssd1 vccd1 vccd1 _17013_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_305_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14225_ _15110_/S vssd1 vssd1 vccd1 vccd1 _15114_/S sky130_fd_sc_hd__buf_2
XFILLER_156_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11437_ _11497_/A _11437_/B vssd1 vssd1 vccd1 vccd1 _11437_/X sky130_fd_sc_hd__or2_1
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14156_ _16941_/B _16941_/A _14415_/S vssd1 vssd1 vccd1 vccd1 _16949_/A sky130_fd_sc_hd__and3b_1
XFILLER_152_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_342_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_298_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11368_ _23492_/Q _23588_/Q _22552_/Q _22356_/Q _11461_/A _11365_/X vssd1 vssd1 vccd1
+ vccd1 _11369_/B sky130_fd_sc_hd__mux4_1
XFILLER_125_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_313_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13107_ _13107_/A _13107_/B vssd1 vssd1 vccd1 vccd1 _13107_/Y sky130_fd_sc_hd__nor2_1
XFILLER_298_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14087_ _14087_/A vssd1 vssd1 vccd1 vccd1 _14087_/Y sky130_fd_sc_hd__inv_2
X_18964_ _16838_/X _23180_/Q _18968_/S vssd1 vssd1 vccd1 vccd1 _18965_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11299_ _13121_/A vssd1 vssd1 vccd1 vccd1 _11343_/A sky130_fd_sc_hd__buf_4
XFILLER_26_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17915_ _17933_/A vssd1 vssd1 vccd1 vccd1 _17915_/X sky130_fd_sc_hd__clkbuf_2
X_13038_ _22804_/Q _22772_/Q _22673_/Q _22740_/Q _11432_/A _13037_/X vssd1 vssd1 vccd1
+ vccd1 _13039_/B sky130_fd_sc_hd__mux4_1
XFILLER_224_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18895_ _18895_/A vssd1 vssd1 vccd1 vccd1 _23149_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17846_ _22795_/Q _17604_/X _17848_/S vssd1 vssd1 vccd1 vccd1 _17847_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14989_ _22951_/Q vssd1 vssd1 vccd1 vccd1 _14989_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_281_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17777_ _17777_/A vssd1 vssd1 vccd1 vccd1 _22764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19516_ _19210_/X _23411_/Q _19516_/S vssd1 vssd1 vccd1 vccd1 _19517_/A sky130_fd_sc_hd__mux2_1
XFILLER_263_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16728_ _16728_/A vssd1 vssd1 vccd1 vccd1 _22496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_520 _13883_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_531 _14127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_542 _23946_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19447_ _23380_/Q _18820_/X _19455_/S vssd1 vssd1 vccd1 vccd1 _19448_/A sky130_fd_sc_hd__mux2_1
X_16659_ _16659_/A vssd1 vssd1 vccd1 vccd1 _22476_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_553 _13679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_320_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_564 _21871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19378_ _19378_/A vssd1 vssd1 vccd1 vccd1 _23349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_349_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_309_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18329_ _15833_/X _18332_/C _18292_/X vssd1 vssd1 vccd1 vccd1 _18329_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_194_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_336_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21340_ _21340_/A _21615_/A vssd1 vssd1 vccd1 vccd1 _21340_/X sky130_fd_sc_hd__and2_1
XFILLER_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_96_wb_clk_i _22899_/CLK vssd1 vssd1 vccd1 vccd1 _23554_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_135_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21271_ _21078_/B _21242_/X _21269_/Y _21270_/X vssd1 vssd1 vccd1 vccd1 _23904_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_351_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_25_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23459_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_333_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23010_ _23599_/CLK _23010_/D vssd1 vssd1 vccd1 vccd1 _23010_/Q sky130_fd_sc_hd__dfxtp_2
X_20222_ _20192_/X _21500_/B _20218_/Y _20221_/X vssd1 vssd1 vccd1 vccd1 _20604_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_305_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_304_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_305_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_304_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20153_ _20214_/A _20214_/B vssd1 vssd1 vccd1 vccd1 _20168_/A sky130_fd_sc_hd__or2_1
XFILLER_320_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_350_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_320_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20084_ _20090_/C _20090_/D _23636_/Q vssd1 vssd1 vccd1 vccd1 _20086_/B sky130_fd_sc_hd__a21oi_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23912_ _23916_/CLK _23912_/D vssd1 vssd1 vccd1 vccd1 _23912_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23843_ _23876_/CLK _23843_/D vssd1 vssd1 vccd1 vccd1 _23843_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23774_ _23776_/CLK _23774_/D vssd1 vssd1 vccd1 vccd1 _23774_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20986_ _20986_/A _20986_/B vssd1 vssd1 vccd1 vccd1 _21047_/A sky130_fd_sc_hd__or2_4
XFILLER_53_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22725_ _22789_/CLK _22725_/D vssd1 vssd1 vccd1 vccd1 _22725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22656_ _23567_/CLK _22656_/D vssd1 vssd1 vccd1 vccd1 _22656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_328_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_327_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21607_ _21690_/B _21614_/B vssd1 vssd1 vccd1 vccd1 _21607_/X sky130_fd_sc_hd__xor2_4
XFILLER_279_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22587_ _22968_/CLK _22587_/D vssd1 vssd1 vccd1 vccd1 _22587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12340_ _13514_/A _12340_/B vssd1 vssd1 vccd1 vccd1 _13334_/C sky130_fd_sc_hd__xnor2_1
XFILLER_343_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21538_ _21663_/A _21529_/X _21537_/X _21361_/A _21479_/A vssd1 vssd1 vccd1 vccd1
+ _21538_/X sky130_fd_sc_hd__o221a_1
XFILLER_126_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_315_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12271_ _12397_/A _12270_/X _11819_/X vssd1 vssd1 vccd1 vccd1 _12271_/Y sky130_fd_sc_hd__o21ai_1
X_21469_ _23916_/Q _21474_/A vssd1 vssd1 vccd1 vccd1 _21470_/B sky130_fd_sc_hd__nand2_1
XFILLER_182_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _13715_/A _14083_/A _13793_/B _14009_/X input226/X vssd1 vssd1 vccd1 vccd1
+ _14010_/X sky130_fd_sc_hd__a32o_4
X_11222_ _11424_/A _11222_/B vssd1 vssd1 vccd1 vccd1 _11222_/Y sky130_fd_sc_hd__nor2_1
XFILLER_175_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23208_ _23528_/CLK _23208_/D vssd1 vssd1 vccd1 vccd1 _23208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_342_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_323_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_296_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11153_ _12750_/S vssd1 vssd1 vccd1 vccd1 _13089_/A sky130_fd_sc_hd__clkbuf_2
XTAP_6110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23139_ _23459_/CLK _23139_/D vssd1 vssd1 vccd1 vccd1 _23139_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_296_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15961_ _16109_/A _15961_/B vssd1 vssd1 vccd1 vccd1 _15961_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11084_ _11084_/A vssd1 vssd1 vccd1 vccd1 _14195_/A sky130_fd_sc_hd__clkbuf_4
XTAP_6165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput220 localMemory_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input220/X sky130_fd_sc_hd__buf_6
XTAP_5431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput231 localMemory_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 input231/X sky130_fd_sc_hd__buf_8
XFILLER_310_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17700_ _22730_/Q _17601_/X _17704_/S vssd1 vssd1 vccd1 vccd1 _17701_/A sky130_fd_sc_hd__mux2_1
XTAP_6198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput242 localMemory_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input242/X sky130_fd_sc_hd__buf_4
XFILLER_76_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14912_ _14912_/A vssd1 vssd1 vccd1 vccd1 _14913_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput253 manufacturerID[0] vssd1 vssd1 vccd1 vccd1 input253/X sky130_fd_sc_hd__clkbuf_4
XFILLER_237_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18680_ _23069_/Q _17623_/X _18680_/S vssd1 vssd1 vccd1 vccd1 _18681_/A sky130_fd_sc_hd__mux2_1
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15892_ _15891_/A _15866_/Y _15889_/X _15891_/Y _15818_/A vssd1 vssd1 vccd1 vccd1
+ _15892_/X sky130_fd_sc_hd__o311a_1
Xinput264 partID[0] vssd1 vssd1 vccd1 vccd1 input264/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput275 partID[5] vssd1 vssd1 vccd1 vccd1 input275/X sky130_fd_sc_hd__clkbuf_1
XTAP_5486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17631_ _22704_/Q _17630_/X _17640_/S vssd1 vssd1 vccd1 vccd1 _17632_/A sky130_fd_sc_hd__mux2_1
XFILLER_341_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ _15088_/S _14843_/B vssd1 vssd1 vccd1 vccd1 _14843_/X sky130_fd_sc_hd__and2_1
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17562_ _18788_/A vssd1 vssd1 vccd1 vccd1 _17562_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14774_ _14774_/A vssd1 vssd1 vccd1 vccd1 _14774_/Y sky130_fd_sc_hd__clkinv_2
X_11986_ _11986_/A _11986_/B vssd1 vssd1 vccd1 vccd1 _11986_/X sky130_fd_sc_hd__or2_1
XFILLER_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19301_ _19301_/A vssd1 vssd1 vccd1 vccd1 _23315_/D sky130_fd_sc_hd__clkbuf_1
X_16513_ _15936_/X _22413_/Q _16513_/S vssd1 vssd1 vccd1 vccd1 _16514_/A sky130_fd_sc_hd__mux2_1
X_13725_ _14015_/A _13728_/B _14019_/C vssd1 vssd1 vccd1 vccd1 _13726_/A sky130_fd_sc_hd__and3_4
X_17493_ _17493_/A vssd1 vssd1 vccd1 vccd1 _22654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16444_ _16444_/A vssd1 vssd1 vccd1 vccd1 _22382_/D sky130_fd_sc_hd__clkbuf_1
X_19232_ _19232_/A vssd1 vssd1 vccd1 vccd1 _23289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13656_ _13765_/C _14089_/B vssd1 vssd1 vccd1 vccd1 _13657_/A sky130_fd_sc_hd__or2_1
XFILLER_90_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19163_ _19163_/A vssd1 vssd1 vccd1 vccd1 _19163_/X sky130_fd_sc_hd__clkbuf_2
X_12607_ _12289_/Y _13354_/B _13353_/B _13928_/A vssd1 vssd1 vccd1 vccd1 _15122_/A
+ sky130_fd_sc_hd__o2bb2a_2
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16375_ _16089_/X _22353_/Q _16377_/S vssd1 vssd1 vccd1 vccd1 _16376_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13587_ _13587_/A vssd1 vssd1 vccd1 vccd1 _13588_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_346_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_318_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18114_ _22877_/Q _18051_/A _18113_/X _18105_/X vssd1 vssd1 vccd1 vccd1 _22877_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_307_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15326_ _15324_/X _22271_/Q _15524_/S vssd1 vssd1 vccd1 vccd1 _15327_/A sky130_fd_sc_hd__mux2_1
X_19094_ _23237_/Q _18769_/X _19102_/S vssd1 vssd1 vccd1 vccd1 _19095_/A sky130_fd_sc_hd__mux2_1
X_12538_ _12538_/A _12538_/B vssd1 vssd1 vccd1 vccd1 _12538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_319_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_293_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18045_ _18105_/A vssd1 vssd1 vccd1 vccd1 _18045_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_334_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_333_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_318_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15257_ _13379_/B _15867_/S _15256_/X _20138_/B vssd1 vssd1 vccd1 vccd1 _15257_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12469_ _23887_/Q _13472_/A _12344_/X vssd1 vssd1 vccd1 vccd1 _12469_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_333_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_333_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14208_ _14820_/A _21193_/A _19922_/D _13763_/A vssd1 vssd1 vccd1 vccd1 _21287_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_99_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15188_ _15484_/B vssd1 vssd1 vccd1 vccd1 _15432_/B sky130_fd_sc_hd__buf_2
XFILLER_235_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_334_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14139_ _23011_/Q vssd1 vssd1 vccd1 vccd1 _18536_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_301_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19996_ _23611_/Q _19992_/B _19995_/Y vssd1 vssd1 vccd1 vccd1 _23611_/D sky130_fd_sc_hd__o21a_1
XFILLER_298_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_298_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18947_ _19003_/A vssd1 vssd1 vccd1 vccd1 _19016_/S sky130_fd_sc_hd__buf_6
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_301_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18878_ _18878_/A vssd1 vssd1 vccd1 vccd1 _23141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_143_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _22961_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17829_ _22787_/Q _17578_/X _17837_/S vssd1 vssd1 vccd1 vccd1 _17830_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20840_ _20843_/A _20840_/B vssd1 vssd1 vccd1 vccd1 _20841_/A sky130_fd_sc_hd__and2_1
XFILLER_70_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20771_ _20864_/A vssd1 vssd1 vccd1 vccd1 _20810_/A sky130_fd_sc_hd__buf_4
XINSDIODE2_350 _17217_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_361 _23794_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22510_ _23693_/CLK _22510_/D vssd1 vssd1 vccd1 vccd1 _22510_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_211_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_372 _23465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23490_ _23522_/CLK _23490_/D vssd1 vssd1 vccd1 vccd1 _23490_/Q sky130_fd_sc_hd__dfxtp_2
XINSDIODE2_383 _22491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_394 _14090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22441_ _23480_/CLK _22441_/D vssd1 vssd1 vccd1 vccd1 _22441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_349_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22372_ _23572_/CLK _22372_/D vssd1 vssd1 vccd1 vccd1 _22372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21323_ _21575_/A vssd1 vssd1 vccd1 vccd1 _21712_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_191_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_352_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21254_ _11483_/X _15717_/X _21257_/S vssd1 vssd1 vccd1 vccd1 _21255_/B sky130_fd_sc_hd__mux2_1
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_305_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_333_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20205_ _20205_/A _20532_/D vssd1 vssd1 vccd1 vccd1 _20262_/A sky130_fd_sc_hd__nor2_1
XFILLER_289_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21185_ _21185_/A vssd1 vssd1 vccd1 vccd1 _21281_/A sky130_fd_sc_hd__buf_2
XFILLER_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20136_ _23652_/Q _23651_/Q _20136_/C vssd1 vssd1 vccd1 vccd1 _20137_/C sky130_fd_sc_hd__and3_1
XFILLER_278_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_10 _17303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20067_ _20067_/A vssd1 vssd1 vccd1 vccd1 _21122_/A sky130_fd_sc_hd__buf_6
XFILLER_292_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_21 _22254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_32 _18647_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_43 _21165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_54 _20711_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_65 _21607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_76 _14815_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_87 _14179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_98 _12110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11840_ _11840_/A vssd1 vssd1 vccd1 vccd1 _11840_/X sky130_fd_sc_hd__buf_6
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23826_ _23877_/CLK _23826_/D vssd1 vssd1 vccd1 vccd1 _23826_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _22367_/Q _22399_/Q _22688_/Q _23055_/Q _12070_/S _11613_/A vssd1 vssd1 vccd1
+ vccd1 _11772_/B sky130_fd_sc_hd__mux4_1
X_23757_ _23824_/CLK _23757_/D vssd1 vssd1 vccd1 vccd1 _23757_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20969_ _20969_/A vssd1 vssd1 vccd1 vccd1 _20969_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _13510_/A _13510_/B vssd1 vssd1 vccd1 vccd1 _13511_/B sky130_fd_sc_hd__nand2_1
XFILLER_213_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22708_ _23491_/CLK _22708_/D vssd1 vssd1 vccd1 vccd1 _22708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14490_ _15066_/B _20409_/A vssd1 vssd1 vccd1 vccd1 _14491_/A sky130_fd_sc_hd__or2_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23688_ _23696_/CLK _23688_/D vssd1 vssd1 vccd1 vccd1 _23688_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13441_ _23890_/Q _23889_/Q _23887_/Q vssd1 vssd1 vccd1 vccd1 _13442_/C sky130_fd_sc_hd__or3_1
X_22639_ _23549_/CLK _22639_/D vssd1 vssd1 vccd1 vccd1 _22639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16160_ _18868_/A vssd1 vssd1 vccd1 vccd1 _19261_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_355_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13372_ _13375_/A _13372_/B vssd1 vssd1 vccd1 vccd1 _13372_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15111_ _14074_/D _14246_/B _15110_/X _13688_/A _22502_/Q vssd1 vssd1 vccd1 vccd1
+ _15111_/X sky130_fd_sc_hd__o32a_1
XFILLER_166_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12323_ _11819_/X _12316_/X _12318_/X _12322_/X vssd1 vssd1 vccd1 vccd1 _12323_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_316_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16091_ _16091_/A vssd1 vssd1 vccd1 vccd1 _22289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15042_ _14987_/X _14530_/X _15039_/X _21474_/A _15041_/X vssd1 vssd1 vccd1 vccd1
+ _18788_/A sky130_fd_sc_hd__a32o_4
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12254_ _12291_/A _12253_/X _11713_/A vssd1 vssd1 vccd1 vccd1 _12254_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_331_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11205_ _11205_/A vssd1 vssd1 vccd1 vccd1 _13032_/S sky130_fd_sc_hd__buf_6
XFILLER_269_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19850_ _16214_/X _23559_/Q _19854_/S vssd1 vssd1 vccd1 vccd1 _19851_/A sky130_fd_sc_hd__mux2_1
X_12185_ _12196_/A _12184_/X _11844_/A vssd1 vssd1 vccd1 vccd1 _12185_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_295_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_312_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_311_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_312_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18801_ _18801_/A vssd1 vssd1 vccd1 vccd1 _18801_/X sky130_fd_sc_hd__clkbuf_2
X_11136_ _23901_/Q vssd1 vssd1 vccd1 vccd1 _12534_/A sky130_fd_sc_hd__clkbuf_4
X_19781_ _19781_/A vssd1 vssd1 vccd1 vccd1 _23528_/D sky130_fd_sc_hd__clkbuf_1
X_16993_ _11069_/C _16990_/X _17009_/S vssd1 vssd1 vccd1 vccd1 _16993_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18732_ _18754_/A vssd1 vssd1 vccd1 vccd1 _18741_/S sky130_fd_sc_hd__buf_6
XFILLER_249_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15944_ _13188_/A _15583_/X _15196_/X _13543_/A vssd1 vssd1 vccd1 vccd1 _15944_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_11067_ _11069_/C _11069_/D vssd1 vssd1 vccd1 vccd1 _14814_/C sky130_fd_sc_hd__and2_4
XTAP_5261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18663_ _23061_/Q _17598_/X _18669_/S vssd1 vssd1 vccd1 vccd1 _18664_/A sky130_fd_sc_hd__mux2_1
X_15875_ _22969_/Q _16070_/A vssd1 vssd1 vccd1 vccd1 _15875_/X sky130_fd_sc_hd__or2_1
XTAP_5294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17614_ _18840_/A vssd1 vssd1 vccd1 vccd1 _17614_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_224_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14826_ _22506_/Q _14219_/X _13887_/A _14825_/X vssd1 vssd1 vccd1 vccd1 _15331_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18594_ _18594_/A vssd1 vssd1 vccd1 vccd1 _23030_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ _19091_/A _18625_/B vssd1 vssd1 vccd1 vccd1 _17627_/A sky130_fd_sc_hd__nor2_8
XFILLER_189_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14757_ _14757_/A _15256_/B vssd1 vssd1 vccd1 vccd1 _14757_/X sky130_fd_sc_hd__or2_1
X_11969_ _12130_/A _11969_/B vssd1 vssd1 vccd1 vccd1 _11969_/Y sky130_fd_sc_hd__nor2_1
XFILLER_301_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13708_ _13781_/A vssd1 vssd1 vccd1 vccd1 _13709_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17476_ _17476_/A vssd1 vssd1 vccd1 vccd1 _22646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_338_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14688_ _13476_/A _15079_/B _14686_/Y _14687_/X vssd1 vssd1 vccd1 vccd1 _14688_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19215_ _19213_/X _23284_/Q _19227_/S vssd1 vssd1 vccd1 vccd1 _19216_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16427_ _15710_/X _22375_/Q _16429_/S vssd1 vssd1 vccd1 vccd1 _16428_/A sky130_fd_sc_hd__mux2_1
X_13639_ _14220_/A _14224_/A _13639_/C vssd1 vssd1 vccd1 vccd1 _13640_/A sky130_fd_sc_hd__nor3_4
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19146_ _23261_/Q _18849_/X _19146_/S vssd1 vssd1 vccd1 vccd1 _19147_/A sky130_fd_sc_hd__mux2_1
X_16358_ _15785_/X _22345_/Q _16366_/S vssd1 vssd1 vccd1 vccd1 _16359_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_347_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_346_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_334_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15309_ _22956_/Q _15308_/X _16028_/A vssd1 vssd1 vccd1 vccd1 _15309_/X sky130_fd_sc_hd__mux2_1
X_16289_ _22318_/Q _16287_/X _16301_/S vssd1 vssd1 vccd1 vccd1 _16290_/A sky130_fd_sc_hd__mux2_1
X_19077_ _19077_/A vssd1 vssd1 vccd1 vccd1 _23230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18028_ hold2/A _18017_/X _18020_/X _22980_/Q _18023_/X vssd1 vssd1 vccd1 vccd1 _18028_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_160_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19979_ _20008_/A _19979_/B _20005_/C vssd1 vssd1 vccd1 vccd1 _23606_/D sky130_fd_sc_hd__nor3_1
XFILLER_262_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22990_ _23009_/CLK _22990_/D vssd1 vssd1 vccd1 vccd1 _22990_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_262_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21941_ _23801_/Q _21683_/X _21940_/Y _21346_/X vssd1 vssd1 vccd1 vccd1 _21942_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21872_ _21869_/X _21871_/Y _21847_/A vssd1 vssd1 vccd1 vccd1 _21872_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23611_ _23643_/CLK _23611_/D vssd1 vssd1 vccd1 vccd1 _23611_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_231_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20823_ _20823_/A vssd1 vssd1 vccd1 vccd1 _23761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23542_ _23542_/CLK _23542_/D vssd1 vssd1 vccd1 vccd1 _23542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20754_ _20754_/A _20759_/B vssd1 vssd1 vccd1 vccd1 _20757_/B sky130_fd_sc_hd__and2_1
XINSDIODE2_180 _13720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_287_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_191 _13939_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23473_ _23504_/CLK _23473_/D vssd1 vssd1 vccd1 vccd1 _23473_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_338_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20685_ _20895_/A vssd1 vssd1 vccd1 vccd1 _20744_/B sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_40_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _22789_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_211_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22424_ _23555_/CLK _22424_/D vssd1 vssd1 vccd1 vccd1 _22424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22355_ _23491_/CLK _22355_/D vssd1 vssd1 vccd1 vccd1 _22355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_305_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_353_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21306_ _21379_/A vssd1 vssd1 vccd1 vccd1 _21663_/A sky130_fd_sc_hd__clkbuf_2
X_22286_ _23582_/CLK _22286_/D vssd1 vssd1 vccd1 vccd1 _22286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_317_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_306_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21237_ _15081_/A _21229_/X _21235_/Y _21236_/X vssd1 vssd1 vccd1 vccd1 _23891_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_277_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21168_ _21168_/A vssd1 vssd1 vccd1 vccd1 _21168_/X sky130_fd_sc_hd__buf_2
XFILLER_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20119_ _20119_/A _20126_/D vssd1 vssd1 vccd1 vccd1 _20122_/B sky130_fd_sc_hd__and2_1
X_21099_ _23847_/Q _21096_/X _21098_/X _20547_/A vssd1 vssd1 vccd1 vccd1 _21100_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_13990_ _13990_/A _14087_/A vssd1 vssd1 vccd1 vccd1 _13990_/Y sky130_fd_sc_hd__nor2_8
XFILLER_77_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12941_ _13455_/A _12667_/X _11403_/A _12940_/Y vssd1 vssd1 vccd1 vccd1 _13022_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15660_ _21856_/A _15701_/C vssd1 vssd1 vccd1 vccd1 _15661_/B sky130_fd_sc_hd__xnor2_4
XFILLER_45_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _22314_/Q _23450_/Q _12977_/S vssd1 vssd1 vccd1 vccd1 _12872_/X sky130_fd_sc_hd__mux2_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _14922_/A vssd1 vssd1 vccd1 vccd1 _15222_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _23407_/Q _23023_/Q _23375_/Q _23343_/Q _11814_/X _11800_/A vssd1 vssd1 vccd1
+ vccd1 _11824_/B sky130_fd_sc_hd__mux4_1
X_23809_ _23810_/CLK _23809_/D vssd1 vssd1 vccd1 vccd1 _23809_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _23605_/Q _15589_/X _15590_/X _23637_/Q vssd1 vssd1 vccd1 vccd1 _15591_/X
+ sky130_fd_sc_hd__o22a_2
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _17330_/A vssd1 vssd1 vccd1 vccd1 _22587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _16936_/B vssd1 vssd1 vccd1 vccd1 _21294_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_199_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _11754_/A vssd1 vssd1 vccd1 vccd1 _11755_/A sky130_fd_sc_hd__buf_2
XFILLER_159_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_348_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _22116_/A _17260_/X _17292_/S vssd1 vssd1 vccd1 vccd1 _17261_/X sky130_fd_sc_hd__mux2_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14473_ _14473_/A _20989_/A vssd1 vssd1 vccd1 vccd1 _14474_/A sky130_fd_sc_hd__nor2_1
XFILLER_14_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11685_ _12156_/A _11685_/B _11685_/C vssd1 vssd1 vccd1 vccd1 _20303_/A sky130_fd_sc_hd__nand3_4
XFILLER_230_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_347_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19000_ _19000_/A vssd1 vssd1 vccd1 vccd1 _23196_/D sky130_fd_sc_hd__clkbuf_1
X_16212_ _22294_/Q _16211_/X _16221_/S vssd1 vssd1 vccd1 vccd1 _16213_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13424_ _14760_/A _14251_/A _14388_/C vssd1 vssd1 vccd1 vccd1 _13428_/B sky130_fd_sc_hd__mux2_1
XFILLER_347_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17192_ _23480_/Q _17113_/X _17114_/X _17181_/X _15738_/Y vssd1 vssd1 vccd1 vccd1
+ _17192_/X sky130_fd_sc_hd__a32o_1
XFILLER_316_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_329_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_356_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_328_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16143_ _15440_/X _16136_/X _16142_/X _14497_/A vssd1 vssd1 vccd1 vccd1 _16143_/X
+ sky130_fd_sc_hd__o22a_1
X_13355_ _13355_/A vssd1 vssd1 vccd1 vccd1 _13906_/A sky130_fd_sc_hd__inv_2
XFILLER_316_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12306_ _22266_/Q _23082_/Q _23498_/Q _22427_/Q _11113_/A _11565_/A vssd1 vssd1 vccd1
+ vccd1 _12307_/B sky130_fd_sc_hd__mux4_1
X_16074_ _14215_/A _21276_/A _16073_/X _11099_/A vssd1 vssd1 vccd1 vccd1 _16074_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_316_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13286_ _23233_/Q _23201_/Q _23169_/Q _23137_/Q _11461_/A _11365_/X vssd1 vssd1 vccd1
+ vccd1 _13287_/B sky130_fd_sc_hd__mux4_1
XFILLER_288_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19902_ _19902_/A vssd1 vssd1 vccd1 vccd1 _23582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15025_ _15010_/Y _15024_/X _14520_/A vssd1 vssd1 vccd1 vccd1 _15025_/Y sky130_fd_sc_hd__o21ai_2
X_12237_ _13510_/A vssd1 vssd1 vccd1 vccd1 _13928_/A sky130_fd_sc_hd__buf_2
XFILLER_297_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_297_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_300_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19833_ _23552_/Q _19252_/A _19837_/S vssd1 vssd1 vccd1 vccd1 _19834_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_296_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12168_ _12168_/A _12168_/B vssd1 vssd1 vccd1 vccd1 _12168_/Y sky130_fd_sc_hd__nand2_1
XFILLER_311_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_300_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11119_ _11595_/A _20533_/B vssd1 vssd1 vccd1 vccd1 _12468_/B sky130_fd_sc_hd__nor2_8
XFILLER_300_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19764_ _19764_/A vssd1 vssd1 vccd1 vccd1 _23521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16976_ _23944_/Q _17648_/B _17022_/A vssd1 vssd1 vccd1 vccd1 _16976_/X sky130_fd_sc_hd__a21o_1
X_12099_ _11631_/A _12091_/X _12093_/X _12098_/X _11657_/A vssd1 vssd1 vccd1 vccd1
+ _12109_/B sky130_fd_sc_hd__a311o_1
XFILLER_232_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18715_ _16838_/X _23084_/Q _18719_/S vssd1 vssd1 vccd1 vccd1 _18716_/A sky130_fd_sc_hd__mux2_1
Xinput6 coreIndex[5] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15927_ _15752_/X _15926_/X _15480_/A vssd1 vssd1 vccd1 vccd1 _15927_/X sky130_fd_sc_hd__o21a_1
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19695_ _19261_/X _23491_/Q _19697_/S vssd1 vssd1 vccd1 vccd1 _19696_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18646_ _18646_/A vssd1 vssd1 vccd1 vccd1 _23053_/D sky130_fd_sc_hd__clkbuf_1
X_15858_ _23000_/Q _15931_/A _15932_/A input229/X vssd1 vssd1 vccd1 vccd1 _22003_/A
+ sky130_fd_sc_hd__a22o_4
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14809_ _14210_/X _21351_/B _14805_/X _14808_/X vssd1 vssd1 vccd1 vccd1 _18779_/A
+ sky130_fd_sc_hd__a2bb2o_4
X_18577_ _18623_/S vssd1 vssd1 vccd1 vccd1 _18586_/S sky130_fd_sc_hd__buf_4
X_15789_ _22999_/Q _15931_/A _15932_/A input228/X vssd1 vssd1 vccd1 vccd1 _21979_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_33_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17528_ _17528_/A vssd1 vssd1 vccd1 vccd1 _22670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_299_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17459_ _22640_/Q _16291_/X _17465_/S vssd1 vssd1 vccd1 vccd1 _17460_/A sky130_fd_sc_hd__mux2_1
XFILLER_339_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20470_ _20470_/A vssd1 vssd1 vccd1 vccd1 _20487_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_319_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19129_ _23253_/Q _18824_/X _19135_/S vssd1 vssd1 vccd1 vccd1 _19130_/A sky130_fd_sc_hd__mux2_1
XFILLER_307_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22140_ _22140_/A _22140_/B vssd1 vssd1 vccd1 vccd1 _22142_/B sky130_fd_sc_hd__nor2_1
XFILLER_195_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput310 _13964_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[15] sky130_fd_sc_hd__buf_2
XFILLER_133_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput321 _13984_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[26] sky130_fd_sc_hd__buf_2
XFILLER_156_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_322_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput332 _13697_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[0] sky130_fd_sc_hd__buf_2
XFILLER_350_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput343 _13701_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[1] sky130_fd_sc_hd__buf_2
X_22071_ _22071_/A _22071_/B vssd1 vssd1 vccd1 vccd1 _23935_/D sky130_fd_sc_hd__nor2_1
XTAP_6709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput354 _13713_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[2] sky130_fd_sc_hd__buf_2
Xoutput365 _13883_/Y vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[1] sky130_fd_sc_hd__buf_2
XFILLER_99_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_288_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput376 _14030_/X vssd1 vssd1 vccd1 vccd1 din0[11] sky130_fd_sc_hd__buf_2
Xoutput387 _14050_/X vssd1 vssd1 vccd1 vccd1 din0[21] sky130_fd_sc_hd__buf_2
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21022_ _23824_/Q _21028_/B vssd1 vssd1 vccd1 vccd1 _21022_/X sky130_fd_sc_hd__or2_1
XFILLER_302_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput398 _14070_/X vssd1 vssd1 vccd1 vccd1 din0[31] sky130_fd_sc_hd__buf_2
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22973_ _22974_/CLK _22973_/D vssd1 vssd1 vccd1 vccd1 _22973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21924_ _21916_/A _21612_/X _21923_/X _21896_/X vssd1 vssd1 vccd1 vccd1 _23930_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21855_ _23798_/Q _21381_/X _21854_/X _21813_/A vssd1 vssd1 vccd1 vccd1 _21855_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_270_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20806_ _20806_/A _20806_/B vssd1 vssd1 vccd1 vccd1 _20807_/A sky130_fd_sc_hd__and2_1
XFILLER_212_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21786_ _21786_/A _21786_/B vssd1 vssd1 vccd1 vccd1 _21787_/B sky130_fd_sc_hd__nor2_1
XFILLER_358_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23525_ _23525_/CLK _23525_/D vssd1 vssd1 vccd1 vccd1 _23525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20737_ _20763_/A vssd1 vssd1 vccd1 vccd1 _20737_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_358_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_345_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_329_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_345_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23456_ _23456_/CLK _23456_/D vssd1 vssd1 vccd1 vccd1 _23456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11470_ _23331_/Q _23299_/Q _23267_/Q _23555_/Q _21771_/A _15616_/A vssd1 vssd1 vccd1
+ vccd1 _11471_/B sky130_fd_sc_hd__mux4_1
X_20668_ _20730_/A vssd1 vssd1 vccd1 vccd1 _20695_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22407_ _23544_/CLK _22407_/D vssd1 vssd1 vccd1 vccd1 _22407_/Q sky130_fd_sc_hd__dfxtp_1
X_23387_ _23545_/CLK _23387_/D vssd1 vssd1 vccd1 vccd1 _23387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_353_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20599_ _13440_/B _20564_/X _20598_/X vssd1 vssd1 vccd1 vccd1 _20599_/X sky130_fd_sc_hd__a21o_1
XFILLER_326_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13140_ _13491_/A _15996_/A vssd1 vssd1 vccd1 vccd1 _13402_/A sky130_fd_sc_hd__or2_2
XFILLER_354_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_341_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22338_ _23538_/CLK _22338_/D vssd1 vssd1 vccd1 vccd1 _22338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_352_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_313_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13071_ _13121_/A _13070_/X _12745_/X vssd1 vssd1 vccd1 vccd1 _13071_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_340_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22269_ _23565_/CLK _22269_/D vssd1 vssd1 vccd1 vccd1 _22269_/Q sky130_fd_sc_hd__dfxtp_1
X_12022_ _12852_/A _12021_/X _11681_/X vssd1 vssd1 vccd1 vccd1 _12022_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_250_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_294_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16830_ _16830_/A vssd1 vssd1 vccd1 vccd1 _22525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_265_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16761_ _16779_/A vssd1 vssd1 vccd1 vccd1 _16777_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13973_ _13973_/A vssd1 vssd1 vccd1 vccd1 _13973_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18500_ _22995_/Q _18505_/B vssd1 vssd1 vccd1 vccd1 _18500_/Y sky130_fd_sc_hd__nand2_1
XFILLER_219_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15712_ _15712_/A vssd1 vssd1 vccd1 vccd1 _22279_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_274_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12924_ _13096_/A _12921_/X _12923_/X vssd1 vssd1 vccd1 vccd1 _12924_/Y sky130_fd_sc_hd__a21oi_1
X_19480_ _19480_/A vssd1 vssd1 vccd1 vccd1 _23395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16692_ _16784_/A vssd1 vssd1 vccd1 vccd1 _16730_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_47_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18431_ _22971_/Q _18429_/B _18430_/Y vssd1 vssd1 vccd1 vccd1 _22971_/D sky130_fd_sc_hd__o21a_1
X_12855_ _23228_/Q _23196_/Q _23164_/Q _23132_/Q _12843_/X _12844_/X vssd1 vssd1 vccd1
+ vccd1 _12856_/B sky130_fd_sc_hd__mux4_2
X_15643_ _22931_/Q _14752_/X _14753_/X _15644_/A vssd1 vssd1 vccd1 vccd1 _15643_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _12097_/A _11806_/B vssd1 vssd1 vccd1 vccd1 _11806_/X sky130_fd_sc_hd__or2_1
XFILLER_349_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18362_ _14729_/X _18366_/C _18337_/X vssd1 vssd1 vccd1 vccd1 _18362_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15574_ _15574_/A vssd1 vssd1 vccd1 vccd1 _15574_/X sky130_fd_sc_hd__clkbuf_2
X_12786_ _12906_/A _12785_/X _12721_/A vssd1 vssd1 vccd1 vccd1 _12786_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _22583_/Q _17091_/A _17028_/A _17312_/X vssd1 vssd1 vccd1 vccd1 _22583_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_30_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _15478_/A vssd1 vssd1 vccd1 vccd1 _14529_/A sky130_fd_sc_hd__buf_2
X_11737_ _11742_/A vssd1 vssd1 vccd1 vccd1 _12014_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_187_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18293_ _18296_/A _18296_/C _18292_/X vssd1 vssd1 vccd1 vccd1 _18293_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_358_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_308_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14456_ _23589_/Q _14450_/X _14455_/X _23621_/Q vssd1 vssd1 vccd1 vccd1 _14456_/X
+ sky130_fd_sc_hd__o22a_2
X_17244_ _22812_/Q _17244_/B _17244_/C vssd1 vssd1 vccd1 vccd1 _17245_/A sky130_fd_sc_hd__and3_1
XFILLER_187_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11668_ _12024_/A vssd1 vssd1 vccd1 vccd1 _12716_/A sky130_fd_sc_hd__buf_4
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13407_ _13399_/A _13399_/B _13242_/X vssd1 vssd1 vccd1 vccd1 _13408_/B sky130_fd_sc_hd__a21oi_1
X_17175_ _17169_/X _17173_/Y _17174_/Y _17024_/X vssd1 vssd1 vccd1 vccd1 _17175_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_344_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14387_ _14264_/X _14367_/X _14382_/X _14384_/X _16186_/A vssd1 vssd1 vccd1 vccd1
+ _14389_/B sky130_fd_sc_hd__o221a_2
XFILLER_127_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_317_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11599_ _11141_/A _11597_/X _11598_/X vssd1 vssd1 vccd1 vccd1 _11599_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_127_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16126_ _16126_/A vssd1 vssd1 vccd1 vccd1 _22290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_344_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13338_ _13646_/A _13392_/A vssd1 vssd1 vccd1 vccd1 _13338_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16057_ _16057_/A _16057_/B vssd1 vssd1 vccd1 vccd1 _16057_/X sky130_fd_sc_hd__or2_1
X_13269_ _23489_/Q _23585_/Q _22549_/Q _22353_/Q _11492_/S _11200_/A vssd1 vssd1 vccd1
+ vccd1 _13269_/X sky130_fd_sc_hd__mux4_1
XFILLER_170_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15008_ _16053_/S vssd1 vssd1 vccd1 vccd1 _15867_/S sky130_fd_sc_hd__buf_4
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_312_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19816_ _19816_/A vssd1 vssd1 vccd1 vccd1 _23544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_296_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19747_ _19747_/A vssd1 vssd1 vccd1 vccd1 _23513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16959_ _16962_/A _21294_/C _16936_/B vssd1 vssd1 vccd1 vccd1 _17248_/A sky130_fd_sc_hd__or3b_4
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19678_ _19236_/X _23483_/Q _19682_/S vssd1 vssd1 vccd1 vccd1 _19679_/A sky130_fd_sc_hd__mux2_1
XFILLER_271_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18629_ _18629_/A vssd1 vssd1 vccd1 vccd1 _23045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21640_ _21640_/A _21640_/B vssd1 vssd1 vccd1 vccd1 _21640_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_162_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21571_ _23919_/Q _21576_/A vssd1 vssd1 vccd1 vccd1 _21572_/B sky130_fd_sc_hd__and2_1
XFILLER_178_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23310_ _23534_/CLK _23310_/D vssd1 vssd1 vccd1 vccd1 _23310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20522_ _23709_/Q _20523_/B _20522_/C vssd1 vssd1 vccd1 vccd1 _20525_/B sky130_fd_sc_hd__and3_1
XFILLER_339_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_327_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23241_ _23529_/CLK _23241_/D vssd1 vssd1 vccd1 vccd1 _23241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_319_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20453_ _21033_/A _20463_/B vssd1 vssd1 vccd1 vccd1 _20453_/Y sky130_fd_sc_hd__nand2_1
XFILLER_307_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23172_ _23578_/CLK _23172_/D vssd1 vssd1 vccd1 vccd1 _23172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_350_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20384_ _20320_/X _20382_/Y _20383_/X _22171_/A _20294_/X vssd1 vssd1 vccd1 vccd1
+ _20749_/A sky130_fd_sc_hd__a32o_4
XFILLER_107_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_7207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_350_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22123_ _22114_/A _21984_/X _22121_/Y _22122_/X vssd1 vssd1 vccd1 vccd1 _23937_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22054_ _23805_/Q _21560_/X _22053_/Y _21613_/X vssd1 vssd1 vccd1 vccd1 _22054_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_82_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21005_ _20585_/A _20988_/X _21004_/X _20997_/X vssd1 vssd1 vccd1 vccd1 _23817_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_287_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22956_ _22956_/CLK _22956_/D vssd1 vssd1 vccd1 vccd1 _22956_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_244_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21907_ _21933_/B _21907_/B vssd1 vssd1 vccd1 vccd1 _21907_/X sky130_fd_sc_hd__xor2_1
XFILLER_83_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22887_ _23552_/CLK _22887_/D vssd1 vssd1 vccd1 vccd1 _22887_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_203_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12640_ _11584_/A _12639_/X _12656_/A vssd1 vssd1 vccd1 vccd1 _12640_/X sky130_fd_sc_hd__a21o_1
XFILLER_102_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21838_ _21838_/A _21838_/B vssd1 vssd1 vccd1 vccd1 _21838_/Y sky130_fd_sc_hd__nand2_1
XPHY_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_358_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_321_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12571_ _12196_/X _12568_/X _12570_/X _11844_/X vssd1 vssd1 vccd1 vccd1 _12571_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21769_ _21307_/X _21753_/X _21760_/Y _21768_/X _21329_/X vssd1 vssd1 vccd1 vccd1
+ _21769_/Y sky130_fd_sc_hd__o2111ai_2
XFILLER_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14310_ _14308_/Y _14309_/X _14310_/S vssd1 vssd1 vccd1 vccd1 _14310_/X sky130_fd_sc_hd__mux2_1
XPHY_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23508_ _23510_/CLK _23508_/D vssd1 vssd1 vccd1 vccd1 _23508_/Q sky130_fd_sc_hd__dfxtp_1
X_11522_ _13229_/A vssd1 vssd1 vccd1 vccd1 _13218_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_196_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15290_ _13383_/X _13948_/Y _15867_/S vssd1 vssd1 vccd1 vccd1 _15290_/X sky130_fd_sc_hd__mux2_1
XFILLER_346_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14241_ _14241_/A _15112_/A vssd1 vssd1 vccd1 vccd1 _15179_/A sky130_fd_sc_hd__nor2_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23439_ _23503_/CLK _23439_/D vssd1 vssd1 vccd1 vccd1 _23439_/Q sky130_fd_sc_hd__dfxtp_1
X_11453_ _14175_/A _16005_/A _11403_/X _11452_/Y vssd1 vssd1 vccd1 vccd1 _13306_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_328_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_314_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14172_ _14132_/A _14172_/B _14172_/C vssd1 vssd1 vccd1 vccd1 _14524_/B sky130_fd_sc_hd__and3b_1
XFILLER_354_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_298_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11384_ _12283_/B vssd1 vssd1 vccd1 vccd1 _12415_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_124_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13123_ _13131_/A _13122_/X _11352_/A vssd1 vssd1 vccd1 vccd1 _13123_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_340_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_313_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18980_ _18980_/A vssd1 vssd1 vccd1 vccd1 _23187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17931_ _22822_/Q _17914_/X _17929_/X _17930_/X vssd1 vssd1 vccd1 vccd1 _22822_/D
+ sky130_fd_sc_hd__o211a_1
X_13054_ _13046_/Y _13049_/Y _13051_/Y _13053_/Y _11247_/A vssd1 vssd1 vccd1 vccd1
+ _13054_/X sky130_fd_sc_hd__o221a_1
XFILLER_112_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12005_ _12171_/A _12170_/A vssd1 vssd1 vccd1 vccd1 _12005_/Y sky130_fd_sc_hd__nand2_1
X_17862_ _22802_/Q _17626_/X _17870_/S vssd1 vssd1 vccd1 vccd1 _17863_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_294_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19601_ _19612_/A vssd1 vssd1 vccd1 vccd1 _19610_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_282_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16813_ _19163_/A vssd1 vssd1 vccd1 vccd1 _16813_/X sky130_fd_sc_hd__buf_2
XFILLER_4_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17793_ _17793_/A vssd1 vssd1 vccd1 vccd1 _22771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_266_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19532_ _19233_/X _23418_/Q _19538_/S vssd1 vssd1 vccd1 vccd1 _19533_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16744_ _22501_/Q _16729_/X _16730_/X input15/X vssd1 vssd1 vccd1 vccd1 _16745_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_219_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13956_ _13956_/A _13967_/B vssd1 vssd1 vccd1 vccd1 _13957_/A sky130_fd_sc_hd__and2_1
XFILLER_185_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19463_ _19463_/A vssd1 vssd1 vccd1 vccd1 _23387_/D sky130_fd_sc_hd__clkbuf_1
X_12907_ _23322_/Q _23290_/Q _23258_/Q _23546_/Q _12792_/X _12793_/X vssd1 vssd1 vccd1
+ vccd1 _12907_/X sky130_fd_sc_hd__mux4_2
XFILLER_290_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13887_ _13887_/A vssd1 vssd1 vccd1 vccd1 _13888_/B sky130_fd_sc_hd__buf_6
X_16675_ _22484_/Q _16303_/X _16677_/S vssd1 vssd1 vccd1 vccd1 _16676_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18414_ _22965_/Q _18412_/B _18413_/Y vssd1 vssd1 vccd1 vccd1 _22965_/D sky130_fd_sc_hd__o21a_1
X_15626_ _15625_/X _22277_/Q _15750_/S vssd1 vssd1 vccd1 vccd1 _15627_/A sky130_fd_sc_hd__mux2_1
X_12838_ _11218_/A _12828_/X _12837_/X _11124_/A vssd1 vssd1 vccd1 vccd1 _12839_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19394_ _23357_/Q _18849_/X _19394_/S vssd1 vssd1 vccd1 vccd1 _19395_/A sky130_fd_sc_hd__mux2_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18345_ _22941_/Q _18343_/B _18344_/Y vssd1 vssd1 vccd1 vccd1 _22941_/D sky130_fd_sc_hd__o21a_1
X_12769_ _12886_/A _12769_/B vssd1 vssd1 vccd1 vccd1 _12769_/Y sky130_fd_sc_hd__nor2_1
X_15557_ _15835_/B _15557_/B vssd1 vssd1 vccd1 vccd1 _15557_/Y sky130_fd_sc_hd__nand2_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_348_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_168_wb_clk_i _23917_/CLK vssd1 vssd1 vccd1 vccd1 _23714_/CLK sky130_fd_sc_hd__clkbuf_16
X_14508_ _14752_/A vssd1 vssd1 vccd1 vccd1 _14509_/A sky130_fd_sc_hd__clkbuf_2
X_18276_ _18315_/A _18276_/B _18276_/C vssd1 vssd1 vccd1 vccd1 _22919_/D sky130_fd_sc_hd__nor3_1
X_15488_ _15488_/A vssd1 vssd1 vccd1 vccd1 _15488_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_336_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17227_ _22575_/Q _17199_/X _17190_/X _17226_/X vssd1 vssd1 vccd1 vccd1 _22575_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_308_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput20 core_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_1
X_14439_ _14588_/A vssd1 vssd1 vccd1 vccd1 _16168_/B sky130_fd_sc_hd__clkbuf_2
Xinput31 core_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
XFILLER_317_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 core_wb_error_i vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 dout0[19] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_2
XFILLER_317_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput64 dout0[29] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_2
XFILLER_7_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17158_ _14167_/X _15606_/Y _17009_/S _17157_/Y vssd1 vssd1 vccd1 vccd1 _17158_/X
+ sky130_fd_sc_hd__o211a_1
Xinput75 dout0[39] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__clkbuf_1
XFILLER_289_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput86 dout0[49] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_318_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput97 dout0[59] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16109_ _16109_/A _16109_/B vssd1 vssd1 vccd1 vccd1 _16109_/Y sky130_fd_sc_hd__nand2_1
X_17089_ _17070_/X _17084_/X _17088_/X _17057_/X vssd1 vssd1 vccd1 vccd1 _17089_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_171_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_331_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_297_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22810_ _22968_/CLK _22810_/D vssd1 vssd1 vccd1 vccd1 _22810_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23790_ _23862_/CLK _23790_/D vssd1 vssd1 vccd1 vccd1 _23790_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_203_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22741_ _23073_/CLK _22741_/D vssd1 vssd1 vccd1 vccd1 _22741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_344_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22672_ _23583_/CLK _22672_/D vssd1 vssd1 vccd1 vccd1 _22672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_279_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21623_ _21624_/A _21624_/C _21624_/B vssd1 vssd1 vccd1 vccd1 _21625_/A sky130_fd_sc_hd__o21ai_1
XFILLER_178_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21554_ _20234_/A _21841_/A _15234_/B _21842_/A vssd1 vssd1 vccd1 vccd1 _21554_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_328_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20505_ _23713_/Q _20524_/B _20505_/C vssd1 vssd1 vccd1 vccd1 _20509_/A sky130_fd_sc_hd__and3_1
XFILLER_308_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21485_ _21485_/A _21485_/B vssd1 vssd1 vccd1 vccd1 _21543_/C sky130_fd_sc_hd__nand2_1
XFILLER_354_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_308_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23224_ _23420_/CLK _23224_/D vssd1 vssd1 vccd1 vccd1 _23224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_314_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20436_ _23693_/Q _20448_/B vssd1 vssd1 vccd1 vccd1 _20436_/X sky130_fd_sc_hd__or2_1
XFILLER_165_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23155_ _23507_/CLK _23155_/D vssd1 vssd1 vccd1 vccd1 _23155_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_7026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20367_ _20333_/X _20731_/A _20366_/X _20360_/X vssd1 vssd1 vccd1 vccd1 _23678_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_7037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22106_ _22082_/A _22082_/B _22081_/A vssd1 vssd1 vccd1 vccd1 _22110_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_7059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23086_ _23502_/CLK _23086_/D vssd1 vssd1 vccd1 vccd1 _23086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20298_ _20227_/X _20296_/Y _20187_/X vssd1 vssd1 vccd1 vccd1 _20298_/X sky130_fd_sc_hd__o21a_1
XFILLER_322_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_314_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22037_ _21989_/A _22037_/B vssd1 vssd1 vccd1 vccd1 _22038_/C sky130_fd_sc_hd__and2b_1
XTAP_6369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ _13821_/A _13810_/B vssd1 vssd1 vccd1 vccd1 _13857_/B sky130_fd_sc_hd__or2_1
XFILLER_263_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14790_ _14780_/X _14789_/X _15341_/S vssd1 vssd1 vccd1 vccd1 _14790_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13741_ _13786_/A _13741_/B vssd1 vssd1 vccd1 vccd1 _13742_/A sky130_fd_sc_hd__and2_4
X_22939_ _23649_/CLK _22939_/D vssd1 vssd1 vccd1 vccd1 _22939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_290_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13672_ _13993_/A _13657_/A _13671_/Y vssd1 vssd1 vccd1 vccd1 _14080_/A sky130_fd_sc_hd__o21a_1
X_16460_ _16528_/S vssd1 vssd1 vccd1 vccd1 _16469_/S sky130_fd_sc_hd__buf_8
XFILLER_71_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12623_ _12900_/A _12622_/X _11285_/A vssd1 vssd1 vccd1 vccd1 _12623_/Y sky130_fd_sc_hd__o21ai_1
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15411_ _15379_/Y _15410_/X _20493_/B vssd1 vssd1 vccd1 vccd1 _15412_/B sky130_fd_sc_hd__mux2_1
X_16391_ _16391_/A vssd1 vssd1 vccd1 vccd1 _22358_/D sky130_fd_sc_hd__clkbuf_1
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_346_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18130_ _18116_/A _14107_/X _22881_/Q vssd1 vssd1 vccd1 vccd1 _18130_/X sky130_fd_sc_hd__a21o_1
XPHY_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15342_ _13621_/A _14676_/B _14942_/A _13646_/A _13439_/A vssd1 vssd1 vccd1 vccd1
+ _15342_/X sky130_fd_sc_hd__o221a_1
XPHY_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12554_ _22458_/Q _22618_/Q _12554_/S vssd1 vssd1 vccd1 vccd1 _12554_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_339_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_346_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11505_ _22290_/Q _23106_/Q _23522_/Q _22451_/Q _11432_/X _11435_/X vssd1 vssd1 vccd1
+ vccd1 _11506_/B sky130_fd_sc_hd__mux4_2
XFILLER_12_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18061_ hold8/A _18051_/X _18059_/X _18060_/X vssd1 vssd1 vccd1 vccd1 _22858_/D sky130_fd_sc_hd__o211a_1
X_15273_ _14215_/X _21227_/A _15272_/X _14882_/X vssd1 vssd1 vccd1 vccd1 _15273_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_12485_ _12485_/A _12485_/B vssd1 vssd1 vccd1 vccd1 _12485_/X sky130_fd_sc_hd__or2_1
XFILLER_156_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14224_ _14224_/A _14224_/B vssd1 vssd1 vccd1 vccd1 _15110_/S sky130_fd_sc_hd__or2_4
X_17012_ _17237_/A vssd1 vssd1 vccd1 vccd1 _17012_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11436_ _22807_/Q _22775_/Q _22676_/Q _22743_/Q _11432_/X _11435_/X vssd1 vssd1 vccd1
+ vccd1 _11437_/B sky130_fd_sc_hd__mux4_1
XFILLER_298_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14155_ _22910_/Q _14159_/A _14151_/X _22603_/Q vssd1 vssd1 vccd1 vccd1 _16941_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_125_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11367_ _13278_/A _11367_/B vssd1 vssd1 vccd1 vccd1 _11367_/X sky130_fd_sc_hd__or2_1
XFILLER_98_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ _22287_/Q _23103_/Q _23519_/Q _22448_/Q _13190_/S _11207_/A vssd1 vssd1 vccd1
+ vccd1 _13107_/B sky130_fd_sc_hd__mux4_2
XFILLER_286_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14086_ _22590_/Q _14081_/X _14085_/Y _14083_/X vssd1 vssd1 vccd1 vccd1 _14086_/X
+ sky130_fd_sc_hd__a22o_4
X_18963_ _18963_/A vssd1 vssd1 vccd1 vccd1 _23179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_301_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11298_ _13225_/A vssd1 vssd1 vccd1 vccd1 _13121_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_286_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17914_ _17932_/A vssd1 vssd1 vccd1 vccd1 _17914_/X sky130_fd_sc_hd__clkbuf_2
X_13037_ _13037_/A vssd1 vssd1 vccd1 vccd1 _13037_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_279_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18894_ _23149_/Q _18798_/X _18896_/S vssd1 vssd1 vccd1 vccd1 _18895_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17845_ _17845_/A vssd1 vssd1 vccd1 vccd1 _22794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_282_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17776_ _22764_/Q _17607_/X _17776_/S vssd1 vssd1 vccd1 vccd1 _17777_/A sky130_fd_sc_hd__mux2_1
X_14988_ _22919_/Q _14988_/B vssd1 vssd1 vccd1 vccd1 _14988_/X sky130_fd_sc_hd__and2_1
XFILLER_240_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19515_ _19515_/A vssd1 vssd1 vccd1 vccd1 _23410_/D sky130_fd_sc_hd__clkbuf_1
X_16727_ _16741_/A _16727_/B vssd1 vssd1 vccd1 vccd1 _16728_/A sky130_fd_sc_hd__or2_1
XFILLER_241_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13939_ _13951_/A _13939_/B vssd1 vssd1 vccd1 vccd1 _13939_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_510 _15914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_521 _14045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19446_ _19468_/A vssd1 vssd1 vccd1 vccd1 _19455_/S sky130_fd_sc_hd__clkbuf_4
XINSDIODE2_532 _14127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16658_ _22476_/Q _16278_/X _16662_/S vssd1 vssd1 vccd1 vccd1 _16659_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_543 _14076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_554 _15914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_565 _22601_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15609_ _23927_/Q vssd1 vssd1 vccd1 vccd1 _21826_/A sky130_fd_sc_hd__clkbuf_2
X_19377_ _23349_/Q _18824_/X _19383_/S vssd1 vssd1 vccd1 vccd1 _19378_/A sky130_fd_sc_hd__mux2_1
XFILLER_304_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16589_ _16589_/A vssd1 vssd1 vccd1 vccd1 _22445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_349_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18328_ _22935_/Q _18326_/B _18327_/Y vssd1 vssd1 vccd1 vccd1 _22935_/D sky130_fd_sc_hd__o21a_1
XFILLER_176_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_336_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18259_ _18277_/A vssd1 vssd1 vccd1 vccd1 _20067_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_200_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_318_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21270_ _21281_/A vssd1 vssd1 vccd1 vccd1 _21270_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_351_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20221_ _20275_/A _20217_/Y _20320_/A vssd1 vssd1 vccd1 vccd1 _20221_/X sky130_fd_sc_hd__o21a_1
XFILLER_305_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_304_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_332_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20152_ _17149_/A _20499_/B _20197_/S vssd1 vssd1 vccd1 vccd1 _20152_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_65_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23511_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_304_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_311_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20083_ _20090_/C _20090_/D _20082_/X vssd1 vssd1 vccd1 vccd1 _23635_/D sky130_fd_sc_hd__o21ba_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23911_ _23911_/CLK _23911_/D vssd1 vssd1 vccd1 vccd1 _23911_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23842_ _23876_/CLK _23842_/D vssd1 vssd1 vccd1 vccd1 _23842_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_245_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23773_ _23841_/CLK _23773_/D vssd1 vssd1 vccd1 vccd1 _23773_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20985_ _23812_/Q _20925_/A _20984_/X _20978_/X vssd1 vssd1 vccd1 vccd1 _23812_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22724_ _23058_/CLK _22724_/D vssd1 vssd1 vccd1 vccd1 _22724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_300_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_300_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22655_ _23566_/CLK _22655_/D vssd1 vssd1 vccd1 vccd1 _22655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_328_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21606_ _21559_/A _21559_/B _21605_/X vssd1 vssd1 vccd1 vccd1 _21614_/B sky130_fd_sc_hd__o21ba_1
XFILLER_279_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22586_ _22968_/CLK _22586_/D vssd1 vssd1 vccd1 vccd1 _22586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21537_ _21530_/Y _21535_/X _22214_/S vssd1 vssd1 vccd1 vccd1 _21537_/X sky130_fd_sc_hd__mux2_2
XFILLER_279_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_343_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12270_ _22267_/Q _23083_/Q _23499_/Q _22428_/Q _11920_/X _12269_/X vssd1 vssd1 vccd1
+ vccd1 _12270_/X sky130_fd_sc_hd__mux4_2
X_21468_ _23916_/Q _21474_/A vssd1 vssd1 vccd1 vccd1 _21468_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11221_ _23332_/Q _23300_/Q _23268_/Q _23556_/Q _13434_/A _11170_/X vssd1 vssd1 vccd1
+ vccd1 _11222_/B sky130_fd_sc_hd__mux4_1
XFILLER_181_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23207_ _23367_/CLK _23207_/D vssd1 vssd1 vccd1 vccd1 _23207_/Q sky130_fd_sc_hd__dfxtp_1
X_20419_ _23687_/Q _20429_/B vssd1 vssd1 vccd1 vccd1 _20419_/X sky130_fd_sc_hd__or2_1
XFILLER_175_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21399_ _21400_/A _21406_/A vssd1 vssd1 vccd1 vccd1 _21401_/A sky130_fd_sc_hd__nor2_1
XFILLER_325_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11152_ _12751_/S vssd1 vssd1 vccd1 vccd1 _12750_/S sky130_fd_sc_hd__buf_6
XFILLER_323_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23138_ _23489_/CLK _23138_/D vssd1 vssd1 vccd1 vccd1 _23138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_350_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_296_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23069_ _23073_/CLK _23069_/D vssd1 vssd1 vccd1 vccd1 _23069_/Q sky130_fd_sc_hd__dfxtp_1
X_15960_ _14592_/A _15953_/X _15959_/Y _15652_/X vssd1 vssd1 vccd1 vccd1 _15961_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_11083_ _21335_/A _14187_/A _21335_/C vssd1 vssd1 vccd1 vccd1 _11084_/A sky130_fd_sc_hd__and3_1
XTAP_6166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput210 localMemory_wb_adr_i[6] vssd1 vssd1 vccd1 vccd1 input210/X sky130_fd_sc_hd__clkbuf_1
XFILLER_310_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput221 localMemory_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input221/X sky130_fd_sc_hd__buf_6
Xinput232 localMemory_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 input232/X sky130_fd_sc_hd__buf_8
XTAP_6188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14911_ _14911_/A vssd1 vssd1 vccd1 vccd1 _14911_/X sky130_fd_sc_hd__buf_2
XTAP_6199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput243 localMemory_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input243/X sky130_fd_sc_hd__buf_4
XFILLER_209_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput254 manufacturerID[10] vssd1 vssd1 vccd1 vccd1 input254/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15891_ _15891_/A _15891_/B vssd1 vssd1 vccd1 vccd1 _15891_/Y sky130_fd_sc_hd__nand2_2
Xinput265 partID[10] vssd1 vssd1 vccd1 vccd1 input265/X sky130_fd_sc_hd__clkbuf_1
XTAP_5476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput276 partID[6] vssd1 vssd1 vccd1 vccd1 input276/X sky130_fd_sc_hd__clkbuf_1
X_17630_ _18856_/A vssd1 vssd1 vccd1 vccd1 _17630_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_248_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ _14840_/X _15133_/B _15133_/A vssd1 vssd1 vccd1 vccd1 _14843_/B sky130_fd_sc_hd__mux2_1
XFILLER_75_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17561_ _17561_/A vssd1 vssd1 vccd1 vccd1 _22682_/D sky130_fd_sc_hd__clkbuf_1
X_11985_ _23476_/Q _23572_/Q _22536_/Q _22340_/Q _11637_/X _12793_/A vssd1 vssd1 vccd1
+ vccd1 _11986_/B sky130_fd_sc_hd__mux4_1
XFILLER_263_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14773_ _14772_/X _14626_/X _15132_/S vssd1 vssd1 vccd1 vccd1 _14774_/A sky130_fd_sc_hd__mux2_2
XFILLER_95_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19300_ _19210_/X _23315_/Q _19300_/S vssd1 vssd1 vccd1 vccd1 _19301_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16512_ _16512_/A vssd1 vssd1 vccd1 vccd1 _22412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13724_ _13724_/A _14089_/A vssd1 vssd1 vccd1 vccd1 _14019_/C sky130_fd_sc_hd__nor2_2
X_17492_ _22654_/Q _16233_/X _17494_/S vssd1 vssd1 vccd1 vccd1 _17493_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19231_ _19229_/X _23289_/Q _19243_/S vssd1 vssd1 vccd1 vccd1 _19232_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16443_ _15975_/X _22382_/Q _16451_/S vssd1 vssd1 vccd1 vccd1 _16444_/A sky130_fd_sc_hd__mux2_1
X_13655_ _13655_/A vssd1 vssd1 vccd1 vccd1 _13765_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_204_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19162_ _19162_/A vssd1 vssd1 vccd1 vccd1 _23268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12606_ _12606_/A _12606_/B vssd1 vssd1 vccd1 vccd1 _13353_/B sky130_fd_sc_hd__or2_1
X_16374_ _16374_/A vssd1 vssd1 vccd1 vccd1 _22352_/D sky130_fd_sc_hd__clkbuf_1
X_13586_ _23934_/Q vssd1 vssd1 vccd1 vccd1 _17229_/A sky130_fd_sc_hd__buf_4
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18113_ _22876_/Q _17956_/A _18053_/A _23009_/Q _18054_/A vssd1 vssd1 vccd1 vccd1
+ _18113_/X sky130_fd_sc_hd__a221o_1
X_15325_ _16198_/S vssd1 vssd1 vccd1 vccd1 _15524_/S sky130_fd_sc_hd__buf_4
X_12537_ _22293_/Q _23429_/Q _12537_/S vssd1 vssd1 vccd1 vccd1 _12538_/B sky130_fd_sc_hd__mux2_1
XFILLER_318_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_307_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19093_ _19161_/S vssd1 vssd1 vccd1 vccd1 _19102_/S sky130_fd_sc_hd__buf_6
XFILLER_346_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_318_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18044_ _21220_/A vssd1 vssd1 vccd1 vccd1 _18105_/A sky130_fd_sc_hd__clkbuf_4
X_15256_ _15256_/A _15256_/B vssd1 vssd1 vccd1 vccd1 _15256_/X sky130_fd_sc_hd__or2_1
X_12468_ _12544_/B _12468_/B _13699_/B vssd1 vssd1 vccd1 vccd1 _12468_/X sky130_fd_sc_hd__or3_1
XFILLER_315_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11419_ _22291_/Q _23107_/Q _23523_/Q _22452_/Q _11157_/X _11418_/X vssd1 vssd1 vccd1
+ vccd1 _11420_/B sky130_fd_sc_hd__mux4_1
X_14207_ _14207_/A _14207_/B vssd1 vssd1 vccd1 vccd1 _19922_/D sky130_fd_sc_hd__nor2_8
X_15187_ _15187_/A _15187_/B vssd1 vssd1 vccd1 vccd1 _15484_/B sky130_fd_sc_hd__nand2_2
XFILLER_299_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12399_ _12406_/A _12398_/X _11282_/A vssd1 vssd1 vccd1 vccd1 _12399_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_299_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_334_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_298_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_302_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14138_ _14138_/A vssd1 vssd1 vccd1 vccd1 _15416_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_334_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19995_ _20027_/A _20009_/B vssd1 vssd1 vccd1 vccd1 _19995_/Y sky130_fd_sc_hd__nor2_1
XFILLER_302_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_301_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_330_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18946_ _19164_/A _19018_/B vssd1 vssd1 vccd1 vccd1 _19003_/A sky130_fd_sc_hd__or2_4
X_14069_ _14074_/B _14069_/B _14069_/C vssd1 vssd1 vccd1 vccd1 _14069_/X sky130_fd_sc_hd__or3_1
XTAP_7390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18877_ _23141_/Q _18769_/X _18885_/S vssd1 vssd1 vccd1 vccd1 _18878_/A sky130_fd_sc_hd__mux2_1
XFILLER_254_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17828_ _17874_/S vssd1 vssd1 vccd1 vccd1 _17837_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_227_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17759_ _22756_/Q _17582_/X _17765_/S vssd1 vssd1 vccd1 vccd1 _17760_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_183_wb_clk_i _23931_/CLK vssd1 vssd1 vccd1 vccd1 _23934_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20770_ _20770_/A _21097_/B vssd1 vssd1 vccd1 vccd1 _20864_/A sky130_fd_sc_hd__nor2_8
XFILLER_223_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_340 _17129_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_112_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23005_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XINSDIODE2_351 _22029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19429_ _23372_/Q _18795_/X _19433_/S vssd1 vssd1 vccd1 vccd1 _19430_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_362 _23785_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_373 _23465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_384 _22492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_356_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_395 _14090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22440_ _23511_/CLK _22440_/D vssd1 vssd1 vccd1 vccd1 _22440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_309_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22371_ _23444_/CLK _22371_/D vssd1 vssd1 vccd1 vccd1 _22371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21322_ _21466_/A vssd1 vssd1 vccd1 vccd1 _21575_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21253_ _15671_/X _21196_/X _21252_/X vssd1 vssd1 vccd1 vccd1 _23897_/D sky130_fd_sc_hd__o21ba_2
XFILLER_191_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_305_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20204_ _20146_/X _20585_/A _20202_/X _20203_/X vssd1 vssd1 vccd1 vccd1 _23657_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21184_ _20759_/A _21158_/X _21142_/A _20520_/C _21150_/A vssd1 vssd1 vccd1 vccd1
+ _21184_/X sky130_fd_sc_hd__a221o_1
XFILLER_278_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20135_ _23651_/Q _20136_/C _23652_/Q vssd1 vssd1 vccd1 vccd1 _20137_/B sky130_fd_sc_hd__a21oi_1
XFILLER_131_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20066_ _20066_/A _20066_/B _20066_/C _20076_/D vssd1 vssd1 vccd1 vccd1 _20071_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_286_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_11 _22217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_22 _22254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_33 _18708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_44 _20749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_55 _21400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_66 _21625_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_77 _21898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_88 _20387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23825_ _23878_/CLK _23825_/D vssd1 vssd1 vccd1 vccd1 _23825_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_99 _21648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23756_ _23824_/CLK _23756_/D vssd1 vssd1 vccd1 vccd1 _23756_/Q sky130_fd_sc_hd__dfxtp_2
X_11770_ _11770_/A vssd1 vssd1 vccd1 vccd1 _12070_/S sky130_fd_sc_hd__buf_4
XFILLER_199_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20968_ _23805_/Q _20953_/X _20967_/X _20964_/X vssd1 vssd1 vccd1 vccd1 _23805_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22707_ _23586_/CLK _22707_/D vssd1 vssd1 vccd1 vccd1 _22707_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23687_ _23696_/CLK _23687_/D vssd1 vssd1 vccd1 vccd1 _23687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20899_ _23781_/Q _20893_/X _20898_/X _20788_/X vssd1 vssd1 vccd1 vccd1 _23781_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13440_ _13440_/A _13440_/B _13440_/C _21335_/A vssd1 vssd1 vccd1 vccd1 _20214_/B
+ sky130_fd_sc_hd__nand4_4
X_22638_ _23581_/CLK _22638_/D vssd1 vssd1 vccd1 vccd1 _22638_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13371_ _13371_/A _13371_/B _13371_/C vssd1 vssd1 vccd1 vccd1 _13372_/B sky130_fd_sc_hd__and3_1
X_22569_ _23646_/CLK _22569_/D vssd1 vssd1 vccd1 vccd1 _22569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15110_ input148/X input113/X _15110_/S vssd1 vssd1 vccd1 vccd1 _15110_/X sky130_fd_sc_hd__mux2_8
X_12322_ _12318_/A _12319_/X _12321_/X _11347_/A vssd1 vssd1 vccd1 vccd1 _12322_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_315_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16090_ _16089_/X _22289_/Q _16125_/S vssd1 vssd1 vccd1 vccd1 _16091_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15041_ _15746_/A vssd1 vssd1 vccd1 vccd1 _15041_/X sky130_fd_sc_hd__buf_2
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12253_ _23403_/Q _23019_/Q _23371_/Q _23339_/Q _11113_/A _12199_/X vssd1 vssd1 vccd1
+ vccd1 _12253_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11204_ _13089_/A vssd1 vssd1 vccd1 vccd1 _11205_/A sky130_fd_sc_hd__buf_4
XFILLER_79_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12184_ _22784_/Q _22752_/Q _22653_/Q _22720_/Q _11112_/A _12458_/A vssd1 vssd1 vccd1
+ vccd1 _12184_/X sky130_fd_sc_hd__mux4_2
XFILLER_351_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18800_ _18800_/A vssd1 vssd1 vccd1 vccd1 _23117_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11135_ _11135_/A vssd1 vssd1 vccd1 vccd1 _15864_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_150_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19780_ _23528_/Q _19175_/A _19782_/S vssd1 vssd1 vccd1 vccd1 _19781_/A sky130_fd_sc_hd__mux2_1
X_16992_ _17222_/B vssd1 vssd1 vccd1 vccd1 _17009_/S sky130_fd_sc_hd__buf_2
XFILLER_205_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18731_ _18731_/A vssd1 vssd1 vccd1 vccd1 _23091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15943_ _15575_/X _15243_/Y _15942_/X vssd1 vssd1 vccd1 vccd1 _21269_/A sky130_fd_sc_hd__a21oi_4
X_11066_ _23879_/Q vssd1 vssd1 vccd1 vccd1 _11069_/D sky130_fd_sc_hd__buf_4
XFILLER_62_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18662_ _18662_/A vssd1 vssd1 vccd1 vccd1 _23060_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15874_ _22937_/Q _15000_/X _15001_/X _18427_/A vssd1 vssd1 vccd1 vccd1 _15874_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_5295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_292_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17613_ _17613_/A vssd1 vssd1 vccd1 vccd1 _22698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14825_ input153/X _13650_/A _14719_/S input117/X _14235_/X vssd1 vssd1 vccd1 vccd1
+ _14825_/X sky130_fd_sc_hd__a221o_4
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18593_ _16870_/X _23030_/Q _18597_/S vssd1 vssd1 vccd1 vccd1 _18594_/A sky130_fd_sc_hd__mux2_1
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17544_ _18769_/A vssd1 vssd1 vccd1 vccd1 _17544_/X sky130_fd_sc_hd__clkbuf_2
X_14756_ _14727_/X _14728_/X _14751_/X _14754_/X _14755_/X vssd1 vssd1 vccd1 vccd1
+ _14756_/X sky130_fd_sc_hd__o32a_4
XFILLER_233_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11968_ _23316_/Q _23284_/Q _23252_/Q _23540_/Q _12825_/A _12756_/A vssd1 vssd1 vccd1
+ vccd1 _11969_/B sky130_fd_sc_hd__mux4_2
XFILLER_189_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13707_ _14970_/S vssd1 vssd1 vccd1 vccd1 _13781_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17475_ _22646_/Q _16200_/X _17483_/S vssd1 vssd1 vccd1 vccd1 _17476_/A sky130_fd_sc_hd__mux2_1
X_11899_ _11890_/Y _11892_/Y _11896_/Y _11898_/Y _11215_/A vssd1 vssd1 vccd1 vccd1
+ _11909_/B sky130_fd_sc_hd__o221a_1
X_14687_ _14687_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14687_/X sky130_fd_sc_hd__and2_1
X_19214_ _19246_/A vssd1 vssd1 vccd1 vccd1 _19227_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_340_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16426_ _16426_/A vssd1 vssd1 vccd1 vccd1 _22374_/D sky130_fd_sc_hd__clkbuf_1
X_13638_ _22611_/Q _13718_/D _14089_/B vssd1 vssd1 vccd1 vccd1 _13639_/C sky130_fd_sc_hd__or3_1
XFILLER_301_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19145_ _19145_/A vssd1 vssd1 vccd1 vccd1 _23260_/D sky130_fd_sc_hd__clkbuf_1
X_16357_ _16368_/A vssd1 vssd1 vccd1 vccd1 _16366_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13569_ _13569_/A _13569_/B vssd1 vssd1 vccd1 vccd1 _13570_/B sky130_fd_sc_hd__xnor2_4
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15308_ _14592_/X _15301_/X _15307_/X _14498_/X vssd1 vssd1 vccd1 vccd1 _15308_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19076_ _16895_/X _23230_/Q _19084_/S vssd1 vssd1 vccd1 vccd1 _19077_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16288_ _16288_/A vssd1 vssd1 vccd1 vccd1 _16301_/S sky130_fd_sc_hd__buf_6
XFILLER_172_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18027_ hold2/A _18016_/X _18026_/X _18000_/X vssd1 vssd1 vccd1 vccd1 _22847_/D sky130_fd_sc_hd__o211a_1
X_15239_ _18798_/A vssd1 vssd1 vccd1 vccd1 _19191_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_315_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_303_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_303_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19978_ _23606_/Q _23605_/Q _19978_/C _19978_/D vssd1 vssd1 vccd1 vccd1 _20005_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_262_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18929_ _23165_/Q _18849_/X _18929_/S vssd1 vssd1 vccd1 vccd1 _18930_/A sky130_fd_sc_hd__mux2_1
XFILLER_262_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21940_ _22038_/A _21940_/B vssd1 vssd1 vccd1 vccd1 _21940_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_83_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21871_ _21871_/A _22045_/A vssd1 vssd1 vccd1 vccd1 _21871_/Y sky130_fd_sc_hd__nand2_1
XFILLER_243_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23610_ _23643_/CLK _23610_/D vssd1 vssd1 vccd1 vccd1 _23610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_282_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20822_ _20825_/A _20822_/B vssd1 vssd1 vccd1 vccd1 _20823_/A sky130_fd_sc_hd__and2_1
XFILLER_54_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23541_ _23541_/CLK _23541_/D vssd1 vssd1 vccd1 vccd1 _23541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20753_ _23745_/Q _20729_/X _20752_/X _20737_/X vssd1 vssd1 vccd1 vccd1 _23745_/D
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_170 _17385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_181 _14043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_192 _13939_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23472_ _23951_/A _23472_/D vssd1 vssd1 vccd1 vccd1 _23472_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_126_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20684_ _23734_/Q _20667_/X _20683_/X _20673_/X vssd1 vssd1 vccd1 vccd1 _23734_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_338_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22423_ _23494_/CLK _22423_/D vssd1 vssd1 vccd1 vccd1 _22423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_338_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_353_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22354_ _23554_/CLK _22354_/D vssd1 vssd1 vccd1 vccd1 _22354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_80_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23422_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21305_ _21984_/A vssd1 vssd1 vccd1 vccd1 _21305_/X sky130_fd_sc_hd__buf_2
XFILLER_136_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_353_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22285_ _23547_/CLK _22285_/D vssd1 vssd1 vccd1 vccd1 _22285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_317_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21236_ _21281_/A vssd1 vssd1 vccd1 vccd1 _21236_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_305_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_321_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21167_ _23870_/Q _21147_/X _21165_/Y _21166_/X _18192_/X vssd1 vssd1 vccd1 vccd1
+ _23870_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_320_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20118_ _23646_/Q _23645_/Q vssd1 vssd1 vccd1 vccd1 _20126_/D sky130_fd_sc_hd__and2_1
XFILLER_293_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21098_ _21124_/A vssd1 vssd1 vccd1 vccd1 _21098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20049_ _20086_/A _20049_/B _20063_/C vssd1 vssd1 vccd1 vccd1 _23626_/D sky130_fd_sc_hd__nor3_1
XFILLER_274_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12940_ _13212_/A _12940_/B vssd1 vssd1 vccd1 vccd1 _12940_/Y sky130_fd_sc_hd__nand2_1
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _12871_/A _12871_/B vssd1 vssd1 vccd1 vccd1 _12871_/Y sky130_fd_sc_hd__nor2_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _14610_/A vssd1 vssd1 vccd1 vccd1 _14922_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _23311_/Q _23279_/Q _23247_/Q _23535_/Q _11821_/X _11317_/A vssd1 vssd1 vccd1
+ vccd1 _11822_/X sky130_fd_sc_hd__mux4_1
X_23808_ _23810_/CLK _23808_/D vssd1 vssd1 vccd1 vccd1 _23808_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _15590_/A vssd1 vssd1 vccd1 vccd1 _15590_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_233_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14541_ _23888_/Q vssd1 vssd1 vccd1 vccd1 _14541_/X sky130_fd_sc_hd__buf_4
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _12269_/A vssd1 vssd1 vccd1 vccd1 _11754_/A sky130_fd_sc_hd__buf_4
XFILLER_324_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23739_ _23874_/CLK _23739_/D vssd1 vssd1 vccd1 vccd1 _23739_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _21078_/B _17259_/X _17291_/S vssd1 vssd1 vccd1 vccd1 _17260_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11684_ _11666_/X _11671_/X _11674_/X _11682_/X _11683_/X vssd1 vssd1 vccd1 vccd1
+ _11685_/C sky130_fd_sc_hd__a221o_2
XFILLER_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14472_ _23717_/Q _23847_/Q _15354_/S vssd1 vssd1 vccd1 vccd1 _14472_/X sky130_fd_sc_hd__mux2_2
XFILLER_41_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_329_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_329_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16211_ _18776_/A vssd1 vssd1 vccd1 vccd1 _16211_/X sky130_fd_sc_hd__buf_2
XFILLER_197_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13423_ _13436_/A _20305_/A vssd1 vssd1 vccd1 vccd1 _14251_/A sky130_fd_sc_hd__nor2_2
X_17191_ input89/X input53/X _17200_/S vssd1 vssd1 vccd1 vccd1 _17191_/X sky130_fd_sc_hd__mux2_8
XFILLER_328_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16142_ _23715_/Q _14905_/A _16141_/X vssd1 vssd1 vccd1 vccd1 _16142_/X sky130_fd_sc_hd__o21a_4
X_13354_ _13510_/B _13354_/B vssd1 vssd1 vccd1 vccd1 _15079_/A sky130_fd_sc_hd__xnor2_1
XFILLER_139_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_347_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12305_ _12565_/A _12304_/X _11844_/X vssd1 vssd1 vccd1 vccd1 _12305_/Y sky130_fd_sc_hd__o21ai_1
X_13285_ _13278_/Y _13280_/Y _13282_/Y _13284_/Y _21898_/A vssd1 vssd1 vccd1 vccd1
+ _13295_/B sky130_fd_sc_hd__o221a_1
XFILLER_154_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16073_ _14690_/X _16058_/X _17289_/A _15436_/X vssd1 vssd1 vccd1 vccd1 _16073_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_108_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19901_ _16287_/X _23582_/Q _19909_/S vssd1 vssd1 vccd1 vccd1 _19902_/A sky130_fd_sc_hd__mux2_1
X_15024_ _14632_/A _15013_/X _15023_/X vssd1 vssd1 vccd1 vccd1 _15024_/X sky130_fd_sc_hd__o21ba_2
X_12236_ _12234_/X _12236_/B vssd1 vssd1 vccd1 vccd1 _13510_/A sky130_fd_sc_hd__and2b_1
XFILLER_30_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19832_ _19832_/A vssd1 vssd1 vccd1 vccd1 _23551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12167_ _12162_/Y _12159_/A _12163_/Y _12166_/X _12112_/A vssd1 vssd1 vccd1 vccd1
+ _12167_/Y sky130_fd_sc_hd__a32oi_1
XFILLER_257_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11118_ _12465_/A _11840_/A _21079_/C vssd1 vssd1 vccd1 vccd1 _20533_/B sky130_fd_sc_hd__or3_4
XFILLER_296_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19763_ _19255_/X _23521_/Q _19765_/S vssd1 vssd1 vccd1 vccd1 _19764_/A sky130_fd_sc_hd__mux2_1
X_12098_ _12091_/A _12095_/X _12097_/X _11681_/A vssd1 vssd1 vccd1 vccd1 _12098_/X
+ sky130_fd_sc_hd__o211a_1
X_16975_ input69/X input54/X _17219_/S vssd1 vssd1 vccd1 vccd1 _16975_/X sky130_fd_sc_hd__mux2_8
XFILLER_283_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18714_ _18714_/A vssd1 vssd1 vccd1 vccd1 _23083_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15926_ _15940_/B _15926_/B vssd1 vssd1 vccd1 vccd1 _15926_/X sky130_fd_sc_hd__or2_2
X_19694_ _19694_/A vssd1 vssd1 vccd1 vccd1 _23490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 coreIndex[6] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_4
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_292_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18645_ _23053_/Q _17572_/X _18647_/S vssd1 vssd1 vccd1 vccd1 _18646_/A sky130_fd_sc_hd__mux2_1
XFILLER_280_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _21077_/B _15672_/X _15855_/X _15856_/X vssd1 vssd1 vccd1 vccd1 _15857_/X
+ sky130_fd_sc_hd__o22a_4
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14808_ _14713_/A _14987_/B _15048_/A vssd1 vssd1 vccd1 vccd1 _14808_/X sky130_fd_sc_hd__o21a_1
XFILLER_18_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18576_ _18576_/A vssd1 vssd1 vccd1 vccd1 _23022_/D sky130_fd_sc_hd__clkbuf_1
X_15788_ _15788_/A vssd1 vssd1 vccd1 vccd1 _22281_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17527_ _22670_/Q _16284_/X _17527_/S vssd1 vssd1 vccd1 vccd1 _17528_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14739_ _23815_/Q _15066_/B _20986_/A vssd1 vssd1 vccd1 vccd1 _14739_/X sky130_fd_sc_hd__or3_1
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17458_ _17458_/A vssd1 vssd1 vccd1 vccd1 _22639_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16409_ _16455_/S vssd1 vssd1 vccd1 vccd1 _16418_/S sky130_fd_sc_hd__buf_4
XFILLER_193_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17389_ _21185_/A vssd1 vssd1 vccd1 vccd1 _22122_/A sky130_fd_sc_hd__buf_12
XFILLER_347_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_353_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_307_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19128_ _19128_/A vssd1 vssd1 vccd1 vccd1 _23252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_319_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_334_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19059_ _19059_/A vssd1 vssd1 vccd1 vccd1 _23222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput300 _13998_/Y vssd1 vssd1 vccd1 vccd1 addr1[6] sky130_fd_sc_hd__buf_2
XFILLER_322_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput311 _13965_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[16] sky130_fd_sc_hd__buf_2
Xoutput322 _13986_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[27] sky130_fd_sc_hd__buf_2
XFILLER_133_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22070_ _22064_/A _21329_/X _18012_/X vssd1 vssd1 vccd1 vccd1 _22071_/B sky130_fd_sc_hd__o21ai_1
Xoutput333 _13754_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[10] sky130_fd_sc_hd__buf_2
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_322_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput344 _13813_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[20] sky130_fd_sc_hd__buf_2
XFILLER_350_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput355 _13873_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[30] sky130_fd_sc_hd__buf_2
XFILLER_259_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput366 _13889_/X vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[2] sky130_fd_sc_hd__buf_2
X_21021_ _20630_/A _21008_/X _21020_/X _21010_/X vssd1 vssd1 vccd1 vccd1 _23823_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_288_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput377 _14033_/X vssd1 vssd1 vccd1 vccd1 din0[12] sky130_fd_sc_hd__buf_2
Xoutput388 _14053_/X vssd1 vssd1 vccd1 vccd1 din0[22] sky130_fd_sc_hd__buf_2
XFILLER_303_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput399 _14016_/X vssd1 vssd1 vccd1 vccd1 din0[3] sky130_fd_sc_hd__buf_2
XFILLER_87_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22972_ _22974_/CLK _22972_/D vssd1 vssd1 vccd1 vccd1 _22972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_347_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21923_ _21081_/A _21908_/X _21914_/X _22061_/A _21922_/Y vssd1 vssd1 vccd1 vccd1
+ _21923_/X sky130_fd_sc_hd__a221o_1
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21854_ _21934_/B _21854_/B vssd1 vssd1 vccd1 vccd1 _21854_/X sky130_fd_sc_hd__xor2_4
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20805_ _20620_/B _20791_/X _20792_/X _23757_/Q vssd1 vssd1 vccd1 vccd1 _20806_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_298_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21785_ _23828_/Q _23762_/Q vssd1 vssd1 vccd1 vccd1 _21786_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_358_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23524_ _23556_/CLK _23524_/D vssd1 vssd1 vccd1 vccd1 _23524_/Q sky130_fd_sc_hd__dfxtp_1
X_20736_ _20757_/A _20736_/B _20736_/C vssd1 vssd1 vccd1 vccd1 _20736_/X sky130_fd_sc_hd__or3_1
XFILLER_298_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_329_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23455_ _23582_/CLK _23455_/D vssd1 vssd1 vccd1 vccd1 _23455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20667_ _20729_/A vssd1 vssd1 vccd1 vccd1 _20667_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_338_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22406_ _23542_/CLK _22406_/D vssd1 vssd1 vccd1 vccd1 _22406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23386_ _23420_/CLK _23386_/D vssd1 vssd1 vccd1 vccd1 _23386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_337_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20598_ _20662_/A vssd1 vssd1 vccd1 vccd1 _20598_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_192_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22337_ _23504_/CLK _22337_/D vssd1 vssd1 vccd1 vccd1 _22337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_313_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13070_ _22384_/Q _22416_/Q _22705_/Q _23072_/Q _11311_/A _11323_/A vssd1 vssd1 vccd1
+ vccd1 _13070_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22268_ _23500_/CLK _22268_/D vssd1 vssd1 vccd1 vccd1 _22268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12021_ _23411_/Q _23027_/Q _23379_/Q _23347_/Q _12013_/X _12717_/A vssd1 vssd1 vccd1
+ vccd1 _12021_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21219_ _13440_/A _21202_/X _21217_/Y _21218_/X vssd1 vssd1 vccd1 vccd1 _23885_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22199_ _21307_/X _22184_/X _22191_/X _22198_/X _21410_/X vssd1 vssd1 vccd1 vccd1
+ _22199_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_333_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_294_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16760_ _16760_/A vssd1 vssd1 vccd1 vccd1 _22505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13972_ _13972_/A _13979_/B vssd1 vssd1 vccd1 vccd1 _13973_/A sky130_fd_sc_hd__and2_1
XFILLER_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15711_ _15710_/X _22279_/Q _15750_/S vssd1 vssd1 vccd1 vccd1 _15712_/A sky130_fd_sc_hd__mux2_1
XFILLER_247_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12923_ _11195_/A _12922_/X _12683_/A vssd1 vssd1 vccd1 vccd1 _12923_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16691_ _16691_/A _16806_/B vssd1 vssd1 vccd1 vccd1 _16784_/A sky130_fd_sc_hd__or2_4
XFILLER_46_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_261_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18430_ _18441_/A _18435_/C vssd1 vssd1 vccd1 vccd1 _18430_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15642_ _22963_/Q vssd1 vssd1 vccd1 vccd1 _15644_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _12707_/X _12846_/X _12849_/X _12853_/X _11378_/A vssd1 vssd1 vccd1 vccd1
+ _12864_/B sky130_fd_sc_hd__a311o_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _22947_/Q _18359_/B _18360_/Y vssd1 vssd1 vccd1 vccd1 _22947_/D sky130_fd_sc_hd__o21a_1
X_11805_ _23215_/Q _23183_/Q _23151_/Q _23119_/Q _11799_/X _11800_/X vssd1 vssd1 vccd1
+ vccd1 _11806_/B sky130_fd_sc_hd__mux4_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _15573_/A vssd1 vssd1 vccd1 vccd1 _22276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _23415_/Q _23031_/Q _23383_/Q _23351_/Q _11308_/A _11320_/A vssd1 vssd1 vccd1
+ vccd1 _12785_/X sky130_fd_sc_hd__mux4_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_348_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _17242_/A _17305_/X _17311_/X _16997_/X vssd1 vssd1 vccd1 vccd1 _17312_/X
+ sky130_fd_sc_hd__o211a_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ _14815_/C _14524_/B vssd1 vssd1 vccd1 vccd1 _15478_/A sky130_fd_sc_hd__and2_2
X_18292_ _18423_/A vssd1 vssd1 vccd1 vccd1 _18292_/X sky130_fd_sc_hd__clkbuf_4
X_11736_ _12139_/A _11736_/B vssd1 vssd1 vccd1 vccd1 _11736_/Y sky130_fd_sc_hd__nor2_1
XFILLER_187_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17243_ input94/X input59/X _17266_/S vssd1 vssd1 vccd1 vccd1 _17243_/X sky130_fd_sc_hd__mux2_8
X_14455_ _14455_/A vssd1 vssd1 vccd1 vccd1 _14455_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11667_ _11745_/A vssd1 vssd1 vccd1 vccd1 _12024_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_179_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13406_ _13561_/A _13406_/B vssd1 vssd1 vccd1 vccd1 _13406_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_127_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17174_ _21846_/A _17174_/B vssd1 vssd1 vccd1 vccd1 _17174_/Y sky130_fd_sc_hd__nand2_1
XFILLER_316_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11598_ _12371_/A vssd1 vssd1 vccd1 vccd1 _11598_/X sky130_fd_sc_hd__buf_2
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14386_ _15346_/B vssd1 vssd1 vccd1 vccd1 _16186_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_316_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16125_ _16124_/X _22290_/Q _16125_/S vssd1 vssd1 vccd1 vccd1 _16126_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13337_ _13337_/A vssd1 vssd1 vccd1 vccd1 _13646_/A sky130_fd_sc_hd__buf_6
XFILLER_316_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16056_ _16097_/A _14861_/X _16055_/X _13301_/A vssd1 vssd1 vccd1 vccd1 _16056_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_288_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13268_ _13268_/A _13268_/B vssd1 vssd1 vccd1 vccd1 _13268_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15007_ _15918_/S vssd1 vssd1 vccd1 vccd1 _16053_/S sky130_fd_sc_hd__clkbuf_2
X_12219_ _12208_/X _12212_/X _12214_/X _12218_/X _11375_/A vssd1 vssd1 vccd1 vccd1
+ _12229_/B sky130_fd_sc_hd__a221o_1
XFILLER_331_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13199_ _13199_/A _13199_/B vssd1 vssd1 vccd1 vccd1 _13199_/X sky130_fd_sc_hd__or2_1
XFILLER_170_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_296_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19815_ _23544_/Q _19226_/A _19815_/S vssd1 vssd1 vccd1 vccd1 _19816_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19746_ _19229_/X _23513_/Q _19754_/S vssd1 vssd1 vccd1 vccd1 _19747_/A sky130_fd_sc_hd__mux2_1
X_16958_ _22249_/D _16958_/B _22246_/A vssd1 vssd1 vccd1 vccd1 _21294_/C sky130_fd_sc_hd__or3_1
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_323_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15909_ _23837_/Q _14907_/A _15905_/X _15908_/X _14923_/A vssd1 vssd1 vccd1 vccd1
+ _15909_/X sky130_fd_sc_hd__a221o_1
X_19677_ _19677_/A vssd1 vssd1 vccd1 vccd1 _23482_/D sky130_fd_sc_hd__clkbuf_1
X_16889_ _19239_/A vssd1 vssd1 vccd1 vccd1 _16889_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_225_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18628_ _23045_/Q _17544_/X _18636_/S vssd1 vssd1 vccd1 vccd1 _18629_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_307_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18559_ _18559_/A vssd1 vssd1 vccd1 vccd1 _23014_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_19_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23559_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_162_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21570_ _21570_/A _21576_/A vssd1 vssd1 vccd1 vccd1 _21572_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20521_ _23712_/Q _20523_/B _20521_/C vssd1 vssd1 vccd1 vccd1 _20525_/A sky130_fd_sc_hd__and3_1
XFILLER_166_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_308_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23240_ _23528_/CLK _23240_/D vssd1 vssd1 vccd1 vccd1 _23240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20452_ _20660_/A _20447_/X _20451_/X _20445_/X vssd1 vssd1 vccd1 vccd1 _23699_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_354_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23171_ _23459_/CLK _23171_/D vssd1 vssd1 vccd1 vccd1 _23171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20383_ _20396_/A _20383_/B vssd1 vssd1 vccd1 vccd1 _20383_/X sky130_fd_sc_hd__or2_1
XFILLER_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_334_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22122_ _22122_/A vssd1 vssd1 vccd1 vccd1 _22122_/X sky130_fd_sc_hd__clkbuf_2
XTAP_7219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22053_ _22053_/A _22155_/A vssd1 vssd1 vccd1 vccd1 _22053_/Y sky130_fd_sc_hd__xnor2_1
XTAP_6529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_294_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21004_ _23817_/Q _21009_/B vssd1 vssd1 vccd1 vccd1 _21004_/X sky130_fd_sc_hd__or2_1
XFILLER_287_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22955_ _23602_/CLK _22955_/D vssd1 vssd1 vccd1 vccd1 _22955_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_260_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21906_ _21936_/A _21936_/B _21879_/A _21879_/B vssd1 vssd1 vccd1 vccd1 _21907_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22886_ _23552_/CLK _22886_/D vssd1 vssd1 vccd1 vccd1 _22886_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_204_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21837_ _21837_/A _21837_/B vssd1 vssd1 vccd1 vccd1 _21838_/B sky130_fd_sc_hd__xnor2_1
XPHY_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ _12570_/A _12570_/B vssd1 vssd1 vccd1 vccd1 _12570_/X sky130_fd_sc_hd__or2_1
XFILLER_358_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21768_ _21515_/B _21765_/X _21766_/Y _21767_/X vssd1 vssd1 vccd1 vccd1 _21768_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23507_ _23507_/CLK _23507_/D vssd1 vssd1 vccd1 vccd1 _23507_/Q sky130_fd_sc_hd__dfxtp_1
X_11521_ _13064_/A _11521_/B vssd1 vssd1 vccd1 vccd1 _11521_/X sky130_fd_sc_hd__or2_1
XFILLER_212_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20719_ _15864_/X _20692_/X _20702_/X vssd1 vssd1 vccd1 vccd1 _20719_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_358_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21699_ _21942_/A _21699_/B vssd1 vssd1 vccd1 vccd1 _21699_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14240_ input141/X input169/X _15052_/S vssd1 vssd1 vccd1 vccd1 _14240_/X sky130_fd_sc_hd__mux2_8
X_11452_ _13273_/A _11452_/B vssd1 vssd1 vccd1 vccd1 _11452_/Y sky130_fd_sc_hd__nand2_1
XFILLER_345_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23438_ _23502_/CLK _23438_/D vssd1 vssd1 vccd1 vccd1 _23438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14171_ _14745_/A vssd1 vssd1 vccd1 vccd1 _15440_/A sky130_fd_sc_hd__clkbuf_8
X_23369_ _23369_/CLK _23369_/D vssd1 vssd1 vccd1 vccd1 _23369_/Q sky130_fd_sc_hd__dfxtp_1
X_11383_ _12520_/S vssd1 vssd1 vccd1 vccd1 _12283_/B sky130_fd_sc_hd__buf_4
XFILLER_341_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_353_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_298_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13122_ _23423_/Q _23039_/Q _23391_/Q _23359_/Q _11311_/A _11323_/A vssd1 vssd1 vccd1
+ vccd1 _13122_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17930_ _22254_/A vssd1 vssd1 vccd1 vccd1 _17930_/X sky130_fd_sc_hd__clkbuf_2
X_13053_ _13095_/A _13052_/X _12816_/X vssd1 vssd1 vccd1 vccd1 _13053_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_97_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12004_ _12171_/A _12170_/A vssd1 vssd1 vccd1 vccd1 _13531_/A sky130_fd_sc_hd__nor2_1
XFILLER_239_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17861_ _17861_/A vssd1 vssd1 vccd1 vccd1 _17870_/S sky130_fd_sc_hd__buf_6
XFILLER_120_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19600_ _19600_/A vssd1 vssd1 vccd1 vccd1 _23448_/D sky130_fd_sc_hd__clkbuf_1
X_16812_ _16808_/C _16811_/X _16704_/A vssd1 vssd1 vccd1 vccd1 _22520_/D sky130_fd_sc_hd__a21oi_1
X_17792_ _22771_/Q _17630_/X _17798_/S vssd1 vssd1 vccd1 vccd1 _17793_/A sky130_fd_sc_hd__mux2_1
XFILLER_289_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19531_ _19531_/A vssd1 vssd1 vccd1 vccd1 _23417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16743_ _16779_/A vssd1 vssd1 vccd1 vccd1 _16759_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13955_ _14224_/B _13965_/B vssd1 vssd1 vccd1 vccd1 _13955_/Y sky130_fd_sc_hd__nor2_1
XFILLER_253_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19462_ _23387_/Q _18843_/X _19466_/S vssd1 vssd1 vccd1 vccd1 _19463_/A sky130_fd_sc_hd__mux2_1
X_12906_ _12906_/A _12906_/B vssd1 vssd1 vccd1 vccd1 _12906_/X sky130_fd_sc_hd__or2_1
X_16674_ _16674_/A vssd1 vssd1 vccd1 vccd1 _22483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13886_ _15119_/A vssd1 vssd1 vccd1 vccd1 _13887_/A sky130_fd_sc_hd__buf_4
XFILLER_59_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18413_ _18441_/A _18418_/C vssd1 vssd1 vccd1 vccd1 _18413_/Y sky130_fd_sc_hd__nor2_1
XFILLER_185_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15625_ _19217_/A vssd1 vssd1 vccd1 vccd1 _15625_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_234_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19393_ _19393_/A vssd1 vssd1 vccd1 vccd1 _23356_/D sky130_fd_sc_hd__clkbuf_1
X_12837_ _12830_/Y _12832_/Y _12834_/Y _12836_/Y _11559_/X vssd1 vssd1 vccd1 vccd1
+ _12837_/X sky130_fd_sc_hd__o221a_1
XFILLER_34_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _18360_/A _18349_/C vssd1 vssd1 vccd1 vccd1 _18344_/Y sky130_fd_sc_hd__nor2_1
X_15556_ _14730_/A _15549_/X _15555_/Y _15150_/A vssd1 vssd1 vccd1 vccd1 _15557_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_187_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _22279_/Q _23095_/Q _23511_/Q _22440_/Q _12755_/X _12756_/X vssd1 vssd1 vccd1
+ vccd1 _12769_/B sky130_fd_sc_hd__mux4_2
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14931_/A vssd1 vssd1 vccd1 vccd1 _14752_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_203_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18275_ _18275_/A _22919_/Q _18275_/C vssd1 vssd1 vccd1 vccd1 _18276_/C sky130_fd_sc_hd__and3_1
X_11719_ _11719_/A vssd1 vssd1 vccd1 vccd1 _11777_/S sky130_fd_sc_hd__buf_4
XFILLER_348_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15487_ _14833_/A _15483_/Y _15486_/Y _15183_/A vssd1 vssd1 vccd1 vccd1 _21240_/A
+ sky130_fd_sc_hd__a22o_4
X_12699_ _23480_/Q _23576_/Q _22540_/Q _22344_/Q _12750_/S _12041_/X vssd1 vssd1 vccd1
+ vccd1 _12699_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17226_ _17167_/A _17219_/X _18449_/B _16996_/X _17109_/A vssd1 vssd1 vccd1 vccd1
+ _17226_/X sky130_fd_sc_hd__o221a_4
X_14438_ _14500_/A _14506_/B _15068_/C vssd1 vssd1 vccd1 vccd1 _14588_/A sky130_fd_sc_hd__nor3_2
XFILLER_175_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput10 core_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput21 core_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_1
Xinput32 core_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
Xinput43 dout0[0] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_2
XFILLER_317_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput54 dout0[1] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__buf_2
XFILLER_128_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17157_ _23477_/Q _17170_/B vssd1 vssd1 vccd1 vccd1 _17157_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14369_ _14369_/A _14373_/A vssd1 vssd1 vccd1 vccd1 _14369_/X sky130_fd_sc_hd__or2b_1
Xinput65 dout0[2] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__buf_2
Xinput76 dout0[3] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__buf_2
XFILLER_332_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput87 dout0[4] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__buf_2
X_16108_ _14592_/A _16101_/X _16107_/Y _15652_/X vssd1 vssd1 vccd1 vccd1 _16109_/B
+ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_leaf_137_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _23693_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput98 dout0[5] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__buf_2
X_17088_ _17073_/X _17087_/X _16968_/X _17078_/X vssd1 vssd1 vccd1 vccd1 _17088_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_143_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_289_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16039_ _23938_/Q _17267_/A _16039_/C vssd1 vssd1 vccd1 vccd1 _16077_/B sky130_fd_sc_hd__and3_1
XFILLER_276_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_297_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19729_ _19729_/A vssd1 vssd1 vccd1 vccd1 _23505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22740_ _23391_/CLK _22740_/D vssd1 vssd1 vccd1 vccd1 _22740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_344_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22671_ _23549_/CLK _22671_/D vssd1 vssd1 vccd1 vccd1 _22671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21622_ _21689_/A _21689_/B vssd1 vssd1 vccd1 vccd1 _21624_/B sky130_fd_sc_hd__or2_1
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21553_ _21553_/A vssd1 vssd1 vccd1 vccd1 _21842_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_165_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20504_ _21549_/A vssd1 vssd1 vccd1 vccd1 _21605_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_166_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21484_ _21480_/X _21481_/X _21526_/C vssd1 vssd1 vccd1 vccd1 _21542_/A sky130_fd_sc_hd__mux2_2
X_23223_ _23511_/CLK _23223_/D vssd1 vssd1 vccd1 vccd1 _23223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_342_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20435_ _20470_/A vssd1 vssd1 vccd1 vccd1 _20448_/B sky130_fd_sc_hd__buf_2
XFILLER_308_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_351_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23154_ _23538_/CLK _23154_/D vssd1 vssd1 vccd1 vccd1 _23154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_351_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_350_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20366_ _23678_/Q _20391_/B vssd1 vssd1 vccd1 vccd1 _20366_/X sky130_fd_sc_hd__or2_1
XTAP_7016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22105_ _23807_/Q _21746_/X _22104_/Y _21395_/X vssd1 vssd1 vccd1 vccd1 _22105_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_7049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_350_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23085_ _23565_/CLK _23085_/D vssd1 vssd1 vccd1 vccd1 _23085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20297_ _15606_/Y _20295_/X _20296_/Y vssd1 vssd1 vccd1 vccd1 _20297_/Y sky130_fd_sc_hd__o21ai_1
XTAP_6326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22036_ _22029_/A _21984_/X _22035_/X _21896_/X vssd1 vssd1 vccd1 vccd1 _23934_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_6359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_330_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13740_ _13778_/A _13730_/X _13771_/B _13739_/X _14006_/C vssd1 vssd1 vccd1 vccd1
+ _13741_/B sky130_fd_sc_hd__a32o_4
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22938_ _23649_/CLK _22938_/D vssd1 vssd1 vccd1 vccd1 _22938_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13671_ _14002_/A _16534_/B vssd1 vssd1 vccd1 vccd1 _13671_/Y sky130_fd_sc_hd__nand2_1
X_22869_ _23632_/CLK _22869_/D vssd1 vssd1 vccd1 vccd1 _22869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15410_ _14569_/A _21235_/A _15409_/X _15698_/A vssd1 vssd1 vccd1 vccd1 _15410_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_12622_ _22277_/Q _23093_/Q _23509_/Q _22438_/Q _12013_/X _12710_/A vssd1 vssd1 vccd1
+ vccd1 _12622_/X sky130_fd_sc_hd__mux4_2
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16390_ _14706_/X _22358_/Q _16396_/S vssd1 vssd1 vccd1 vccd1 _16391_/A sky130_fd_sc_hd__mux2_1
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15341_ _14947_/Y _15340_/Y _15341_/S vssd1 vssd1 vccd1 vccd1 _15341_/X sky130_fd_sc_hd__mux2_2
XPHY_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12553_ _12565_/A _12553_/B vssd1 vssd1 vccd1 vccd1 _12553_/X sky130_fd_sc_hd__or2_1
XFILLER_346_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_345_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18060_ _18105_/A vssd1 vssd1 vccd1 vccd1 _18060_/X sky130_fd_sc_hd__clkbuf_2
X_11504_ _11497_/A _11503_/X _11135_/A vssd1 vssd1 vccd1 vccd1 _11504_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_185_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15272_ _15097_/S _15258_/Y _15271_/X _14587_/X vssd1 vssd1 vccd1 vccd1 _15272_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_346_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12484_ _22358_/Q _22390_/Q _22679_/Q _23046_/Q _11919_/A _12216_/A vssd1 vssd1 vccd1
+ vccd1 _12485_/B sky130_fd_sc_hd__mux4_2
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17011_ _17005_/X _17006_/X _17007_/Y _17010_/X _16996_/A vssd1 vssd1 vccd1 vccd1
+ _17011_/X sky130_fd_sc_hd__a221o_1
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14223_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14223_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11435_ _11435_/A vssd1 vssd1 vccd1 vccd1 _11435_/X sky130_fd_sc_hd__buf_6
XFILLER_138_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_326_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14154_ _13670_/C _14151_/X _14152_/X _14153_/X vssd1 vssd1 vccd1 vccd1 _16941_/B
+ sky130_fd_sc_hd__a22o_1
X_11366_ _22292_/Q _23108_/Q _23524_/Q _22453_/Q _11461_/A _11365_/X vssd1 vssd1 vccd1
+ vccd1 _11367_/B sky130_fd_sc_hd__mux4_1
XFILLER_171_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13105_ _13149_/A _13104_/X _12816_/A vssd1 vssd1 vccd1 vccd1 _13105_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_98_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_342_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11297_ _11515_/A vssd1 vssd1 vccd1 vccd1 _13225_/A sky130_fd_sc_hd__clkbuf_8
X_14085_ _14085_/A vssd1 vssd1 vccd1 vccd1 _14085_/Y sky130_fd_sc_hd__inv_2
X_18962_ _16835_/X _23179_/Q _18968_/S vssd1 vssd1 vccd1 vccd1 _18963_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17913_ _22817_/Q _17891_/X _17911_/X _17912_/X vssd1 vssd1 vccd1 vccd1 _22817_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_301_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13036_ _11196_/A _13032_/X _13035_/X vssd1 vssd1 vccd1 vccd1 _13036_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_267_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18893_ _18893_/A vssd1 vssd1 vccd1 vccd1 _23148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17844_ _22794_/Q _17601_/X _17848_/S vssd1 vssd1 vccd1 vccd1 _17845_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17775_ _17775_/A vssd1 vssd1 vccd1 vccd1 _22763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_304_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14987_ _15037_/A _14987_/B vssd1 vssd1 vccd1 vccd1 _14987_/X sky130_fd_sc_hd__or2_1
XFILLER_19_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19514_ _19207_/X _23410_/Q _19516_/S vssd1 vssd1 vccd1 vccd1 _19515_/A sky130_fd_sc_hd__mux2_1
X_16726_ _22496_/Q _16711_/X _16712_/X input41/X vssd1 vssd1 vccd1 vccd1 _16727_/B
+ sky130_fd_sc_hd__o22a_1
X_13938_ _21570_/A vssd1 vssd1 vccd1 vccd1 _13939_/B sky130_fd_sc_hd__buf_8
XFILLER_75_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_500 _15005_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_511 _17143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19445_ _19445_/A vssd1 vssd1 vccd1 vccd1 _23379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_522 _14050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16657_ _16657_/A vssd1 vssd1 vccd1 vccd1 _22475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_533 _23943_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13869_ _13768_/Y _13864_/B _13863_/B _13821_/Y vssd1 vssd1 vccd1 vccd1 _13871_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_320_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_544 _14079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_555 _23473_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15608_ _14822_/X _15579_/X _15607_/Y _14882_/A vssd1 vssd1 vccd1 vccd1 _15608_/X
+ sky130_fd_sc_hd__a22o_1
X_19376_ _19376_/A vssd1 vssd1 vccd1 vccd1 _23348_/D sky130_fd_sc_hd__clkbuf_1
X_16588_ _15898_/X _22445_/Q _16590_/S vssd1 vssd1 vccd1 vccd1 _16589_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18327_ _18360_/A _18332_/C vssd1 vssd1 vccd1 vccd1 _18327_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15539_ _15490_/S _15132_/X _15491_/S vssd1 vssd1 vccd1 vccd1 _15539_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_337_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_349_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18258_ _18263_/A _18263_/B _18257_/Y vssd1 vssd1 vccd1 vccd1 _22915_/D sky130_fd_sc_hd__o21a_1
XFILLER_176_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_318_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17209_ _17276_/A vssd1 vssd1 vccd1 vccd1 _17266_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_352_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18189_ _18195_/A _18195_/C vssd1 vssd1 vccd1 vccd1 _18191_/C sky130_fd_sc_hd__nor2_1
XFILLER_191_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_345_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20220_ _20220_/A vssd1 vssd1 vccd1 vccd1 _20320_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_351_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_333_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20151_ _20216_/A vssd1 vssd1 vccd1 vccd1 _20197_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_170_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_332_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20082_ _20090_/C _20072_/B _20085_/D _18516_/A vssd1 vssd1 vccd1 vccd1 _20082_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_350_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23910_ _23910_/CLK _23910_/D vssd1 vssd1 vccd1 vccd1 _23910_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23841_ _23841_/CLK _23841_/D vssd1 vssd1 vccd1 vccd1 _23841_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_34_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _22666_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23772_ _23776_/CLK _23772_/D vssd1 vssd1 vccd1 vccd1 _23772_/Q sky130_fd_sc_hd__dfxtp_4
X_20984_ _17315_/X _21085_/A _20888_/B _20926_/A vssd1 vssd1 vccd1 vccd1 _20984_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22723_ _23567_/CLK _22723_/D vssd1 vssd1 vccd1 vccd1 _22723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22654_ _23559_/CLK _22654_/D vssd1 vssd1 vccd1 vccd1 _22654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21605_ _21605_/A _21605_/B _21605_/C vssd1 vssd1 vccd1 vccd1 _21605_/X sky130_fd_sc_hd__and3_1
X_22585_ _23693_/CLK _22585_/D vssd1 vssd1 vccd1 vccd1 _22585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_328_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_328_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21536_ _21816_/A vssd1 vssd1 vccd1 vccd1 _22214_/S sky130_fd_sc_hd__buf_4
XFILLER_127_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_327_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21467_ _22171_/B vssd1 vssd1 vccd1 vccd1 _21829_/B sky130_fd_sc_hd__buf_2
XFILLER_147_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11220_ _15864_/A _11172_/Y _11188_/Y _11211_/X _15929_/A vssd1 vssd1 vccd1 vccd1
+ _11249_/B sky130_fd_sc_hd__o311a_1
XFILLER_308_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20418_ _20491_/B vssd1 vssd1 vccd1 vccd1 _20429_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_23206_ _23494_/CLK _23206_/D vssd1 vssd1 vccd1 vccd1 _23206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21398_ _21676_/B vssd1 vssd1 vccd1 vccd1 _21398_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_324_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11151_ _11151_/A vssd1 vssd1 vccd1 vccd1 _12751_/S sky130_fd_sc_hd__buf_6
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23137_ _23553_/CLK _23137_/D vssd1 vssd1 vccd1 vccd1 _23137_/Q sky130_fd_sc_hd__dfxtp_1
X_20349_ _20227_/X _20347_/X _20348_/Y _20320_/X vssd1 vssd1 vccd1 vccd1 _20349_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_323_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_296_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23068_ _23068_/CLK _23068_/D vssd1 vssd1 vccd1 vccd1 _23068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11082_ _13436_/A _13421_/A vssd1 vssd1 vccd1 vccd1 _21335_/C sky130_fd_sc_hd__nand2_4
XFILLER_295_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput200 localMemory_wb_adr_i[19] vssd1 vssd1 vccd1 vccd1 input200/X sky130_fd_sc_hd__clkbuf_1
XTAP_6156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput211 localMemory_wb_adr_i[7] vssd1 vssd1 vccd1 vccd1 input211/X sky130_fd_sc_hd__clkbuf_1
XTAP_6178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput222 localMemory_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input222/X sky130_fd_sc_hd__buf_6
XTAP_5433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22019_ _22019_/A vssd1 vssd1 vccd1 vccd1 _22190_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_48_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14910_ _14910_/A vssd1 vssd1 vccd1 vccd1 _14911_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput233 localMemory_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 input233/X sky130_fd_sc_hd__buf_8
XTAP_6189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15890_ _17229_/A _15924_/C vssd1 vssd1 vccd1 vccd1 _15891_/B sky130_fd_sc_hd__xnor2_2
XFILLER_341_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput244 localMemory_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input244/X sky130_fd_sc_hd__buf_4
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput255 manufacturerID[1] vssd1 vssd1 vccd1 vccd1 input255/X sky130_fd_sc_hd__clkbuf_4
XTAP_5466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput266 partID[11] vssd1 vssd1 vccd1 vccd1 input266/X sky130_fd_sc_hd__clkbuf_1
XFILLER_286_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput277 partID[7] vssd1 vssd1 vccd1 vccd1 input277/X sky130_fd_sc_hd__clkbuf_1
XTAP_5488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ _14664_/X _14653_/A _14841_/S vssd1 vssd1 vccd1 vccd1 _15133_/B sky130_fd_sc_hd__mux2_1
XFILLER_64_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17560_ _22682_/Q _17559_/X _17560_/S vssd1 vssd1 vccd1 vccd1 _17561_/A sky130_fd_sc_hd__mux2_1
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14772_ _14278_/X _14285_/X _14853_/S vssd1 vssd1 vccd1 vccd1 _14772_/X sky130_fd_sc_hd__mux2_1
X_11984_ _12842_/A _11984_/B vssd1 vssd1 vccd1 vccd1 _11984_/X sky130_fd_sc_hd__or2_1
XFILLER_217_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16511_ _15898_/X _22412_/Q _16513_/S vssd1 vssd1 vccd1 vccd1 _16512_/A sky130_fd_sc_hd__mux2_1
X_13723_ _13723_/A vssd1 vssd1 vccd1 vccd1 _13723_/X sky130_fd_sc_hd__clkbuf_1
X_17491_ _17491_/A vssd1 vssd1 vccd1 vccd1 _22653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19230_ _19246_/A vssd1 vssd1 vccd1 vccd1 _19243_/S sky130_fd_sc_hd__clkbuf_4
X_16442_ _16442_/A vssd1 vssd1 vccd1 vccd1 _16451_/S sky130_fd_sc_hd__buf_6
XFILLER_232_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13654_ _14224_/A vssd1 vssd1 vccd1 vccd1 _13993_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_182_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19161_ _23268_/Q _18871_/X _19161_/S vssd1 vssd1 vccd1 vccd1 _19162_/A sky130_fd_sc_hd__mux2_1
X_12605_ _12605_/A vssd1 vssd1 vccd1 vccd1 _12606_/B sky130_fd_sc_hd__clkinv_2
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ _16049_/X _22352_/Q _16377_/S vssd1 vssd1 vccd1 vccd1 _16374_/A sky130_fd_sc_hd__mux2_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _13655_/A vssd1 vssd1 vccd1 vccd1 _13718_/D sky130_fd_sc_hd__clkinv_4
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18112_ _22876_/Q _18051_/A _18111_/X _18105_/X vssd1 vssd1 vccd1 vccd1 _22876_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_223_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_346_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15324_ _19197_/A vssd1 vssd1 vccd1 vccd1 _15324_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19092_ _19148_/A vssd1 vssd1 vccd1 vccd1 _19161_/S sky130_fd_sc_hd__buf_6
X_12536_ _12536_/A _12536_/B vssd1 vssd1 vccd1 vccd1 _12536_/Y sky130_fd_sc_hd__nand2_1
XFILLER_157_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18043_ _22852_/Q _18036_/X _18037_/X _22985_/Q _18038_/X vssd1 vssd1 vccd1 vccd1
+ _18043_/X sky130_fd_sc_hd__a221o_1
XFILLER_333_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15255_ _14264_/X _15251_/X _15850_/B _14384_/X vssd1 vssd1 vccd1 vccd1 _15255_/X
+ sky130_fd_sc_hd__o22a_2
X_12467_ _11241_/A _12454_/X _12461_/X _12466_/X vssd1 vssd1 vccd1 vccd1 _13699_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_8_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14206_ _14206_/A _14207_/B vssd1 vssd1 vccd1 vccd1 _21193_/A sky130_fd_sc_hd__nor2_1
X_11418_ _11418_/A vssd1 vssd1 vccd1 vccd1 _11418_/X sky130_fd_sc_hd__buf_4
X_15186_ _15186_/A _15433_/B vssd1 vssd1 vccd1 vccd1 _15186_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12398_ _23463_/Q _23559_/Q _22523_/Q _22327_/Q _11814_/X _11800_/A vssd1 vssd1 vccd1
+ vccd1 _12398_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14137_ _14137_/A vssd1 vssd1 vccd1 vccd1 _14138_/A sky130_fd_sc_hd__clkbuf_2
X_11349_ _12797_/A vssd1 vssd1 vccd1 vccd1 _12721_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_235_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19994_ _23611_/Q _23610_/Q _19994_/C vssd1 vssd1 vccd1 vccd1 _20009_/B sky130_fd_sc_hd__and3_1
XFILLER_314_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_299_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_298_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18945_ _18945_/A vssd1 vssd1 vccd1 vccd1 _23172_/D sky130_fd_sc_hd__clkbuf_1
X_14068_ _14049_/X _13872_/B _14009_/X input238/X vssd1 vssd1 vccd1 vccd1 _14068_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_113_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_315_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13019_ _13493_/B vssd1 vssd1 vccd1 vccd1 _13019_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18876_ _18944_/S vssd1 vssd1 vccd1 vccd1 _18885_/S sky130_fd_sc_hd__buf_6
XTAP_6690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_267_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17827_ _17827_/A vssd1 vssd1 vccd1 vccd1 _22786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_255_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17758_ _17758_/A vssd1 vssd1 vccd1 vccd1 _22755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16709_ _16723_/A _16709_/B vssd1 vssd1 vccd1 vccd1 _16710_/A sky130_fd_sc_hd__or2_1
XFILLER_235_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17689_ _22725_/Q _17585_/X _17693_/S vssd1 vssd1 vccd1 vccd1 _17690_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_330 _16975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_341 _17133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_352 _22029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19428_ _19428_/A vssd1 vssd1 vccd1 vccd1 _23371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_357_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_363 _23790_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_374 _23467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_385 _22493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_396 _14090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19359_ _23341_/Q _18798_/X _19361_/S vssd1 vssd1 vccd1 vccd1 _19360_/A sky130_fd_sc_hd__mux2_1
XFILLER_349_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22370_ _23570_/CLK _22370_/D vssd1 vssd1 vccd1 vccd1 _22370_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_152_wb_clk_i _23945_/CLK vssd1 vssd1 vccd1 vccd1 _23862_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_176_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_309_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21321_ _21321_/A _21321_/B vssd1 vssd1 vccd1 vccd1 _21466_/A sky130_fd_sc_hd__nand2_2
XFILLER_190_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21252_ _15674_/X _15675_/Y _21242_/A _20058_/X vssd1 vssd1 vccd1 vccd1 _21252_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_340_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_305_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_333_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20203_ _20324_/A vssd1 vssd1 vccd1 vccd1 _20203_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21183_ _23876_/Q _21168_/X _21182_/X _21163_/X vssd1 vssd1 vccd1 vccd1 _23876_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_333_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_321_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20134_ _20134_/A _20134_/B vssd1 vssd1 vccd1 vccd1 _23651_/D sky130_fd_sc_hd__nor2_1
XFILLER_277_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20065_ _23631_/Q vssd1 vssd1 vccd1 vccd1 _20079_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_219_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_12 _17315_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_23 _22254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_34 _18708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_45 _20428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_56 _21400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_67 _21633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_78 _20400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23824_ _23824_/CLK _23824_/D vssd1 vssd1 vccd1 vccd1 _23824_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_89 _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23755_ _23755_/CLK _23755_/D vssd1 vssd1 vccd1 vccd1 _23755_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ _22064_/A _20966_/X _20727_/B _20954_/X vssd1 vssd1 vccd1 vccd1 _20967_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22706_ _23073_/CLK _22706_/D vssd1 vssd1 vccd1 vccd1 _22706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23686_ _23692_/CLK _23686_/D vssd1 vssd1 vccd1 vccd1 _23686_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20898_ _21300_/B _20894_/X _20558_/A _20897_/X vssd1 vssd1 vccd1 vccd1 _20898_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_198_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_328_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22637_ _22666_/CLK _22637_/D vssd1 vssd1 vccd1 vccd1 _22637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13370_ _15079_/A _14940_/A _13370_/C _13370_/D vssd1 vssd1 vccd1 vccd1 _13370_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_142_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22568_ _23646_/CLK _22568_/D vssd1 vssd1 vccd1 vccd1 _22568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12321_ _12321_/A _12321_/B vssd1 vssd1 vccd1 vccd1 _12321_/X sky130_fd_sc_hd__or2_1
XFILLER_355_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21519_ _14195_/X _21518_/X _21615_/A _15161_/B vssd1 vssd1 vccd1 vccd1 _21519_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_357_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22499_ _23704_/CLK _22499_/D vssd1 vssd1 vccd1 vccd1 _22499_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15040_ _22983_/Q _14138_/A _15164_/A input242/X vssd1 vssd1 vccd1 vccd1 _21474_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_170_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12252_ _12256_/A _12252_/B vssd1 vssd1 vccd1 vccd1 _12252_/Y sky130_fd_sc_hd__nor2_1
XFILLER_324_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11203_ _13041_/A vssd1 vssd1 vccd1 vccd1 _13253_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_312_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12183_ _12350_/A _12183_/B vssd1 vssd1 vccd1 vccd1 _12183_/Y sky130_fd_sc_hd__nand2_1
XFILLER_150_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_311_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11134_ _11134_/A vssd1 vssd1 vccd1 vccd1 _11135_/A sky130_fd_sc_hd__buf_4
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16991_ _17248_/A vssd1 vssd1 vccd1 vccd1 _17222_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_296_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18730_ _16860_/X _23091_/Q _18730_/S vssd1 vssd1 vccd1 vccd1 _18731_/A sky130_fd_sc_hd__mux2_1
X_11065_ _23880_/Q vssd1 vssd1 vccd1 vccd1 _11069_/C sky130_fd_sc_hd__buf_4
X_15942_ _15942_/A vssd1 vssd1 vccd1 vccd1 _15942_/X sky130_fd_sc_hd__buf_4
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_295_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18661_ _23060_/Q _17594_/X _18669_/S vssd1 vssd1 vccd1 vccd1 _18662_/A sky130_fd_sc_hd__mux2_1
XTAP_5274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ _22969_/Q vssd1 vssd1 vccd1 vccd1 _18427_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17612_ _22698_/Q _17610_/X _17624_/S vssd1 vssd1 vccd1 vccd1 _17613_/A sky130_fd_sc_hd__mux2_1
X_14824_ _22514_/Q _13691_/A _14238_/X _14823_/X _15056_/A vssd1 vssd1 vccd1 vccd1
+ _15332_/A sky130_fd_sc_hd__o221ai_4
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18592_ _18592_/A vssd1 vssd1 vccd1 vccd1 _23029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_292_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17543_ _17543_/A vssd1 vssd1 vccd1 vccd1 _22677_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ _14755_/A vssd1 vssd1 vccd1 vccd1 _14755_/X sky130_fd_sc_hd__buf_4
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11967_ _12700_/A _11951_/Y _11956_/Y _11960_/Y _11966_/Y vssd1 vssd1 vccd1 vccd1
+ _11967_/X sky130_fd_sc_hd__o32a_1
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13706_ _13706_/A vssd1 vssd1 vccd1 vccd1 _14970_/S sky130_fd_sc_hd__clkbuf_4
X_17474_ _17542_/S vssd1 vssd1 vccd1 vccd1 _17483_/S sky130_fd_sc_hd__buf_6
XFILLER_339_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14686_ _14687_/A _14687_/B _15256_/B vssd1 vssd1 vccd1 vccd1 _14686_/Y sky130_fd_sc_hd__o21ai_1
X_11898_ _11698_/A _11897_/X _11713_/X vssd1 vssd1 vccd1 vccd1 _11898_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19213_ _19213_/A vssd1 vssd1 vccd1 vccd1 _19213_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16425_ _15668_/X _22374_/Q _16429_/S vssd1 vssd1 vccd1 vccd1 _16426_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13637_ _13977_/A _13970_/A _13975_/A _13636_/X vssd1 vssd1 vccd1 vccd1 _14089_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_347_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19144_ _23260_/Q _18846_/X _19146_/S vssd1 vssd1 vccd1 vccd1 _19145_/A sky130_fd_sc_hd__mux2_1
XFILLER_347_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16356_ _16356_/A vssd1 vssd1 vccd1 vccd1 _22344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13568_ _23937_/Q vssd1 vssd1 vccd1 vccd1 _17267_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15307_ _23695_/Q _15210_/X _15306_/X vssd1 vssd1 vccd1 vccd1 _15307_/X sky130_fd_sc_hd__o21a_2
XFILLER_146_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_347_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19075_ _19075_/A vssd1 vssd1 vccd1 vccd1 _19084_/S sky130_fd_sc_hd__buf_4
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12519_ _12519_/A _12519_/B _12519_/C vssd1 vssd1 vccd1 vccd1 _20499_/B sky130_fd_sc_hd__and3_4
XFILLER_118_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16287_ _18852_/A vssd1 vssd1 vccd1 vccd1 _16287_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_334_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13499_ _13499_/A vssd1 vssd1 vccd1 vccd1 _13618_/B sky130_fd_sc_hd__inv_2
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18026_ hold1/A _18017_/X _18020_/X _22979_/Q _18023_/X vssd1 vssd1 vccd1 vccd1 _18026_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_172_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15238_ _11935_/X _15048_/X _15235_/X _21576_/A _15041_/X vssd1 vssd1 vccd1 vccd1
+ _18798_/A sky130_fd_sc_hd__a32o_4
XFILLER_315_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_2_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ _15168_/X _22268_/Q _15284_/S vssd1 vssd1 vccd1 vccd1 _15170_/A sky130_fd_sc_hd__mux2_1
XFILLER_314_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_299_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_287_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19977_ _23600_/Q _19977_/B _19977_/C vssd1 vssd1 vccd1 vccd1 _19978_/D sky130_fd_sc_hd__and3_1
XFILLER_302_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_330_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_302_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18928_ _18928_/A vssd1 vssd1 vccd1 vccd1 _23164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_262_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18859_ _18859_/A vssd1 vssd1 vccd1 vccd1 _18859_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_228_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21870_ _21870_/A vssd1 vssd1 vccd1 vccd1 _22045_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20821_ _20652_/B _20810_/X _20811_/X _23761_/Q vssd1 vssd1 vccd1 vccd1 _20822_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_211_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23540_ _23542_/CLK _23540_/D vssd1 vssd1 vccd1 vccd1 _23540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20752_ _20757_/A _20752_/B _20752_/C vssd1 vssd1 vccd1 vccd1 _20752_/X sky130_fd_sc_hd__or3_1
XFILLER_51_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_160 _13979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_171 _17029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_357_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_182 _14056_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23471_ _23538_/CLK _23471_/D vssd1 vssd1 vccd1 vccd1 _23471_/Q sky130_fd_sc_hd__dfxtp_4
XINSDIODE2_193 _14095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20683_ _20695_/A _20683_/B _20683_/C vssd1 vssd1 vccd1 vccd1 _20683_/X sky130_fd_sc_hd__or3_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22422_ _23903_/CLK _22422_/D vssd1 vssd1 vccd1 vccd1 _22422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_338_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_353_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22353_ _23073_/CLK _22353_/D vssd1 vssd1 vccd1 vccd1 _22353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_353_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21304_ _21410_/A vssd1 vssd1 vccd1 vccd1 _21984_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_352_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22284_ _23100_/CLK _22284_/D vssd1 vssd1 vccd1 vccd1 _22284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_317_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_353_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21235_ _21235_/A _21240_/B vssd1 vssd1 vccd1 vccd1 _21235_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21166_ _21083_/X _20515_/D _21150_/X vssd1 vssd1 vccd1 vccd1 _21166_/X sky130_fd_sc_hd__a21o_1
XFILLER_132_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_321_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20117_ _23645_/Q _20119_/A _23646_/Q vssd1 vssd1 vccd1 vccd1 _20120_/B sky130_fd_sc_hd__a21oi_1
XFILLER_266_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21097_ _21097_/A _21097_/B _21148_/A vssd1 vssd1 vccd1 vccd1 _21124_/A sky130_fd_sc_hd__or3_4
XFILLER_292_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20048_ _23624_/Q _20048_/B _20048_/C _20056_/D vssd1 vssd1 vccd1 vccd1 _20063_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_19_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _22798_/Q _22766_/Q _22667_/Q _22734_/Q _12922_/S _12756_/X vssd1 vssd1 vccd1
+ vccd1 _12871_/B sky130_fd_sc_hd__mux4_2
XFILLER_73_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23807_ _23810_/CLK _23807_/D vssd1 vssd1 vccd1 vccd1 _23807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11821_/A vssd1 vssd1 vccd1 vccd1 _11821_/X sky130_fd_sc_hd__buf_4
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21999_ _21999_/A _22003_/A vssd1 vssd1 vccd1 vccd1 _22000_/B sky130_fd_sc_hd__or2_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _18770_/A vssd1 vssd1 vccd1 vccd1 _17471_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _12139_/A _11751_/X _11284_/A vssd1 vssd1 vccd1 vccd1 _11752_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23738_ _23915_/CLK _23738_/D vssd1 vssd1 vccd1 vccd1 _23738_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_324_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _15806_/S vssd1 vssd1 vccd1 vccd1 _15354_/S sky130_fd_sc_hd__buf_4
XFILLER_230_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11683_ _11683_/A vssd1 vssd1 vccd1 vccd1 _11683_/X sky130_fd_sc_hd__buf_6
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23669_ _23684_/CLK _23669_/D vssd1 vssd1 vccd1 vccd1 _23669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16210_ _16210_/A vssd1 vssd1 vccd1 vccd1 _22293_/D sky130_fd_sc_hd__clkbuf_1
X_13422_ _15425_/A _15080_/A vssd1 vssd1 vccd1 vccd1 _20305_/A sky130_fd_sc_hd__nand2_4
X_17190_ _17324_/A vssd1 vssd1 vccd1 vccd1 _17190_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16141_ _23843_/Q _14907_/A _16137_/X _16140_/X _14922_/A vssd1 vssd1 vccd1 vccd1
+ _16141_/X sky130_fd_sc_hd__a221o_1
XFILLER_127_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13353_ _13928_/A _13353_/B _13353_/C vssd1 vssd1 vccd1 vccd1 _15122_/B sky130_fd_sc_hd__nand3_1
XFILLER_139_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_347_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12304_ _23402_/Q _23018_/Q _23370_/Q _23338_/Q _12245_/S _12292_/X vssd1 vssd1 vccd1
+ vccd1 _12304_/X sky130_fd_sc_hd__mux4_1
XFILLER_344_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16072_ _14518_/A _16060_/X _16071_/X vssd1 vssd1 vccd1 vccd1 _17289_/A sky130_fd_sc_hd__o21ai_4
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13284_ _11343_/A _13283_/X _11288_/A vssd1 vssd1 vccd1 vccd1 _13284_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19900_ _19900_/A vssd1 vssd1 vccd1 vccd1 _19909_/S sky130_fd_sc_hd__buf_6
X_15023_ _14835_/A _13913_/A _15090_/A _15995_/B _15022_/X vssd1 vssd1 vccd1 vccd1
+ _15023_/X sky130_fd_sc_hd__a221o_1
XFILLER_114_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12235_ _12235_/A _12235_/B vssd1 vssd1 vccd1 vccd1 _12236_/B sky130_fd_sc_hd__or2_1
XFILLER_269_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_331_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19831_ _23551_/Q _19249_/A _19837_/S vssd1 vssd1 vccd1 vccd1 _19832_/A sky130_fd_sc_hd__mux2_1
XFILLER_296_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12166_ _21738_/A _12165_/Y _13234_/S vssd1 vssd1 vccd1 vccd1 _12166_/X sky130_fd_sc_hd__mux2_8
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ _23903_/Q _23902_/Q vssd1 vssd1 vccd1 vccd1 _21079_/C sky130_fd_sc_hd__or2_2
X_19762_ _19762_/A vssd1 vssd1 vccd1 vccd1 _23520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16974_ _22553_/Q _16922_/X _16970_/X _16973_/X vssd1 vssd1 vccd1 vccd1 _22553_/D
+ sky130_fd_sc_hd__a211o_1
X_12097_ _12097_/A _12097_/B vssd1 vssd1 vccd1 vccd1 _12097_/X sky130_fd_sc_hd__or2_1
XFILLER_49_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18713_ _16835_/X _23083_/Q _18719_/S vssd1 vssd1 vccd1 vccd1 _18714_/A sky130_fd_sc_hd__mux2_1
XFILLER_283_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15925_ _17229_/A _15924_/C _17246_/A vssd1 vssd1 vccd1 vccd1 _15926_/B sky130_fd_sc_hd__a21oi_1
XFILLER_65_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19693_ _19258_/X _23490_/Q _19693_/S vssd1 vssd1 vccd1 vccd1 _19694_/A sky130_fd_sc_hd__mux2_1
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 coreIndex[7] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_4
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18644_ _18644_/A vssd1 vssd1 vccd1 vccd1 _23052_/D sky130_fd_sc_hd__clkbuf_1
X_15856_ _15162_/A _13601_/Y _14529_/A vssd1 vssd1 vccd1 vccd1 _15856_/X sky130_fd_sc_hd__a21o_1
XFILLER_225_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14807_ _14807_/A vssd1 vssd1 vccd1 vccd1 _14987_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_36_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15787_ _15785_/X _22281_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15788_/A sky130_fd_sc_hd__mux2_1
X_18575_ _16844_/X _23022_/Q _18575_/S vssd1 vssd1 vccd1 vccd1 _18576_/A sky130_fd_sc_hd__mux2_1
X_12999_ _11515_/A _12996_/X _12998_/X _12721_/X vssd1 vssd1 vccd1 vccd1 _12999_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17526_ _17526_/A vssd1 vssd1 vccd1 vccd1 _22669_/D sky130_fd_sc_hd__clkbuf_1
X_14738_ _14922_/A vssd1 vssd1 vccd1 vccd1 _14738_/X sky130_fd_sc_hd__buf_4
XFILLER_339_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_339_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17457_ _22639_/Q _16287_/X _17465_/S vssd1 vssd1 vccd1 vccd1 _17458_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14669_ _14659_/X _14667_/Y _14855_/A vssd1 vssd1 vccd1 vccd1 _14669_/X sky130_fd_sc_hd__mux2_2
XFILLER_221_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16408_ _16408_/A vssd1 vssd1 vccd1 vccd1 _22366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17388_ _20808_/A vssd1 vssd1 vccd1 vccd1 _21185_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_353_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_307_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19127_ _23252_/Q _18820_/X _19135_/S vssd1 vssd1 vccd1 vccd1 _19128_/A sky130_fd_sc_hd__mux2_1
X_16339_ _16339_/A vssd1 vssd1 vccd1 vccd1 _22336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_257_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_346_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_334_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19058_ _16870_/X _23222_/Q _19062_/S vssd1 vssd1 vccd1 vccd1 _19059_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput301 _13999_/Y vssd1 vssd1 vccd1 vccd1 addr1[7] sky130_fd_sc_hd__buf_2
XFILLER_133_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput312 _13966_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[17] sky130_fd_sc_hd__buf_2
X_18009_ _18198_/A _18009_/B _18009_/C _14125_/Y vssd1 vssd1 vccd1 vccd1 _18009_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_322_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput323 _13900_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[2] sky130_fd_sc_hd__buf_2
XFILLER_273_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput334 _13757_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[11] sky130_fd_sc_hd__buf_2
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput345 _13818_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[21] sky130_fd_sc_hd__buf_2
Xoutput356 _13878_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[31] sky130_fd_sc_hd__buf_2
X_21020_ _23823_/Q _21028_/B vssd1 vssd1 vccd1 vccd1 _21020_/X sky130_fd_sc_hd__or2_1
XFILLER_299_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput367 _13892_/Y vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[3] sky130_fd_sc_hd__buf_2
XFILLER_302_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput378 _14035_/X vssd1 vssd1 vccd1 vccd1 din0[13] sky130_fd_sc_hd__buf_2
XFILLER_288_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput389 _14054_/X vssd1 vssd1 vccd1 vccd1 din0[23] sky130_fd_sc_hd__buf_2
XFILLER_87_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22971_ _22971_/CLK _22971_/D vssd1 vssd1 vccd1 vccd1 _22971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21922_ _21922_/A _21922_/B vssd1 vssd1 vccd1 vccd1 _21922_/Y sky130_fd_sc_hd__nand2_1
XFILLER_228_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21853_ _21876_/A _21853_/B vssd1 vssd1 vccd1 vccd1 _21854_/B sky130_fd_sc_hd__nor2_2
XFILLER_70_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20804_ _20804_/A vssd1 vssd1 vccd1 vccd1 _23756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21784_ _23828_/Q _23762_/Q vssd1 vssd1 vccd1 vccd1 _21786_/A sky130_fd_sc_hd__and2_1
XFILLER_212_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23523_ _23902_/CLK _23523_/D vssd1 vssd1 vccd1 vccd1 _23523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20735_ _13165_/Y _20732_/X _20734_/Y vssd1 vssd1 vccd1 vccd1 _20736_/C sky130_fd_sc_hd__a21oi_2
XFILLER_243_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_357_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23454_ _23550_/CLK _23454_/D vssd1 vssd1 vccd1 vccd1 _23454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20666_ _23731_/Q _20628_/X _20665_/X _20637_/X vssd1 vssd1 vccd1 vccd1 _23731_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_338_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22405_ _23573_/CLK _22405_/D vssd1 vssd1 vccd1 vccd1 _22405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23385_ _23545_/CLK _23385_/D vssd1 vssd1 vccd1 vccd1 _23385_/Q sky130_fd_sc_hd__dfxtp_1
X_20597_ _20597_/A _20631_/B vssd1 vssd1 vccd1 vccd1 _20601_/B sky130_fd_sc_hd__nor2_2
XFILLER_167_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_326_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22336_ _23440_/CLK _22336_/D vssd1 vssd1 vccd1 vccd1 _22336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_352_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_313_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_341_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22267_ _23466_/CLK _22267_/D vssd1 vssd1 vccd1 vccd1 _22267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12020_ _12020_/A vssd1 vssd1 vccd1 vccd1 _12717_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21218_ _21281_/A vssd1 vssd1 vccd1 vccd1 _21218_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22198_ _21398_/X _22195_/X _22196_/Y _22197_/Y _21677_/X vssd1 vssd1 vccd1 vccd1
+ _22198_/X sky130_fd_sc_hd__a311o_2
XFILLER_132_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_333_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21149_ _21149_/A _21177_/B vssd1 vssd1 vccd1 vccd1 _21149_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13971_ _13971_/A vssd1 vssd1 vccd1 vccd1 _13971_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15710_ _19223_/A vssd1 vssd1 vccd1 vccd1 _15710_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12922_ _22474_/Q _22634_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12922_/X sky130_fd_sc_hd__mux2_1
X_16690_ _22519_/Q _16679_/A vssd1 vssd1 vccd1 vccd1 _16806_/B sky130_fd_sc_hd__or2b_1
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15641_ _14839_/X _15489_/X _15637_/X _15640_/Y vssd1 vssd1 vccd1 vccd1 _15641_/X
+ sky130_fd_sc_hd__o211a_2
X_12853_ _12904_/A _12850_/X _12852_/X _12797_/X vssd1 vssd1 vccd1 vccd1 _12853_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_261_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _18360_/A _18366_/C vssd1 vssd1 vccd1 vccd1 _18360_/Y sky130_fd_sc_hd__nor2_1
X_11804_ _12318_/A vssd1 vssd1 vccd1 vccd1 _12097_/A sky130_fd_sc_hd__buf_2
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15572_ _15570_/X _22276_/Q _15750_/S vssd1 vssd1 vccd1 vccd1 _15573_/A sky130_fd_sc_hd__mux2_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _12784_/A _12784_/B vssd1 vssd1 vccd1 vccd1 _12784_/Y sky130_fd_sc_hd__nor2_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _17245_/A _17310_/X _16996_/A _17283_/X vssd1 vssd1 vccd1 vccd1 _17311_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_202_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _23911_/Q vssd1 vssd1 vccd1 vccd1 _21300_/B sky130_fd_sc_hd__buf_4
XFILLER_348_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18291_ _22923_/Q _18287_/C _18290_/Y vssd1 vssd1 vccd1 vccd1 _22923_/D sky130_fd_sc_hd__o21a_1
X_11735_ _23312_/Q _23280_/Q _23248_/Q _23536_/Q _11457_/C _12020_/A vssd1 vssd1 vccd1
+ vccd1 _11736_/B sky130_fd_sc_hd__mux4_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17242_/A vssd1 vssd1 vccd1 vccd1 _17242_/X sky130_fd_sc_hd__buf_2
X_14454_ _15590_/A vssd1 vssd1 vccd1 vccd1 _14455_/A sky130_fd_sc_hd__buf_2
XFILLER_175_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11666_ _12909_/A _11666_/B vssd1 vssd1 vccd1 vccd1 _11666_/X sky130_fd_sc_hd__or2_1
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13405_ _13402_/A _13402_/B _13246_/Y vssd1 vssd1 vccd1 vccd1 _13406_/B sky130_fd_sc_hd__a21oi_1
XFILLER_317_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17173_ _17171_/X _17172_/Y _17163_/B vssd1 vssd1 vccd1 vccd1 _17173_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_127_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14385_ _14385_/A _14385_/B vssd1 vssd1 vccd1 vccd1 _15346_/B sky130_fd_sc_hd__or2_1
X_11597_ _22794_/Q _22762_/Q _22663_/Q _22730_/Q _12755_/A _11568_/A vssd1 vssd1 vccd1
+ vccd1 _11597_/X sky130_fd_sc_hd__mux4_1
XFILLER_316_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16124_ _19258_/A vssd1 vssd1 vccd1 vccd1 _16124_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13336_ _13371_/B _13371_/C _13371_/A vssd1 vssd1 vccd1 vccd1 _13375_/A sky130_fd_sc_hd__a21oi_4
XFILLER_316_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_304_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16055_ _16054_/A _14793_/A _16054_/Y _15583_/A vssd1 vssd1 vccd1 vccd1 _16055_/X
+ sky130_fd_sc_hd__o211a_1
X_13267_ _22289_/Q _23105_/Q _23521_/Q _22450_/Q _11206_/X _11208_/X vssd1 vssd1 vccd1
+ vccd1 _13268_/B sky130_fd_sc_hd__mux4_1
XFILLER_332_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15006_ _14385_/B _14371_/Y _14175_/Y vssd1 vssd1 vccd1 vccd1 _15918_/S sky130_fd_sc_hd__o21ai_4
XFILLER_29_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12218_ _11330_/A _12217_/X _11346_/A vssd1 vssd1 vccd1 vccd1 _12218_/X sky130_fd_sc_hd__o21a_1
XFILLER_130_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_307_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13198_ _23229_/Q _23197_/Q _23165_/Q _23133_/Q _13090_/S _13195_/X vssd1 vssd1 vccd1
+ vccd1 _13199_/B sky130_fd_sc_hd__mux4_2
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19814_ _19814_/A vssd1 vssd1 vccd1 vccd1 _23543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_285_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_297_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12149_ _22369_/Q _22401_/Q _22690_/Q _23057_/Q _11741_/X _12025_/A vssd1 vssd1 vccd1
+ vccd1 _12149_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19745_ _19756_/A vssd1 vssd1 vccd1 vccd1 _19754_/S sky130_fd_sc_hd__buf_2
X_16957_ _23461_/Q _17230_/A _17231_/A _17042_/A _14520_/B vssd1 vssd1 vccd1 vccd1
+ _16957_/X sky130_fd_sc_hd__a32o_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15908_ _23773_/Q _14911_/A _14913_/A _15906_/X _15907_/X vssd1 vssd1 vccd1 vccd1
+ _15908_/X sky130_fd_sc_hd__a221o_1
XFILLER_323_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19676_ _19233_/X _23482_/Q _19682_/S vssd1 vssd1 vccd1 vccd1 _19677_/A sky130_fd_sc_hd__mux2_1
XFILLER_253_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16888_ _16888_/A vssd1 vssd1 vccd1 vccd1 _22543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_292_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18627_ _18695_/S vssd1 vssd1 vccd1 vccd1 _18636_/S sky130_fd_sc_hd__buf_8
XFILLER_225_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15839_ _23803_/Q _14917_/X _15067_/X vssd1 vssd1 vccd1 vccd1 _15839_/X sky130_fd_sc_hd__a21o_1
XFILLER_227_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18558_ _16819_/X _23014_/Q _18564_/S vssd1 vssd1 vccd1 vccd1 _18559_/A sky130_fd_sc_hd__mux2_1
XFILLER_252_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_307_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17509_ _17509_/A vssd1 vssd1 vccd1 vccd1 _22661_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18489_ _20067_/A vssd1 vssd1 vccd1 vccd1 _18516_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20520_ _20520_/A _20520_/B _20520_/C _20520_/D vssd1 vssd1 vccd1 vccd1 _20526_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_220_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_348_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_59_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23542_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20451_ _23699_/Q _20468_/B vssd1 vssd1 vccd1 vccd1 _20451_/X sky130_fd_sc_hd__or2_1
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_335_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_323_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23170_ _23489_/CLK _23170_/D vssd1 vssd1 vccd1 vccd1 _23170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20382_ _17289_/A _20261_/X _20383_/B vssd1 vssd1 vccd1 vccd1 _20382_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_334_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_335_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22121_ _21307_/X _22105_/X _22112_/X _22120_/X _21410_/X vssd1 vssd1 vccd1 vccd1
+ _22121_/Y sky130_fd_sc_hd__o2111ai_2
XTAP_7209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22052_ _22052_/A _22052_/B vssd1 vssd1 vccd1 vccd1 _22155_/A sky130_fd_sc_hd__and2_1
XTAP_6519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_314_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21003_ _20579_/A _20988_/X _21002_/X _20997_/X vssd1 vssd1 vccd1 vccd1 _23816_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_276_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_303_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22954_ _23599_/CLK _22954_/D vssd1 vssd1 vccd1 vccd1 _22954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21905_ _21936_/C _21937_/A vssd1 vssd1 vccd1 vccd1 _21933_/B sky130_fd_sc_hd__nand2_1
X_22885_ _23584_/CLK _22885_/D vssd1 vssd1 vccd1 vccd1 _22885_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_71_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21836_ _21836_/A _21836_/B vssd1 vssd1 vccd1 vccd1 _21837_/B sky130_fd_sc_hd__nor2_1
XPHY_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21767_ _21767_/A vssd1 vssd1 vccd1 vccd1 _21767_/X sky130_fd_sc_hd__buf_2
XPHY_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11520_ _22290_/Q _23106_/Q _23522_/Q _22451_/Q _11517_/X _11519_/X vssd1 vssd1 vccd1
+ vccd1 _11521_/B sky130_fd_sc_hd__mux4_1
XFILLER_212_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23506_ _23538_/CLK _23506_/D vssd1 vssd1 vccd1 vccd1 _23506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_346_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20718_ _21165_/A _20744_/B vssd1 vssd1 vccd1 vccd1 _20721_/B sky130_fd_sc_hd__nor2_4
XFILLER_157_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21698_ _23793_/Q _21683_/X _21697_/Y _21346_/X vssd1 vssd1 vccd1 vccd1 _21699_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11451_ _13718_/A _11451_/B _11451_/C vssd1 vssd1 vccd1 vccd1 _11452_/B sky130_fd_sc_hd__and3_2
X_23437_ _23565_/CLK _23437_/D vssd1 vssd1 vccd1 vccd1 _23437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20649_ _20733_/A vssd1 vssd1 vccd1 vccd1 _20649_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_354_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14170_ _15066_/B vssd1 vssd1 vccd1 vccd1 _14745_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_301_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23368_ _23368_/CLK _23368_/D vssd1 vssd1 vccd1 vccd1 _23368_/Q sky130_fd_sc_hd__dfxtp_1
X_11382_ _14172_/C _11382_/B _11382_/C vssd1 vssd1 vccd1 vccd1 _12520_/S sky130_fd_sc_hd__nand3_4
XFILLER_152_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_341_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13121_ _13121_/A _13121_/B vssd1 vssd1 vccd1 vccd1 _13121_/Y sky130_fd_sc_hd__nor2_1
XFILLER_194_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22319_ _23582_/CLK _22319_/D vssd1 vssd1 vccd1 vccd1 _22319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_341_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23299_ _23491_/CLK _23299_/D vssd1 vssd1 vccd1 vccd1 _23299_/Q sky130_fd_sc_hd__dfxtp_1
X_13052_ _23488_/Q _23584_/Q _22548_/Q _22352_/Q _13088_/S _13037_/X vssd1 vssd1 vccd1
+ vccd1 _13052_/X sky130_fd_sc_hd__mux4_1
XFILLER_313_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12003_ _13616_/A _21773_/A _12739_/A vssd1 vssd1 vccd1 vccd1 _12170_/A sky130_fd_sc_hd__mux2_2
XFILLER_78_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17860_ _17860_/A vssd1 vssd1 vccd1 vccd1 _22801_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_289_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_289_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16811_ _13457_/A _13934_/A _16810_/B _16808_/D _16810_/Y vssd1 vssd1 vccd1 vccd1
+ _16811_/X sky130_fd_sc_hd__a221o_1
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17791_ _17791_/A vssd1 vssd1 vccd1 vccd1 _22770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_293_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19530_ _19229_/X _23417_/Q _19538_/S vssd1 vssd1 vccd1 vccd1 _19531_/A sky130_fd_sc_hd__mux2_1
X_16742_ _16742_/A vssd1 vssd1 vccd1 vccd1 _22500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13954_ _16679_/B vssd1 vssd1 vccd1 vccd1 _13965_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_219_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_253_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12905_ _23482_/Q _23578_/Q _22542_/Q _22346_/Q _12776_/X _12777_/X vssd1 vssd1 vccd1
+ vccd1 _12906_/B sky130_fd_sc_hd__mux4_1
XFILLER_74_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19461_ _19461_/A vssd1 vssd1 vccd1 vccd1 _23386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16673_ _22483_/Q _16300_/X _16673_/S vssd1 vssd1 vccd1 vccd1 _16674_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13885_ _14216_/A _13479_/X _13832_/A _14071_/A vssd1 vssd1 vccd1 vccd1 _15119_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_234_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18412_ _22965_/Q _18412_/B vssd1 vssd1 vccd1 vccd1 _18418_/C sky130_fd_sc_hd__and2_1
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15624_ _18824_/A vssd1 vssd1 vccd1 vccd1 _19217_/A sky130_fd_sc_hd__clkbuf_2
X_12836_ _12836_/A _12836_/B vssd1 vssd1 vccd1 vccd1 _12836_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ _23356_/Q _18846_/X _19394_/S vssd1 vssd1 vccd1 vccd1 _19393_/A sky130_fd_sc_hd__mux2_1
XFILLER_262_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18343_ _22941_/Q _18343_/B vssd1 vssd1 vccd1 vccd1 _18349_/C sky130_fd_sc_hd__and2_1
X_15555_ _23700_/Q _15210_/A _15554_/X vssd1 vssd1 vccd1 vccd1 _15555_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _12985_/A _12766_/X _11132_/A vssd1 vssd1 vccd1 vccd1 _12767_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_187_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_349_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14506_ _14510_/A _14506_/B vssd1 vssd1 vccd1 vccd1 _14931_/A sky130_fd_sc_hd__or2_2
XFILLER_202_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_337_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18274_ _18275_/A _18275_/C _22919_/Q vssd1 vssd1 vccd1 vccd1 _18276_/B sky130_fd_sc_hd__a21oi_1
X_11718_ _11723_/A _11718_/B vssd1 vssd1 vccd1 vccd1 _11718_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15486_ _13833_/A _15484_/Y _15830_/B _13737_/A vssd1 vssd1 vccd1 vccd1 _15486_/Y
+ sky130_fd_sc_hd__a22oi_1
X_12698_ _12698_/A vssd1 vssd1 vccd1 vccd1 _12919_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_348_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17225_ _17169_/A _17223_/Y _17224_/Y _17283_/A vssd1 vssd1 vccd1 vccd1 _18449_/B
+ sky130_fd_sc_hd__a31o_4
X_14437_ _14609_/A _20890_/A vssd1 vssd1 vccd1 vccd1 _15068_/C sky130_fd_sc_hd__or2_4
XFILLER_30_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11649_ _12476_/A vssd1 vssd1 vccd1 vccd1 _12216_/A sky130_fd_sc_hd__buf_4
Xinput11 core_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_2
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 core_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_2
XFILLER_329_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput33 core_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_1
X_17156_ input85/X input50/X _17219_/S vssd1 vssd1 vccd1 vccd1 _17156_/X sky130_fd_sc_hd__mux2_8
Xinput44 dout0[10] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_2
X_14368_ _14368_/A vssd1 vssd1 vccd1 vccd1 _15387_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xinput55 dout0[20] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_2
XFILLER_155_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput66 dout0[30] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__buf_2
Xinput77 dout0[40] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16107_ _23714_/Q _15592_/X _16106_/X vssd1 vssd1 vccd1 vccd1 _16107_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_128_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_305_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput88 dout0[50] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13319_ _13319_/A _13319_/B vssd1 vssd1 vccd1 vccd1 _13319_/X sky130_fd_sc_hd__or2_1
Xinput99 dout0[60] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__clkbuf_1
X_17087_ _13945_/B _17086_/X _17087_/S vssd1 vssd1 vccd1 vccd1 _17087_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14299_ _14297_/X _14298_/X _14310_/S vssd1 vssd1 vccd1 vccd1 _14299_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16038_ _14570_/X _21274_/A _16037_/X _15365_/X vssd1 vssd1 vccd1 vccd1 _16038_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_192_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_297_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_177_wb_clk_i _23917_/CLK vssd1 vssd1 vccd1 vccd1 _23915_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_285_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_300_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_106_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23582_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_285_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17989_ _22839_/Q _17981_/X _17988_/X _17979_/X vssd1 vssd1 vccd1 vccd1 _22839_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_300_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19728_ _19204_/X _23505_/Q _19732_/S vssd1 vssd1 vccd1 vccd1 _19729_/A sky130_fd_sc_hd__mux2_1
XFILLER_270_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19659_ _19659_/A vssd1 vssd1 vccd1 vccd1 _23474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22670_ _23581_/CLK _22670_/D vssd1 vssd1 vccd1 vccd1 _22670_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_280_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21621_ _14180_/B _21605_/B _21618_/Y _21619_/X vssd1 vssd1 vccd1 vccd1 _21689_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_179_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21552_ _21716_/B vssd1 vssd1 vccd1 vccd1 _21841_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_178_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20503_ _21555_/A _22046_/A vssd1 vssd1 vccd1 vccd1 _21549_/A sky130_fd_sc_hd__nand2_4
XFILLER_339_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21483_ _20217_/A _21868_/A _21441_/A _21500_/A vssd1 vssd1 vccd1 vccd1 _21526_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23222_ _23573_/CLK _23222_/D vssd1 vssd1 vccd1 vccd1 _23222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20434_ _23692_/Q _20413_/X _20432_/Y _20433_/X vssd1 vssd1 vccd1 vccd1 _23692_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_335_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23153_ _23537_/CLK _23153_/D vssd1 vssd1 vccd1 vccd1 _23153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20365_ _20302_/X _20363_/Y _20364_/X _22116_/B _20307_/X vssd1 vssd1 vccd1 vccd1
+ _20731_/A sky130_fd_sc_hd__a32o_4
XTAP_7017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22104_ _22155_/C _22104_/B vssd1 vssd1 vccd1 vccd1 _22104_/Y sky130_fd_sc_hd__xnor2_2
XTAP_7039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23084_ _23500_/CLK _23084_/D vssd1 vssd1 vccd1 vccd1 _23084_/Q sky130_fd_sc_hd__dfxtp_1
X_20296_ _20296_/A _20394_/B vssd1 vssd1 vccd1 vccd1 _20296_/Y sky130_fd_sc_hd__nand2_1
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_310_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_288_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22035_ _13960_/X _22018_/X _22026_/X _22034_/Y vssd1 vssd1 vccd1 vccd1 _22035_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_6349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_314_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22937_ _23649_/CLK _22937_/D vssd1 vssd1 vccd1 vccd1 _22937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13670_ _13670_/A _13670_/B _13670_/C _14147_/B vssd1 vssd1 vccd1 vccd1 _16534_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_204_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22868_ _23632_/CLK _22868_/D vssd1 vssd1 vccd1 vccd1 _22868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12621_ _12958_/A _12621_/B vssd1 vssd1 vccd1 vccd1 _12621_/Y sky130_fd_sc_hd__nor2_1
XFILLER_232_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21819_ _21819_/A _21819_/B vssd1 vssd1 vccd1 vccd1 _21821_/A sky130_fd_sc_hd__nand2_1
XFILLER_358_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22799_ _22801_/CLK _22799_/D vssd1 vssd1 vccd1 vccd1 _22799_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15340_ _15340_/A vssd1 vssd1 vccd1 vccd1 _15340_/Y sky130_fd_sc_hd__inv_2
XPHY_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12552_ _22781_/Q _22749_/Q _22650_/Q _22717_/Q _12245_/S _12292_/X vssd1 vssd1 vccd1
+ vccd1 _12553_/B sky130_fd_sc_hd__mux4_1
XFILLER_358_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_346_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ _23426_/Q _23042_/Q _23394_/Q _23362_/Q _13255_/S _11418_/A vssd1 vssd1 vccd1
+ vccd1 _11503_/X sky130_fd_sc_hd__mux4_1
XPHY_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15271_ _14431_/X _15259_/X _15269_/X _15270_/X _14937_/X vssd1 vssd1 vccd1 vccd1
+ _15271_/X sky130_fd_sc_hd__o32a_4
XFILLER_345_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12483_ _12474_/X _12478_/X _12480_/X _12482_/X _23898_/Q vssd1 vssd1 vccd1 vccd1
+ _12493_/B sky130_fd_sc_hd__a221o_1
XFILLER_327_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17010_ _17174_/B _17009_/X _16951_/A vssd1 vssd1 vccd1 vccd1 _17010_/X sky130_fd_sc_hd__o21a_1
XFILLER_345_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14222_ _14246_/B vssd1 vssd1 vccd1 vccd1 _14238_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11434_ _13037_/A vssd1 vssd1 vccd1 vccd1 _11435_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_314_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14153_ _14159_/A vssd1 vssd1 vccd1 vccd1 _14153_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11365_ _11365_/A vssd1 vssd1 vccd1 vccd1 _11365_/X sky130_fd_sc_hd__buf_4
XFILLER_314_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_4_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23467_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13104_ _23487_/Q _23583_/Q _22547_/Q _22351_/Q _11205_/A _13085_/X vssd1 vssd1 vccd1
+ vccd1 _13104_/X sky130_fd_sc_hd__mux4_2
XFILLER_302_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14084_ _22589_/Q _14081_/X _14082_/Y _14083_/X vssd1 vssd1 vccd1 vccd1 _14084_/X
+ sky130_fd_sc_hd__a22o_4
X_18961_ _18961_/A vssd1 vssd1 vccd1 vccd1 _23178_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11296_ _12784_/A vssd1 vssd1 vccd1 vccd1 _11515_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_180_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_313_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17912_ _22254_/A vssd1 vssd1 vccd1 vccd1 _17912_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13035_ _11435_/A _13034_/X _13158_/A vssd1 vssd1 vccd1 vccd1 _13035_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18892_ _23148_/Q _18795_/X _18896_/S vssd1 vssd1 vccd1 vccd1 _18893_/A sky130_fd_sc_hd__mux2_1
XTAP_6850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17843_ _17843_/A vssd1 vssd1 vccd1 vccd1 _22793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_310_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17774_ _22763_/Q _17604_/X _17776_/S vssd1 vssd1 vccd1 vccd1 _17775_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14986_ _14986_/A vssd1 vssd1 vccd1 vccd1 _22265_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_281_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19513_ _19513_/A vssd1 vssd1 vccd1 vccd1 _23409_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16725_ _16804_/A vssd1 vssd1 vccd1 vccd1 _16741_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_263_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13937_ _23919_/Q vssd1 vssd1 vccd1 vccd1 _21570_/A sky130_fd_sc_hd__buf_4
XFILLER_93_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_501 _15033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19444_ _23379_/Q _18817_/X _19444_/S vssd1 vssd1 vccd1 vccd1 _19445_/A sky130_fd_sc_hd__mux2_1
XFILLER_234_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_512 _17156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16656_ _22475_/Q _16275_/X _16662_/S vssd1 vssd1 vccd1 vccd1 _16657_/A sky130_fd_sc_hd__mux2_1
X_13868_ _13969_/A vssd1 vssd1 vccd1 vccd1 _13967_/B sky130_fd_sc_hd__clkbuf_4
XINSDIODE2_523 _14063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_534 _23944_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_545 _21186_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_343_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12819_ _22316_/Q _23452_/Q _12819_/S vssd1 vssd1 vccd1 vccd1 _12819_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_556 _23469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15607_ _15345_/A _15586_/X _15606_/Y _15697_/A vssd1 vssd1 vccd1 vccd1 _15607_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_349_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19375_ _23348_/Q _18820_/X _19383_/S vssd1 vssd1 vccd1 vccd1 _19376_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_320_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16587_ _16587_/A vssd1 vssd1 vccd1 vccd1 _22444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13799_ _14241_/A _13711_/B _13798_/Y _15830_/A vssd1 vssd1 vccd1 vccd1 _13799_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18326_ _22935_/Q _18326_/B vssd1 vssd1 vccd1 vccd1 _18332_/C sky130_fd_sc_hd__and2_1
XFILLER_176_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ _15538_/A _15538_/B vssd1 vssd1 vccd1 vccd1 _15538_/Y sky130_fd_sc_hd__nor2_1
XFILLER_175_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18257_ _18263_/A _18263_/B _18175_/X vssd1 vssd1 vccd1 vccd1 _18257_/Y sky130_fd_sc_hd__a21oi_1
X_15469_ _14807_/A _15453_/A _15574_/A vssd1 vssd1 vccd1 vccd1 _15469_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_329_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17208_ _22573_/Q _17199_/X _17190_/X _17207_/X vssd1 vssd1 vccd1 vccd1 _22573_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_318_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18188_ _18188_/A _18188_/B _18178_/B vssd1 vssd1 vccd1 vccd1 _18195_/C sky130_fd_sc_hd__or3b_1
XFILLER_129_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17139_ _17070_/A _17132_/X _17138_/X _17109_/X vssd1 vssd1 vccd1 vccd1 _17139_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_144_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_289_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20150_ _20205_/A _20532_/D vssd1 vssd1 vccd1 vccd1 _20216_/A sky130_fd_sc_hd__or2_1
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_289_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20081_ _23635_/Q vssd1 vssd1 vccd1 vccd1 _20090_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_301_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23840_ _23876_/CLK _23840_/D vssd1 vssd1 vccd1 vccd1 _23840_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_111_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23771_ _23776_/CLK _23771_/D vssd1 vssd1 vccd1 vccd1 _23771_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20983_ _23811_/Q _20925_/A _20982_/X _20978_/X vssd1 vssd1 vccd1 vccd1 _23811_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22722_ _23054_/CLK _22722_/D vssd1 vssd1 vccd1 vccd1 _22722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_74_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23545_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_213_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22653_ _23144_/CLK _22653_/D vssd1 vssd1 vccd1 vccd1 _22653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21604_ _21604_/A _21624_/A vssd1 vssd1 vccd1 vccd1 _21690_/B sky130_fd_sc_hd__nor2_2
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22584_ _23649_/CLK _22584_/D vssd1 vssd1 vccd1 vccd1 _22584_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_194_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_327_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21535_ _21535_/A _21535_/B vssd1 vssd1 vccd1 vccd1 _21535_/X sky130_fd_sc_hd__xor2_1
XFILLER_223_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21466_ _21466_/A vssd1 vssd1 vccd1 vccd1 _22171_/B sky130_fd_sc_hd__buf_2
XFILLER_336_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23205_ _23493_/CLK _23205_/D vssd1 vssd1 vccd1 vccd1 _23205_/Q sky130_fd_sc_hd__dfxtp_1
X_20417_ _23686_/Q _20413_/X _20416_/Y _20392_/X vssd1 vssd1 vccd1 vccd1 _23686_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_162_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21397_ _21575_/A vssd1 vssd1 vccd1 vccd1 _21676_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_135_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23136_ _23264_/CLK _23136_/D vssd1 vssd1 vccd1 vccd1 _23136_/Q sky130_fd_sc_hd__dfxtp_1
X_11150_ _11708_/S vssd1 vssd1 vccd1 vccd1 _11151_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20348_ _17232_/A _20215_/X _20347_/X vssd1 vssd1 vccd1 vccd1 _20348_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_350_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_311_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_325_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23067_ _23581_/CLK _23067_/D vssd1 vssd1 vccd1 vccd1 _23067_/Q sky130_fd_sc_hd__dfxtp_1
X_11081_ _23892_/Q vssd1 vssd1 vccd1 vccd1 _13421_/A sky130_fd_sc_hd__buf_2
XTAP_6146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20279_ _20279_/A _20279_/B vssd1 vssd1 vccd1 vccd1 _20279_/Y sky130_fd_sc_hd__nand2_1
XFILLER_295_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput201 localMemory_wb_adr_i[1] vssd1 vssd1 vccd1 vccd1 input201/X sky130_fd_sc_hd__clkbuf_1
XFILLER_299_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput212 localMemory_wb_adr_i[8] vssd1 vssd1 vccd1 vccd1 input212/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22018_ _21613_/X _22017_/Y _21560_/X _23804_/Q vssd1 vssd1 vccd1 vccd1 _22018_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput223 localMemory_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input223/X sky130_fd_sc_hd__buf_6
XTAP_6179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput234 localMemory_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 input234/X sky130_fd_sc_hd__buf_8
XTAP_5445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 localMemory_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input245/X sky130_fd_sc_hd__buf_6
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput256 manufacturerID[2] vssd1 vssd1 vccd1 vccd1 input256/X sky130_fd_sc_hd__clkbuf_4
XFILLER_291_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput267 partID[12] vssd1 vssd1 vccd1 vccd1 input267/X sky130_fd_sc_hd__clkbuf_1
XTAP_5478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ _14661_/X _14663_/X _14840_/S vssd1 vssd1 vccd1 vccd1 _14840_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput278 partID[8] vssd1 vssd1 vccd1 vccd1 input278/X sky130_fd_sc_hd__clkbuf_1
XTAP_5489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ _15798_/A vssd1 vssd1 vccd1 vccd1 _14839_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11983_ _22276_/Q _23092_/Q _23508_/Q _22437_/Q _11637_/X _12793_/A vssd1 vssd1 vccd1
+ vccd1 _11984_/B sky130_fd_sc_hd__mux4_1
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16510_ _16510_/A vssd1 vssd1 vccd1 vccd1 _22411_/D sky130_fd_sc_hd__clkbuf_1
X_13722_ _13786_/A _13722_/B vssd1 vssd1 vccd1 vccd1 _13723_/A sky130_fd_sc_hd__and2_4
Xclkbuf_4_4_0_wb_clk_i INSDIODE2_358/DIODE vssd1 vssd1 vccd1 vccd1 _23931_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_95_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17490_ _22653_/Q _16230_/X _17494_/S vssd1 vssd1 vccd1 vccd1 _17491_/A sky130_fd_sc_hd__mux2_1
XFILLER_260_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16441_ _16441_/A vssd1 vssd1 vccd1 vccd1 _22381_/D sky130_fd_sc_hd__clkbuf_1
X_13653_ _17385_/B _14224_/B vssd1 vssd1 vccd1 vccd1 _13653_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12604_ _13913_/A _13356_/A _13355_/A _12603_/X vssd1 vssd1 vccd1 vccd1 _13354_/B
+ sky130_fd_sc_hd__o31ai_2
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16372_ _16372_/A vssd1 vssd1 vccd1 vccd1 _22351_/D sky130_fd_sc_hd__clkbuf_1
X_19160_ _19160_/A vssd1 vssd1 vccd1 vccd1 _23267_/D sky130_fd_sc_hd__clkbuf_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ _13686_/A _13686_/B _13985_/A _13584_/D vssd1 vssd1 vccd1 vccd1 _14224_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_358_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_346_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _22875_/Q _17956_/A _18053_/A _23008_/Q _18054_/A vssd1 vssd1 vccd1 vccd1
+ _18111_/X sky130_fd_sc_hd__a221o_1
X_15323_ _18804_/A vssd1 vssd1 vccd1 vccd1 _19197_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _22454_/Q _22614_/Q _12535_/S vssd1 vssd1 vccd1 vccd1 _12536_/B sky130_fd_sc_hd__mux2_1
X_19091_ _19091_/A _19771_/B vssd1 vssd1 vccd1 vccd1 _19148_/A sky130_fd_sc_hd__nor2_8
XFILLER_346_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18042_ _22852_/Q _18035_/X _18041_/X _18029_/X vssd1 vssd1 vccd1 vccd1 _22852_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15254_ _14671_/S _15252_/Y _15253_/X vssd1 vssd1 vccd1 vccd1 _15850_/B sky130_fd_sc_hd__a21o_1
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12466_ _11127_/A _12463_/Y _12465_/Y _11240_/A vssd1 vssd1 vccd1 vccd1 _12466_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_346_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_315_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14205_ _17385_/B _19969_/B vssd1 vssd1 vccd1 vccd1 _14207_/B sky130_fd_sc_hd__or2b_4
X_11417_ _12368_/B vssd1 vssd1 vccd1 vccd1 _13718_/A sky130_fd_sc_hd__buf_6
XFILLER_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_299_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15185_ _15485_/B vssd1 vssd1 vccd1 vccd1 _15433_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_342_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12397_ _12397_/A _12397_/B vssd1 vssd1 vccd1 vccd1 _12397_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_315_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14136_ _23012_/Q _14700_/C vssd1 vssd1 vccd1 vccd1 _14137_/A sky130_fd_sc_hd__and2_4
XFILLER_181_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11348_ _11348_/A vssd1 vssd1 vccd1 vccd1 _12797_/A sky130_fd_sc_hd__buf_4
XFILLER_152_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19993_ _23610_/Q _19994_/C _19992_/Y vssd1 vssd1 vccd1 vccd1 _23610_/D sky130_fd_sc_hd__o21a_1
XFILLER_99_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14067_ input236/X _14058_/X _14066_/X vssd1 vssd1 vccd1 vccd1 _14067_/X sky130_fd_sc_hd__a21bo_4
X_18944_ _23172_/Q _18871_/X _18944_/S vssd1 vssd1 vccd1 vccd1 _18945_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11279_ _23897_/Q vssd1 vssd1 vccd1 vccd1 _11280_/A sky130_fd_sc_hd__inv_2
XTAP_7381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13018_ _13592_/A _13605_/A _13322_/C _13018_/D vssd1 vssd1 vccd1 vccd1 _13018_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_315_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18875_ _18931_/A vssd1 vssd1 vccd1 vccd1 _18944_/S sky130_fd_sc_hd__buf_6
XFILLER_140_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17826_ _22786_/Q _17575_/X _17826_/S vssd1 vssd1 vccd1 vccd1 _17827_/A sky130_fd_sc_hd__mux2_1
XFILLER_251_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_294_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17757_ _22755_/Q _17578_/X _17765_/S vssd1 vssd1 vccd1 vccd1 _17758_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14969_ _14218_/X _15380_/A _15381_/A _13789_/A _14968_/Y vssd1 vssd1 vccd1 vccd1
+ _14969_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_242_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16708_ _22491_/Q _16689_/X _16693_/X input36/X vssd1 vssd1 vccd1 vccd1 _16709_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_208_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17688_ _17688_/A vssd1 vssd1 vccd1 vccd1 _22724_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_320 _16107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_331 _17001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_342 _17139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19427_ _23371_/Q _18792_/X _19433_/S vssd1 vssd1 vccd1 vccd1 _19428_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_353 _17238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16639_ _16639_/A vssd1 vssd1 vccd1 vccd1 _22467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_364 _23703_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_375 _23468_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_356_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_386 _18009_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19358_ _19358_/A vssd1 vssd1 vccd1 vccd1 _23340_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_397 _14090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_349_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18309_ _18317_/A _18314_/C vssd1 vssd1 vccd1 vccd1 _18309_/Y sky130_fd_sc_hd__nor2_1
XFILLER_337_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19289_ _19194_/X _23310_/Q _19289_/S vssd1 vssd1 vccd1 vccd1 _19290_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21320_ _21320_/A _21320_/B vssd1 vssd1 vccd1 vccd1 _21321_/A sky130_fd_sc_hd__nor2_8
XFILLER_176_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_192_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23494_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21251_ _21251_/A vssd1 vssd1 vccd1 vccd1 _23896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_289_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20202_ _23657_/Q _20223_/B vssd1 vssd1 vccd1 vccd1 _20202_/X sky130_fd_sc_hd__or2_1
XFILLER_150_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_121_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23637_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21182_ _20754_/A _21158_/X _21142_/A _20515_/A _21161_/X vssd1 vssd1 vccd1 vccd1
+ _21182_/X sky130_fd_sc_hd__a221o_1
XFILLER_104_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_320_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20133_ _23651_/Q _20136_/C vssd1 vssd1 vccd1 vccd1 _20134_/B sky130_fd_sc_hd__xnor2_1
XFILLER_131_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20064_ _20086_/A _20064_/B _20079_/C vssd1 vssd1 vccd1 vccd1 _23630_/D sky130_fd_sc_hd__nor3_1
XFILLER_286_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_13 _22122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_24 _17682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_35 _19029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_46 _21357_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_57 _21023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_68 _21831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23823_ _23824_/CLK _23823_/D vssd1 vssd1 vccd1 vccd1 _23823_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_261_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_79 _21848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23754_ _23755_/CLK _23754_/D vssd1 vssd1 vccd1 vccd1 _23754_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20966_ _20966_/A vssd1 vssd1 vccd1 vccd1 _20966_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22705_ _23584_/CLK _22705_/D vssd1 vssd1 vccd1 vccd1 _22705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_340_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23685_ _23696_/CLK _23685_/D vssd1 vssd1 vccd1 vccd1 _23685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20897_ _20926_/A vssd1 vssd1 vccd1 vccd1 _20897_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22636_ _23577_/CLK _22636_/D vssd1 vssd1 vccd1 vccd1 _22636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_328_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22567_ _22600_/CLK _22567_/D vssd1 vssd1 vccd1 vccd1 _22567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_328_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ _22459_/Q _22619_/Q _22298_/Q _23434_/Q _11920_/A _11815_/A vssd1 vssd1 vccd1
+ vccd1 _12321_/B sky130_fd_sc_hd__mux4_1
XFILLER_182_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21518_ _21518_/A vssd1 vssd1 vccd1 vccd1 _21518_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22498_ _23704_/CLK _22498_/D vssd1 vssd1 vccd1 vccd1 _22498_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_355_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_336_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ _23307_/Q _23275_/Q _23243_/Q _23531_/Q _11414_/A _11703_/A vssd1 vssd1 vccd1
+ vccd1 _12252_/B sky130_fd_sc_hd__mux4_1
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21449_ _21485_/A _21485_/B vssd1 vssd1 vccd1 vccd1 _21451_/A sky130_fd_sc_hd__and2_1
XFILLER_79_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11202_ _14393_/A _11202_/B vssd1 vssd1 vccd1 vccd1 _11202_/Y sky130_fd_sc_hd__nand2_1
X_12182_ _22300_/Q _23436_/Q _12349_/S vssd1 vssd1 vccd1 vccd1 _12183_/B sky130_fd_sc_hd__mux2_1
XFILLER_351_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_311_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11133_ _11133_/A vssd1 vssd1 vccd1 vccd1 _11134_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_295_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23119_ _23535_/CLK _23119_/D vssd1 vssd1 vccd1 vccd1 _23119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_295_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16990_ _23462_/Q _16987_/X _16988_/X _16989_/X _14619_/X vssd1 vssd1 vccd1 vccd1
+ _16990_/X sky130_fd_sc_hd__a32o_1
XFILLER_352_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_296_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15941_ _16039_/C _15941_/B vssd1 vssd1 vccd1 vccd1 _15941_/X sky130_fd_sc_hd__or2_2
XFILLER_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18660_ _18682_/A vssd1 vssd1 vccd1 vccd1 _18669_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_95_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ _14866_/A _15867_/X _15871_/Y _14896_/A vssd1 vssd1 vccd1 vccd1 _15872_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_77_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17611_ _17627_/A vssd1 vssd1 vccd1 vccd1 _17624_/S sky130_fd_sc_hd__buf_2
X_14823_ input161/X input126/X _15030_/S vssd1 vssd1 vccd1 vccd1 _14823_/X sky130_fd_sc_hd__mux2_8
XFILLER_218_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18591_ _16867_/X _23029_/Q _18597_/S vssd1 vssd1 vccd1 vccd1 _18592_/A sky130_fd_sc_hd__mux2_1
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17542_ _22677_/Q _16306_/X _17542_/S vssd1 vssd1 vccd1 vccd1 _17543_/A sky130_fd_sc_hd__mux2_1
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11966_ _12056_/A _11964_/X _12687_/A vssd1 vssd1 vccd1 vccd1 _11966_/Y sky130_fd_sc_hd__o21ai_1
X_14754_ _22916_/Q _14752_/X _14753_/X _14729_/X vssd1 vssd1 vccd1 vccd1 _14754_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_251_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13705_ _15180_/A vssd1 vssd1 vccd1 vccd1 _13706_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17473_ _17529_/A vssd1 vssd1 vccd1 vccd1 _17542_/S sky130_fd_sc_hd__buf_6
X_14685_ _16131_/B vssd1 vssd1 vccd1 vccd1 _15256_/B sky130_fd_sc_hd__buf_2
XFILLER_260_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11897_ _22785_/Q _22753_/Q _22654_/Q _22721_/Q _11777_/S _11590_/A vssd1 vssd1 vccd1
+ vccd1 _11897_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19212_ _19212_/A vssd1 vssd1 vccd1 vccd1 _23283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_338_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16424_ _16424_/A vssd1 vssd1 vccd1 vccd1 _22373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13636_ _13974_/A _13966_/A _13636_/C _13636_/D vssd1 vssd1 vccd1 vccd1 _13636_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_32_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19143_ _19143_/A vssd1 vssd1 vccd1 vccd1 _23259_/D sky130_fd_sc_hd__clkbuf_1
X_16355_ _15749_/X _22344_/Q _16355_/S vssd1 vssd1 vccd1 vccd1 _16356_/A sky130_fd_sc_hd__mux2_1
X_13567_ _13581_/A _23939_/Q _13490_/A _13566_/Y vssd1 vssd1 vccd1 vccd1 _13583_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_358_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_301_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12518_ _12511_/X _12513_/X _12515_/X _12517_/X _11272_/A vssd1 vssd1 vccd1 vccd1
+ _12519_/C sky130_fd_sc_hd__a221o_1
X_15306_ _23823_/Q _15211_/X _15302_/X _15305_/X _15222_/X vssd1 vssd1 vccd1 vccd1
+ _15306_/X sky130_fd_sc_hd__a221o_2
X_19074_ _19074_/A vssd1 vssd1 vccd1 vccd1 _23229_/D sky130_fd_sc_hd__clkbuf_1
X_16286_ _16286_/A vssd1 vssd1 vccd1 vccd1 _22317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_346_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13498_ _12113_/B _13497_/Y _15460_/A vssd1 vssd1 vccd1 vccd1 _13499_/A sky130_fd_sc_hd__o21bai_1
XFILLER_185_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18025_ hold1/A _18016_/X _18024_/X _18000_/X vssd1 vssd1 vccd1 vccd1 _22846_/D sky130_fd_sc_hd__o211a_1
XFILLER_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12449_ _23900_/Q vssd1 vssd1 vccd1 vccd1 _12449_/X sky130_fd_sc_hd__clkbuf_4
X_15237_ _21591_/B vssd1 vssd1 vccd1 vccd1 _21576_/A sky130_fd_sc_hd__buf_6
XFILLER_299_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_303_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15168_ _19188_/A vssd1 vssd1 vccd1 vccd1 _15168_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14119_ _14119_/A _14119_/B _14119_/C _14119_/D vssd1 vssd1 vccd1 vccd1 _18009_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_299_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19976_ _23604_/Q _19976_/B _19976_/C vssd1 vssd1 vccd1 vccd1 _19977_/C sky130_fd_sc_hd__and3_1
X_15099_ _15367_/A _15099_/B vssd1 vssd1 vccd1 vccd1 _15099_/Y sky130_fd_sc_hd__nor2_1
XFILLER_330_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_286_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18927_ _23164_/Q _18846_/X _18929_/S vssd1 vssd1 vccd1 vccd1 _18928_/A sky130_fd_sc_hd__mux2_1
XFILLER_302_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18858_ _18858_/A vssd1 vssd1 vccd1 vccd1 _23135_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_269_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17809_ _22778_/Q _17550_/X _17815_/S vssd1 vssd1 vccd1 vccd1 _17810_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18789_ _18872_/S vssd1 vssd1 vccd1 vccd1 _18802_/S sky130_fd_sc_hd__buf_4
XFILLER_283_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20820_ _20820_/A vssd1 vssd1 vccd1 vccd1 _23760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20751_ _22166_/A _20632_/X _20750_/X vssd1 vssd1 vccd1 vccd1 _20752_/C sky130_fd_sc_hd__o21a_2
XFILLER_90_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_150 _20353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_161 _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_172 _17029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_183 _14059_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23470_ _23565_/CLK _23470_/D vssd1 vssd1 vccd1 vccd1 _23470_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_357_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_194 _13945_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20682_ _21846_/A _20648_/X _20681_/Y vssd1 vssd1 vccd1 vccd1 _20683_/C sky130_fd_sc_hd__a21oi_4
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22421_ _23851_/CLK _22421_/D vssd1 vssd1 vccd1 vccd1 _22421_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_195_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_287_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22352_ _23552_/CLK _22352_/D vssd1 vssd1 vccd1 vccd1 _22352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_276_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21303_ _21328_/A vssd1 vssd1 vccd1 vccd1 _21410_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22283_ _23453_/CLK _22283_/D vssd1 vssd1 vccd1 vccd1 _22283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_312_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21234_ _14535_/X _21229_/X _21233_/Y _21218_/X vssd1 vssd1 vccd1 vccd1 _23890_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21165_ _21165_/A _21177_/B vssd1 vssd1 vccd1 vccd1 _21165_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20116_ _23645_/Q _20119_/A _20115_/Y vssd1 vssd1 vccd1 vccd1 _23645_/D sky130_fd_sc_hd__a21oi_1
XFILLER_132_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21096_ _21150_/A vssd1 vssd1 vccd1 vccd1 _21096_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_320_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20047_ _23626_/Q _23625_/Q vssd1 vssd1 vccd1 vccd1 _20056_/D sky130_fd_sc_hd__and2_1
XFILLER_283_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11820_ _11863_/A _11813_/X _11817_/X _11819_/X vssd1 vssd1 vccd1 vccd1 _11826_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23806_ _23810_/CLK _23806_/D vssd1 vssd1 vccd1 vccd1 _23806_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21998_ _21999_/A _22003_/A vssd1 vssd1 vccd1 vccd1 _22000_/A sky130_fd_sc_hd__nand2_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _22368_/Q _22400_/Q _22689_/Q _23056_/Q _11745_/X _12014_/A vssd1 vssd1 vccd1
+ vccd1 _11751_/X sky130_fd_sc_hd__mux4_1
XFILLER_198_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23737_ _23874_/CLK _23737_/D vssd1 vssd1 vccd1 vccd1 _23737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20949_ _23799_/Q _20939_/X _20947_/X _20948_/X vssd1 vssd1 vccd1 vccd1 _23799_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _16171_/S vssd1 vssd1 vccd1 vccd1 _15806_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_331_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11682_ _12900_/A _11677_/X _11681_/X vssd1 vssd1 vccd1 vccd1 _11682_/X sky130_fd_sc_hd__o21a_1
X_23668_ _23704_/CLK _23668_/D vssd1 vssd1 vccd1 vccd1 _23668_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13421_ _13421_/A vssd1 vssd1 vccd1 vccd1 _15425_/A sky130_fd_sc_hd__buf_4
XFILLER_230_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22619_ _23530_/CLK _22619_/D vssd1 vssd1 vccd1 vccd1 _22619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23599_ _23599_/CLK _23599_/D vssd1 vssd1 vccd1 vccd1 _23599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16140_ _23779_/Q _14911_/A _14913_/A _16138_/X _16139_/X vssd1 vssd1 vccd1 vccd1
+ _16140_/X sky130_fd_sc_hd__a221o_1
XFILLER_344_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13352_ _13920_/A _13354_/B vssd1 vssd1 vccd1 vccd1 _13353_/C sky130_fd_sc_hd__or2b_1
XFILLER_155_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12303_ _12307_/A _12303_/B vssd1 vssd1 vccd1 vccd1 _12303_/Y sky130_fd_sc_hd__nor2_1
X_16071_ _16059_/X _14728_/B _16061_/X _16070_/Y _15558_/X vssd1 vssd1 vccd1 vccd1
+ _16071_/X sky130_fd_sc_hd__a221o_1
X_13283_ _22289_/Q _23105_/Q _23521_/Q _22450_/Q _13275_/X _13276_/X vssd1 vssd1 vccd1
+ vccd1 _13283_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15022_ _13513_/X _15996_/B _14259_/X _13514_/X _14682_/A vssd1 vssd1 vccd1 vccd1
+ _15022_/X sky130_fd_sc_hd__a221o_1
X_12234_ _12235_/A _12235_/B vssd1 vssd1 vccd1 vccd1 _12234_/X sky130_fd_sc_hd__and2_1
XFILLER_142_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_324_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19830_ _19830_/A vssd1 vssd1 vccd1 vccd1 _23550_/D sky130_fd_sc_hd__clkbuf_1
X_12165_ _21716_/A vssd1 vssd1 vccd1 vccd1 _12165_/Y sky130_fd_sc_hd__inv_2
XFILLER_296_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11116_ _11609_/A vssd1 vssd1 vccd1 vccd1 _11840_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_300_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19761_ _19252_/X _23520_/Q _19765_/S vssd1 vssd1 vccd1 vccd1 _19762_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16973_ _17028_/A vssd1 vssd1 vccd1 vccd1 _16973_/X sky130_fd_sc_hd__clkbuf_2
X_12096_ _23410_/Q _23026_/Q _23378_/Q _23346_/Q _11821_/X _11754_/A vssd1 vssd1 vccd1
+ vccd1 _12097_/B sky130_fd_sc_hd__mux4_1
XFILLER_111_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18712_ _18712_/A vssd1 vssd1 vccd1 vccd1 _23082_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15924_ _17246_/A _17229_/A _15924_/C vssd1 vssd1 vccd1 vccd1 _15940_/B sky130_fd_sc_hd__and3_1
X_19692_ _19692_/A vssd1 vssd1 vccd1 vccd1 _23489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_249_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 core_wb_ack_i vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18643_ _23052_/Q _17569_/X _18647_/S vssd1 vssd1 vccd1 vccd1 _18644_/A sky130_fd_sc_hd__mux2_1
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _16004_/A _15829_/Y _15831_/Y _15854_/X _14807_/A vssd1 vssd1 vccd1 vccd1
+ _15855_/X sky130_fd_sc_hd__o221a_1
XFILLER_264_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14806_ _15565_/A vssd1 vssd1 vccd1 vccd1 _14807_/A sky130_fd_sc_hd__clkbuf_2
X_18574_ _18574_/A vssd1 vssd1 vccd1 vccd1 _23021_/D sky130_fd_sc_hd__clkbuf_1
X_15786_ _15976_/A vssd1 vssd1 vccd1 vccd1 _15937_/S sky130_fd_sc_hd__clkbuf_4
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _12998_/A _12998_/B vssd1 vssd1 vccd1 vccd1 _12998_/X sky130_fd_sc_hd__or2_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17525_ _22669_/Q _16281_/X _17527_/S vssd1 vssd1 vccd1 vccd1 _17526_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14737_ _14745_/A _21084_/A vssd1 vssd1 vccd1 vccd1 _14737_/X sky130_fd_sc_hd__or2_1
X_11949_ _11949_/A vssd1 vssd1 vccd1 vccd1 _12746_/A sky130_fd_sc_hd__buf_4
XFILLER_220_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17456_ _17456_/A vssd1 vssd1 vccd1 vccd1 _17465_/S sky130_fd_sc_hd__buf_6
XFILLER_178_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14668_ _15130_/S vssd1 vssd1 vccd1 vccd1 _14855_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_338_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16407_ _15283_/X _22366_/Q _16407_/S vssd1 vssd1 vccd1 vccd1 _16408_/A sky130_fd_sc_hd__mux2_1
X_13619_ _13619_/A _13619_/B vssd1 vssd1 vccd1 vccd1 _15479_/B sky130_fd_sc_hd__or2_2
XFILLER_299_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17387_ _17326_/A _17326_/B _17394_/A _17325_/B vssd1 vssd1 vccd1 vccd1 _17387_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14599_ _23654_/Q _15353_/B vssd1 vssd1 vccd1 vccd1 _14599_/X sky130_fd_sc_hd__or2_1
XFILLER_257_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19126_ _19148_/A vssd1 vssd1 vccd1 vccd1 _19135_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_192_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16338_ _15372_/X _22336_/Q _16344_/S vssd1 vssd1 vccd1 vccd1 _16339_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19057_ _19057_/A vssd1 vssd1 vccd1 vccd1 _23221_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_307_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16269_ _22312_/Q _16268_/X _16269_/S vssd1 vssd1 vccd1 vccd1 _16270_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_350_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18008_ _22883_/Q vssd1 vssd1 vccd1 vccd1 _18198_/A sky130_fd_sc_hd__clkinv_2
Xoutput302 _14000_/Y vssd1 vssd1 vccd1 vccd1 addr1[8] sky130_fd_sc_hd__buf_2
XFILLER_145_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput313 _13968_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[18] sky130_fd_sc_hd__buf_2
Xoutput324 _13905_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[3] sky130_fd_sc_hd__buf_2
XFILLER_303_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput335 _13760_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[12] sky130_fd_sc_hd__buf_2
XFILLER_288_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput346 _13823_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[22] sky130_fd_sc_hd__buf_2
XFILLER_126_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput357 _13716_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[3] sky130_fd_sc_hd__buf_2
XFILLER_259_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput368 _22486_/Q vssd1 vssd1 vccd1 vccd1 core_wb_stb_o sky130_fd_sc_hd__buf_2
Xoutput379 _14037_/X vssd1 vssd1 vccd1 vccd1 din0[14] sky130_fd_sc_hd__buf_2
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_302_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_288_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19959_ _23602_/Q _19975_/B _19959_/C vssd1 vssd1 vccd1 vccd1 _19960_/B sky130_fd_sc_hd__and3_1
XFILLER_303_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22970_ _22974_/CLK _22970_/D vssd1 vssd1 vccd1 vccd1 _22970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21921_ _21829_/B _21919_/X _21920_/Y _21327_/A vssd1 vssd1 vccd1 vccd1 _21922_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_243_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21852_ _21876_/B _21877_/A vssd1 vssd1 vccd1 vccd1 _21934_/B sky130_fd_sc_hd__nor2_2
XFILLER_71_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20803_ _20806_/A _20803_/B vssd1 vssd1 vccd1 vccd1 _20804_/A sky130_fd_sc_hd__and2_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21783_ _21756_/B _21758_/B _21756_/A vssd1 vssd1 vccd1 vccd1 _21787_/A sky130_fd_sc_hd__o21ba_1
XFILLER_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23522_ _23522_/CLK _23522_/D vssd1 vssd1 vccd1 vccd1 _23522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20734_ _21078_/B _20724_/X _20733_/X vssd1 vssd1 vccd1 vccd1 _20734_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_329_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23453_ _23453_/CLK _23453_/D vssd1 vssd1 vccd1 vccd1 _23453_/Q sky130_fd_sc_hd__dfxtp_1
X_20665_ _20665_/A _20665_/B _20665_/C vssd1 vssd1 vccd1 vccd1 _20665_/X sky130_fd_sc_hd__or3_1
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22404_ _23572_/CLK _22404_/D vssd1 vssd1 vccd1 vccd1 _22404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_326_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23384_ _23575_/CLK _23384_/D vssd1 vssd1 vccd1 vccd1 _23384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_337_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20596_ _20895_/A vssd1 vssd1 vccd1 vccd1 _20631_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_136_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22335_ _23503_/CLK _22335_/D vssd1 vssd1 vccd1 vccd1 _22335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_279_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22266_ _23530_/CLK _22266_/D vssd1 vssd1 vccd1 vccd1 _22266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21217_ _21217_/A _21227_/B vssd1 vssd1 vccd1 vccd1 _21217_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22197_ _22197_/A _22197_/B vssd1 vssd1 vccd1 vccd1 _22197_/Y sky130_fd_sc_hd__nor2_1
XFILLER_183_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21148_ _21148_/A vssd1 vssd1 vccd1 vccd1 _21177_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_132_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_333_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13970_ _13970_/A _13979_/B vssd1 vssd1 vccd1 vccd1 _13971_/A sky130_fd_sc_hd__and2_1
X_21079_ _21079_/A _21079_/B _21079_/C _21079_/D vssd1 vssd1 vccd1 vccd1 _21080_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_281_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12921_ _22313_/Q _23449_/Q _12921_/S vssd1 vssd1 vccd1 vccd1 _12921_/X sky130_fd_sc_hd__mux2_1
XFILLER_246_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15640_ _15995_/A _15491_/X _15639_/X vssd1 vssd1 vccd1 vccd1 _15640_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12852_ _12852_/A _12852_/B vssd1 vssd1 vccd1 vccd1 _12852_/X sky130_fd_sc_hd__or2_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11803_ _12334_/A vssd1 vssd1 vccd1 vccd1 _12318_/A sky130_fd_sc_hd__buf_4
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _23319_/Q _23287_/Q _23255_/Q _23543_/Q _12776_/X _12777_/X vssd1 vssd1 vccd1
+ vccd1 _12784_/B sky130_fd_sc_hd__mux4_2
X_15571_ _15976_/A vssd1 vssd1 vccd1 vccd1 _15750_/S sky130_fd_sc_hd__buf_6
XFILLER_203_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17310_ _22217_/A _17309_/X _17318_/S vssd1 vssd1 vccd1 vccd1 _17310_/X sky130_fd_sc_hd__mux2_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _11742_/A vssd1 vssd1 vccd1 vccd1 _12020_/A sky130_fd_sc_hd__clkbuf_4
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ _14215_/X _21199_/A _14521_/X _14192_/B vssd1 vssd1 vccd1 vccd1 _14522_/X
+ sky130_fd_sc_hd__o211a_1
X_18290_ _18317_/A _18296_/C vssd1 vssd1 vccd1 vccd1 _18290_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _22812_/Q _17241_/B vssd1 vssd1 vccd1 vccd1 _17242_/A sky130_fd_sc_hd__nand2_2
XFILLER_203_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11665_ _23222_/Q _23190_/Q _23158_/Q _23126_/Q _11637_/X _12793_/A vssd1 vssd1 vccd1
+ vccd1 _11666_/B sky130_fd_sc_hd__mux4_2
X_14453_ _14733_/A vssd1 vssd1 vccd1 vccd1 _15590_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13404_ _13404_/A _13404_/B vssd1 vssd1 vccd1 vccd1 _13409_/B sky130_fd_sc_hd__nand2_1
XFILLER_128_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17172_ _17172_/A _17172_/B vssd1 vssd1 vccd1 vccd1 _17172_/Y sky130_fd_sc_hd__nor2_1
X_14384_ _16057_/A vssd1 vssd1 vccd1 vccd1 _14384_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_316_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11596_ _11893_/S vssd1 vssd1 vccd1 vccd1 _12755_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_183_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_317_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16123_ _18865_/A vssd1 vssd1 vccd1 vccd1 _19258_/A sky130_fd_sc_hd__buf_2
X_13335_ _13356_/A _13334_/X _12233_/X vssd1 vssd1 vccd1 vccd1 _13371_/C sky130_fd_sc_hd__o21a_1
XFILLER_182_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_343_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_289_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_331_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_316_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13266_ _13253_/A _13265_/X _11135_/A vssd1 vssd1 vccd1 vccd1 _13266_/Y sky130_fd_sc_hd__o21ai_1
X_16054_ _16054_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16054_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_331_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12217_ _23404_/Q _23020_/Q _23372_/Q _23340_/Q _12215_/X _12216_/X vssd1 vssd1 vccd1
+ vccd1 _12217_/X sky130_fd_sc_hd__mux4_1
X_15005_ _15097_/S _15005_/B vssd1 vssd1 vccd1 vccd1 _15005_/X sky130_fd_sc_hd__or2_1
XFILLER_142_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13197_ _13206_/A _13197_/B vssd1 vssd1 vccd1 vccd1 _13197_/X sky130_fd_sc_hd__or2_1
XFILLER_29_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_307_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19813_ _23543_/Q _19223_/A _19815_/S vssd1 vssd1 vccd1 vccd1 _19814_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12148_ _12780_/A _12148_/B vssd1 vssd1 vccd1 vccd1 _12148_/X sky130_fd_sc_hd__or2_1
XFILLER_97_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_340_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_300_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19744_ _19744_/A vssd1 vssd1 vccd1 vccd1 _23512_/D sky130_fd_sc_hd__clkbuf_1
X_16956_ _17268_/A vssd1 vssd1 vccd1 vccd1 _17042_/A sky130_fd_sc_hd__clkbuf_2
X_12079_ _23410_/Q _23026_/Q _23378_/Q _23346_/Q _11595_/A _11566_/A vssd1 vssd1 vccd1
+ vccd1 _12079_/X sky130_fd_sc_hd__mux4_1
XFILLER_256_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15907_ _23805_/Q _14917_/A _14919_/A vssd1 vssd1 vccd1 vccd1 _15907_/X sky130_fd_sc_hd__a21o_1
X_19675_ _19675_/A vssd1 vssd1 vccd1 vccd1 _23481_/D sky130_fd_sc_hd__clkbuf_1
X_16887_ _16886_/X _22543_/Q _16893_/S vssd1 vssd1 vccd1 vccd1 _16888_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18626_ _18682_/A vssd1 vssd1 vccd1 vccd1 _18695_/S sky130_fd_sc_hd__buf_6
XFILLER_266_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15838_ _23739_/Q _23869_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _15838_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18557_ _18557_/A vssd1 vssd1 vccd1 vccd1 _23013_/D sky130_fd_sc_hd__clkbuf_1
X_15769_ _15769_/A _15769_/B vssd1 vssd1 vccd1 vccd1 _15769_/Y sky130_fd_sc_hd__nand2_1
XFILLER_280_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17508_ _22661_/Q _16255_/X _17516_/S vssd1 vssd1 vccd1 vccd1 _17509_/A sky130_fd_sc_hd__mux2_1
X_18488_ _22991_/Q _18492_/B vssd1 vssd1 vccd1 vccd1 _18488_/Y sky130_fd_sc_hd__nand2_1
XFILLER_205_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17439_ _22631_/Q _16262_/X _17443_/S vssd1 vssd1 vccd1 vccd1 _17440_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_326_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_308_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20450_ _20470_/A vssd1 vssd1 vccd1 vccd1 _20468_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19109_ _23244_/Q _18795_/X _19113_/S vssd1 vssd1 vccd1 vccd1 _19110_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_335_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20381_ _20381_/A _20394_/B vssd1 vssd1 vccd1 vccd1 _20383_/B sky130_fd_sc_hd__nand2_1
XFILLER_284_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_323_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22120_ _21398_/X _22118_/Y _22119_/Y _21767_/X vssd1 vssd1 vccd1 vccd1 _22120_/X
+ sky130_fd_sc_hd__a211o_2
Xclkbuf_leaf_99_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23424_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_307_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_353_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_28_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23893_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22051_ _22100_/A _22051_/B vssd1 vssd1 vccd1 vccd1 _22052_/B sky130_fd_sc_hd__or2_1
XTAP_6509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21002_ _23816_/Q _21009_/B vssd1 vssd1 vccd1 vccd1 _21002_/X sky130_fd_sc_hd__or2_1
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22953_ _23602_/CLK _22953_/D vssd1 vssd1 vccd1 vccd1 _22953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21904_ _21902_/Y _21899_/Y _21898_/Y _21849_/X vssd1 vssd1 vccd1 vccd1 _21937_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_55_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22884_ _23327_/CLK _22884_/D vssd1 vssd1 vccd1 vccd1 _22884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21835_ _23830_/Q _23764_/Q vssd1 vssd1 vccd1 vccd1 _21836_/B sky130_fd_sc_hd__nor2_1
XFILLER_231_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21766_ _21766_/A _22224_/B vssd1 vssd1 vccd1 vccd1 _21766_/Y sky130_fd_sc_hd__nor2_1
XFILLER_321_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23505_ _23505_/CLK _23505_/D vssd1 vssd1 vccd1 vccd1 _23505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20717_ _23739_/Q _20697_/X _20716_/X _20706_/X vssd1 vssd1 vccd1 vccd1 _23739_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21697_ _21801_/A _21697_/B vssd1 vssd1 vccd1 vccd1 _21697_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11450_ _15864_/A _11437_/X _11444_/X _11449_/X vssd1 vssd1 vccd1 vccd1 _11451_/C
+ sky130_fd_sc_hd__a31o_1
X_23436_ _23500_/CLK _23436_/D vssd1 vssd1 vccd1 vccd1 _23436_/Q sky130_fd_sc_hd__dfxtp_1
X_20648_ _20732_/A vssd1 vssd1 vccd1 vccd1 _20648_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_137_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_354_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11381_ _21898_/A _11355_/X _20532_/B _11380_/X vssd1 vssd1 vccd1 vccd1 _20400_/A
+ sky130_fd_sc_hd__o211ai_4
X_23367_ _23367_/CLK _23367_/D vssd1 vssd1 vccd1 vccd1 _23367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_314_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20579_ _20579_/A vssd1 vssd1 vccd1 vccd1 _20580_/A sky130_fd_sc_hd__inv_2
XFILLER_165_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13120_ _23327_/Q _23295_/Q _23263_/Q _23551_/Q _11311_/A _11323_/A vssd1 vssd1 vccd1
+ vccd1 _13121_/B sky130_fd_sc_hd__mux4_1
XFILLER_178_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22318_ _23549_/CLK _22318_/D vssd1 vssd1 vccd1 vccd1 _22318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_314_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23298_ _23426_/CLK _23298_/D vssd1 vssd1 vccd1 vccd1 _23298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_313_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_341_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13051_ _13051_/A _13051_/B vssd1 vssd1 vccd1 vccd1 _13051_/Y sky130_fd_sc_hd__nor2_1
XFILLER_344_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22249_ _21294_/A _21294_/B _22249_/C _22249_/D vssd1 vssd1 vccd1 vccd1 _22249_/X
+ sky130_fd_sc_hd__and4bb_2
XFILLER_133_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12002_ _12864_/A _12002_/B _12002_/C vssd1 vssd1 vccd1 vccd1 _21773_/A sky130_fd_sc_hd__nand3_4
XFILLER_79_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_294_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16810_ input9/X _16810_/B vssd1 vssd1 vccd1 vccd1 _16810_/Y sky130_fd_sc_hd__nor2_1
X_17790_ _22770_/Q _17626_/X _17798_/S vssd1 vssd1 vccd1 vccd1 _17791_/A sky130_fd_sc_hd__mux2_1
XFILLER_289_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16741_ _16741_/A _16741_/B vssd1 vssd1 vccd1 vccd1 _16742_/A sky130_fd_sc_hd__or2_1
XFILLER_207_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13953_ _16679_/B _14099_/A vssd1 vssd1 vccd1 vccd1 _13953_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19460_ _23386_/Q _18840_/X _19466_/S vssd1 vssd1 vccd1 vccd1 _19461_/A sky130_fd_sc_hd__mux2_1
X_12904_ _12904_/A _12904_/B vssd1 vssd1 vccd1 vccd1 _12904_/X sky130_fd_sc_hd__or2_1
XFILLER_207_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16672_ _16672_/A vssd1 vssd1 vccd1 vccd1 _22482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13884_ _13884_/A _13884_/B vssd1 vssd1 vccd1 vccd1 _14071_/A sky130_fd_sc_hd__or2_4
XFILLER_74_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18411_ _19962_/A vssd1 vssd1 vccd1 vccd1 _18441_/A sky130_fd_sc_hd__clkbuf_4
X_15623_ _15615_/X _15619_/Y _15708_/S _21829_/A vssd1 vssd1 vccd1 vccd1 _18824_/A
+ sky130_fd_sc_hd__a2bb2o_4
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19391_ _19391_/A vssd1 vssd1 vccd1 vccd1 _23355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_290_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12835_ _22284_/Q _23100_/Q _23516_/Q _22445_/Q _12825_/X _12685_/X vssd1 vssd1 vccd1
+ vccd1 _12836_/B sky130_fd_sc_hd__mux4_1
XFILLER_262_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _18358_/A _18342_/B _18343_/B vssd1 vssd1 vccd1 vccd1 _22940_/D sky130_fd_sc_hd__nor3_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _23828_/Q _15211_/A _15550_/X _15553_/X _15222_/A vssd1 vssd1 vccd1 vccd1
+ _15554_/X sky130_fd_sc_hd__a221o_2
X_12766_ _23415_/Q _23031_/Q _23383_/Q _23351_/Q _12920_/A _12749_/A vssd1 vssd1 vccd1
+ vccd1 _12766_/X sky130_fd_sc_hd__mux4_2
XFILLER_199_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14505_ _22946_/Q _14499_/X _15360_/A vssd1 vssd1 vccd1 vccd1 _14505_/X sky130_fd_sc_hd__mux2_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _19932_/A vssd1 vssd1 vccd1 vccd1 _18315_/A sky130_fd_sc_hd__clkbuf_4
X_11717_ _23312_/Q _23280_/Q _23248_/Q _23536_/Q _12120_/S _11163_/A vssd1 vssd1 vccd1
+ vccd1 _11718_/B sky130_fd_sc_hd__mux4_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12697_ _12968_/A _12697_/B vssd1 vssd1 vccd1 vccd1 _12697_/Y sky130_fd_sc_hd__nor2_1
XFILLER_187_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15485_ _15485_/A _15485_/B vssd1 vssd1 vccd1 vccd1 _15830_/B sky130_fd_sc_hd__nand2_1
XFILLER_159_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_308_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17224_ _17224_/A _17224_/B vssd1 vssd1 vccd1 vccd1 _17224_/Y sky130_fd_sc_hd__nand2_1
X_11648_ _11648_/A vssd1 vssd1 vccd1 vccd1 _12029_/A sky130_fd_sc_hd__buf_2
X_14436_ _14446_/B _20989_/C vssd1 vssd1 vccd1 vccd1 _20890_/A sky130_fd_sc_hd__or2_4
XFILLER_329_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 core_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_2
XFILLER_122_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput23 core_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_2
Xinput34 core_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17155_ _22811_/Q _17241_/B vssd1 vssd1 vccd1 vccd1 _17167_/A sky130_fd_sc_hd__nand2_2
Xinput45 dout0[11] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_2
X_14367_ _14848_/A _15541_/A _14336_/X _14366_/X vssd1 vssd1 vccd1 vccd1 _14367_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_11579_ _12523_/A vssd1 vssd1 vccd1 vccd1 _12421_/A sky130_fd_sc_hd__buf_2
Xinput56 dout0[21] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__buf_2
XFILLER_183_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput67 dout0[31] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_2
Xinput78 dout0[41] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16106_ _23842_/Q _15593_/X _16102_/X _16105_/X _14738_/X vssd1 vssd1 vccd1 vccd1
+ _16106_/X sky130_fd_sc_hd__a221o_1
XFILLER_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput89 dout0[51] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13318_ _13318_/A vssd1 vssd1 vccd1 vccd1 _13548_/A sky130_fd_sc_hd__inv_2
XFILLER_116_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17086_ _14541_/X _17085_/X _17116_/S vssd1 vssd1 vccd1 vccd1 _17086_/X sky130_fd_sc_hd__mux2_1
X_14298_ _11691_/B _12168_/B _14326_/S vssd1 vssd1 vccd1 vccd1 _14298_/X sky130_fd_sc_hd__mux2_1
XFILLER_318_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_289_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16037_ _15697_/A _17279_/A _16036_/X vssd1 vssd1 vccd1 vccd1 _16037_/X sky130_fd_sc_hd__o21a_1
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13249_ _13249_/A _13249_/B vssd1 vssd1 vccd1 vccd1 _13249_/Y sky130_fd_sc_hd__nand2_1
XFILLER_131_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_297_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17988_ _22838_/Q _17972_/X _17986_/X _17987_/X _17983_/X vssd1 vssd1 vccd1 vccd1
+ _17988_/X sky130_fd_sc_hd__a221o_1
XFILLER_284_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19727_ _19727_/A vssd1 vssd1 vccd1 vccd1 _23504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16939_ _23943_/Q _17648_/B _17022_/A vssd1 vssd1 vccd1 vccd1 _16939_/X sky130_fd_sc_hd__a21o_1
XFILLER_266_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19658_ _19207_/X _23474_/Q _19660_/S vssd1 vssd1 vccd1 vccd1 _19659_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18609_ _18609_/A vssd1 vssd1 vccd1 vccd1 _23037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_252_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19589_ _19589_/A vssd1 vssd1 vccd1 vccd1 _23443_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21620_ _21618_/Y _21619_/X _14180_/B _21550_/B vssd1 vssd1 vccd1 vccd1 _21689_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_339_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21551_ _21619_/B vssd1 vssd1 vccd1 vccd1 _21867_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20502_ _20502_/A vssd1 vssd1 vccd1 vccd1 _22046_/A sky130_fd_sc_hd__buf_2
XFILLER_138_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21482_ _21482_/A vssd1 vssd1 vccd1 vccd1 _21868_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_320_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23221_ _23543_/CLK _23221_/D vssd1 vssd1 vccd1 vccd1 _23221_/Q sky130_fd_sc_hd__dfxtp_1
X_20433_ _20445_/A vssd1 vssd1 vccd1 vccd1 _20433_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_335_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23152_ _23474_/CLK _23152_/D vssd1 vssd1 vccd1 vccd1 _23152_/Q sky130_fd_sc_hd__dfxtp_1
X_20364_ _20396_/A _20364_/B vssd1 vssd1 vccd1 vccd1 _20364_/X sky130_fd_sc_hd__or2_1
XFILLER_323_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22103_ _22053_/A _22155_/A _22155_/B _22102_/Y vssd1 vssd1 vccd1 vccd1 _22104_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_106_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23083_ _23531_/CLK _23083_/D vssd1 vssd1 vccd1 vccd1 _23083_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20295_ _20295_/A vssd1 vssd1 vccd1 vccd1 _20295_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_304_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22034_ _22093_/A _22034_/B vssd1 vssd1 vccd1 vccd1 _22034_/Y sky130_fd_sc_hd__nand2_1
XTAP_6339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22936_ _22971_/CLK _22936_/D vssd1 vssd1 vccd1 vccd1 _22936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_330_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22867_ _23592_/CLK _22867_/D vssd1 vssd1 vccd1 vccd1 _22867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12620_ _23477_/Q _23573_/Q _22537_/Q _22341_/Q _12008_/X _12734_/A vssd1 vssd1 vccd1
+ vccd1 _12621_/B sky130_fd_sc_hd__mux4_2
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21818_ _23829_/Q _23763_/Q vssd1 vssd1 vccd1 vccd1 _21819_/B sky130_fd_sc_hd__or2_1
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22798_ _23448_/CLK _22798_/D vssd1 vssd1 vccd1 vccd1 _22798_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12551_ _13903_/A _13897_/A _13358_/B _12549_/X _12550_/Y vssd1 vssd1 vccd1 vccd1
+ _13356_/A sky130_fd_sc_hd__o311a_2
XFILLER_339_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21749_ _21598_/X _21748_/X _21867_/A _17133_/X vssd1 vssd1 vccd1 vccd1 _21779_/B
+ sky130_fd_sc_hd__a2bb2o_2
XPHY_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11502_ _11502_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11502_/Y sky130_fd_sc_hd__nor2_1
XFILLER_196_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15270_ _22923_/Q _14932_/X _14934_/X _22955_/Q vssd1 vssd1 vccd1 vccd1 _15270_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_196_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12482_ _12334_/A _12481_/X _11346_/A vssd1 vssd1 vccd1 vccd1 _12482_/X sky130_fd_sc_hd__o21a_1
XFILLER_346_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11433_ _13096_/A vssd1 vssd1 vccd1 vccd1 _13037_/A sky130_fd_sc_hd__clkbuf_4
X_14221_ _14234_/A vssd1 vssd1 vccd1 vccd1 _14246_/B sky130_fd_sc_hd__clkbuf_4
X_23419_ _23419_/CLK _23419_/D vssd1 vssd1 vccd1 vccd1 _23419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_327_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_295_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_327_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_314_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14152_ _22913_/Q _22912_/Q _22911_/Q vssd1 vssd1 vccd1 vccd1 _14152_/X sky130_fd_sc_hd__or3_2
XFILLER_193_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11364_ _11364_/A vssd1 vssd1 vccd1 vccd1 _11461_/A sky130_fd_sc_hd__buf_4
XFILLER_164_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13103_ _13149_/A _13102_/X _11134_/A vssd1 vssd1 vccd1 vccd1 _13103_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_217_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14083_ _14083_/A vssd1 vssd1 vccd1 vccd1 _14083_/X sky130_fd_sc_hd__buf_2
X_18960_ _16831_/X _23178_/Q _18968_/S vssd1 vssd1 vccd1 vccd1 _18961_/A sky130_fd_sc_hd__mux2_1
XFILLER_342_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11295_ _12028_/A vssd1 vssd1 vccd1 vccd1 _12784_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_313_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17911_ _22816_/Q _17908_/X _17903_/X input257/X _17899_/X vssd1 vssd1 vccd1 vccd1
+ _17911_/X sky130_fd_sc_hd__a221o_1
X_13034_ _22320_/Q _23456_/Q _13034_/S vssd1 vssd1 vccd1 vccd1 _13034_/X sky130_fd_sc_hd__mux2_1
XFILLER_313_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18891_ _18891_/A vssd1 vssd1 vccd1 vccd1 _23147_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17842_ _22793_/Q _17598_/X _17848_/S vssd1 vssd1 vccd1 vccd1 _17843_/A sky130_fd_sc_hd__mux2_1
XFILLER_294_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_294_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17773_ _17773_/A vssd1 vssd1 vccd1 vccd1 _22762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14985_ _14984_/X _22265_/Q _14985_/S vssd1 vssd1 vccd1 vccd1 _14986_/A sky130_fd_sc_hd__mux2_1
XFILLER_304_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19512_ _19204_/X _23409_/Q _19516_/S vssd1 vssd1 vccd1 vccd1 _19513_/A sky130_fd_sc_hd__mux2_1
X_16724_ _16724_/A vssd1 vssd1 vccd1 vccd1 _22495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13936_ _13942_/B _13936_/B vssd1 vssd1 vccd1 vccd1 _13936_/X sky130_fd_sc_hd__or2_2
XFILLER_240_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_502 _15052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19443_ _19443_/A vssd1 vssd1 vccd1 vccd1 _23378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_263_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_513 _17210_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16655_ _16655_/A vssd1 vssd1 vccd1 vccd1 _22474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13867_ _13892_/A _14066_/C vssd1 vssd1 vccd1 vccd1 _13867_/Y sky130_fd_sc_hd__nor2_1
XFILLER_262_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_524 _14068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_535 _23879_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15606_ _14518_/X _15587_/X _15605_/X vssd1 vssd1 vccd1 vccd1 _15606_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_546 _20234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19374_ _19396_/A vssd1 vssd1 vccd1 vccd1 _19383_/S sky130_fd_sc_hd__clkbuf_4
X_12818_ _12818_/A _12818_/B vssd1 vssd1 vccd1 vccd1 _12818_/Y sky130_fd_sc_hd__nor2_1
XINSDIODE2_557 _23469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16586_ _15861_/X _22444_/Q _16590_/S vssd1 vssd1 vccd1 vccd1 _16587_/A sky130_fd_sc_hd__mux2_1
XFILLER_188_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13798_ _13798_/A _13798_/B vssd1 vssd1 vccd1 vccd1 _13798_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18325_ _19962_/A vssd1 vssd1 vccd1 vccd1 _18360_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_203_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15537_ _13387_/B _13615_/Y _16031_/S vssd1 vssd1 vccd1 vccd1 _15537_/X sky130_fd_sc_hd__mux2_1
X_12749_ _12749_/A vssd1 vssd1 vccd1 vccd1 _12749_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18256_ _18263_/A _20134_/A vssd1 vssd1 vccd1 vccd1 _22914_/D sky130_fd_sc_hd__nor2_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15468_ _15564_/A _15468_/B vssd1 vssd1 vccd1 vccd1 _15468_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17207_ _17167_/X _17200_/X _17206_/X _17176_/X vssd1 vssd1 vccd1 vccd1 _17207_/X
+ sky130_fd_sc_hd__o211a_4
X_14419_ _23905_/Q vssd1 vssd1 vccd1 vccd1 _21526_/A sky130_fd_sc_hd__buf_6
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_329_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18187_ _18187_/A _18187_/B vssd1 vssd1 vccd1 vccd1 _18191_/B sky130_fd_sc_hd__nor2_1
XFILLER_128_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15399_ _23729_/Q _23859_/Q _15729_/S vssd1 vssd1 vccd1 vccd1 _15399_/X sky130_fd_sc_hd__mux2_1
XFILLER_351_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17138_ _17073_/A _17137_/X _17107_/X _17127_/X vssd1 vssd1 vccd1 vccd1 _17138_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_200_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_345_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_304_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_304_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_332_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17069_ _22810_/Q _17241_/B vssd1 vssd1 vccd1 vccd1 _17070_/A sky130_fd_sc_hd__nand2_2
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20080_ _20086_/A _20080_/B _20090_/D vssd1 vssd1 vccd1 vccd1 _23634_/D sky130_fd_sc_hd__nor3_1
XFILLER_298_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_350_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23770_ _23776_/CLK _23770_/D vssd1 vssd1 vccd1 vccd1 _23770_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20982_ _22217_/A _21085_/A _20762_/B _20926_/A vssd1 vssd1 vccd1 vccd1 _20982_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22721_ _23559_/CLK _22721_/D vssd1 vssd1 vccd1 vccd1 _22721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22652_ _23563_/CLK _22652_/D vssd1 vssd1 vccd1 vccd1 _22652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21603_ _16118_/A _21550_/B _21599_/Y _21601_/Y vssd1 vssd1 vccd1 vccd1 _21624_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_22_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22583_ _23649_/CLK _22583_/D vssd1 vssd1 vccd1 vccd1 _22583_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_222_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21534_ _21494_/A _21496_/B _21494_/B vssd1 vssd1 vccd1 vccd1 _21535_/B sky130_fd_sc_hd__a21bo_2
XFILLER_309_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_327_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_43_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23440_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_181_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21465_ _21465_/A vssd1 vssd1 vccd1 vccd1 _21981_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_193_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23204_ _23556_/CLK _23204_/D vssd1 vssd1 vccd1 vccd1 _23204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20416_ _20996_/A _20416_/B vssd1 vssd1 vccd1 vccd1 _20416_/Y sky130_fd_sc_hd__nand2_1
XFILLER_336_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21396_ _23784_/Q _21381_/X _21393_/X _21395_/X vssd1 vssd1 vccd1 vccd1 _21396_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_134_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23135_ _23582_/CLK _23135_/D vssd1 vssd1 vccd1 vccd1 _23135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20347_ _20347_/A _20368_/B vssd1 vssd1 vccd1 vccd1 _20347_/X sky130_fd_sc_hd__or2_1
XFILLER_351_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_296_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_350_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_350_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23066_ _23068_/CLK _23066_/D vssd1 vssd1 vccd1 vccd1 _23066_/Q sky130_fd_sc_hd__dfxtp_1
X_11080_ _11080_/A vssd1 vssd1 vccd1 vccd1 _13436_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_289_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20278_ _20272_/X _20654_/A _20277_/X _20246_/X vssd1 vssd1 vccd1 vccd1 _23666_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_6136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_289_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput202 localMemory_wb_adr_i[20] vssd1 vssd1 vccd1 vccd1 _14148_/B sky130_fd_sc_hd__buf_2
XTAP_6158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22017_ _22017_/A _22037_/B vssd1 vssd1 vccd1 vccd1 _22017_/Y sky130_fd_sc_hd__xnor2_2
XTAP_6169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput213 localMemory_wb_adr_i[9] vssd1 vssd1 vccd1 vccd1 input213/X sky130_fd_sc_hd__clkbuf_1
Xinput224 localMemory_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 input224/X sky130_fd_sc_hd__buf_6
XTAP_5435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput235 localMemory_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 input235/X sky130_fd_sc_hd__buf_8
Xinput246 localMemory_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input246/X sky130_fd_sc_hd__clkbuf_8
XTAP_5457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput257 manufacturerID[3] vssd1 vssd1 vccd1 vccd1 input257/X sky130_fd_sc_hd__buf_2
XTAP_5468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput268 partID[13] vssd1 vssd1 vccd1 vccd1 input268/X sky130_fd_sc_hd__clkbuf_1
XFILLER_276_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput279 partID[9] vssd1 vssd1 vccd1 vccd1 input279/X sky130_fd_sc_hd__clkbuf_1
XFILLER_341_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_291_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14770_ _15801_/A _16097_/B vssd1 vssd1 vccd1 vccd1 _14770_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ _23926_/Q vssd1 vssd1 vccd1 vccd1 _13616_/A sky130_fd_sc_hd__inv_2
XFILLER_327_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13721_ _13764_/A _13721_/B _14089_/A vssd1 vssd1 vccd1 vccd1 _13722_/B sky130_fd_sc_hd__nor3_4
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22919_ _22956_/CLK _22919_/D vssd1 vssd1 vccd1 vccd1 _22919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_272_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23899_ _23902_/CLK _23899_/D vssd1 vssd1 vccd1 vccd1 _23899_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16440_ _15936_/X _22381_/Q _16440_/S vssd1 vssd1 vccd1 vccd1 _16441_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13652_ _13652_/A vssd1 vssd1 vccd1 vccd1 _14224_/B sky130_fd_sc_hd__inv_12
XFILLER_140_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12603_ _13514_/A _12340_/B _13334_/C _12602_/X vssd1 vssd1 vccd1 vccd1 _12603_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _16013_/X _22351_/Q _16377_/S vssd1 vssd1 vccd1 vccd1 _16372_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13583_ _13583_/A _13983_/A _13981_/A _13979_/A vssd1 vssd1 vccd1 vccd1 _13584_/D
+ sky130_fd_sc_hd__or4_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18110_ _22875_/Q _18096_/X _18109_/X _18105_/X vssd1 vssd1 vccd1 vccd1 _22875_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_319_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_346_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15322_ _11828_/X _15048_/X _15319_/X _21641_/A _15321_/X vssd1 vssd1 vccd1 vccd1
+ _18804_/A sky130_fd_sc_hd__a32o_4
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19090_ _19090_/A _19090_/B _18770_/A vssd1 vssd1 vccd1 vccd1 _19771_/B sky130_fd_sc_hd__or3b_4
XFILLER_200_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12534_ _12534_/A _12534_/B vssd1 vssd1 vccd1 vccd1 _12534_/Y sky130_fd_sc_hd__nor2_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18041_ _22851_/Q _18036_/X _18037_/X _22984_/Q _18038_/X vssd1 vssd1 vccd1 vccd1
+ _18041_/X sky130_fd_sc_hd__a221o_1
XFILLER_185_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15253_ _15253_/A vssd1 vssd1 vccd1 vccd1 _15253_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_184_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12465_ _12465_/A _12465_/B vssd1 vssd1 vccd1 vccd1 _12465_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14204_ _14204_/A _16808_/A vssd1 vssd1 vccd1 vccd1 _19969_/B sky130_fd_sc_hd__or2b_4
XFILLER_315_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11416_ _11972_/A _20533_/B vssd1 vssd1 vccd1 vccd1 _12368_/B sky130_fd_sc_hd__or2_1
XFILLER_138_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_326_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15184_ _15119_/A _15187_/B vssd1 vssd1 vccd1 vccd1 _15485_/B sky130_fd_sc_hd__nand2b_1
X_12396_ _22263_/Q _23079_/Q _23495_/Q _22424_/Q _11647_/A _12269_/X vssd1 vssd1 vccd1
+ vccd1 _12397_/B sky130_fd_sc_hd__mux4_1
XFILLER_326_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_342_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14135_ _23011_/Q _23010_/Q vssd1 vssd1 vccd1 vccd1 _14700_/C sky130_fd_sc_hd__nor2_4
X_11347_ _11347_/A vssd1 vssd1 vccd1 vccd1 _11348_/A sky130_fd_sc_hd__buf_2
X_19992_ _20027_/A _19992_/B vssd1 vssd1 vccd1 vccd1 _19992_/Y sky130_fd_sc_hd__nor2_1
XFILLER_180_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_315_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_341_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_330_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11278_ _11278_/A vssd1 vssd1 vccd1 vccd1 _21898_/A sky130_fd_sc_hd__buf_12
X_14066_ _14074_/B _14066_/B _14066_/C vssd1 vssd1 vccd1 vccd1 _14066_/X sky130_fd_sc_hd__or3_1
X_18943_ _18943_/A vssd1 vssd1 vccd1 vccd1 _23171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_330_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13017_ _13601_/A vssd1 vssd1 vccd1 vccd1 _13018_/D sky130_fd_sc_hd__inv_2
X_18874_ _19091_/A _19018_/B vssd1 vssd1 vccd1 vccd1 _18931_/A sky130_fd_sc_hd__nor2_8
XTAP_6670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_315_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17825_ _17825_/A vssd1 vssd1 vccd1 vccd1 _22785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_295_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_227_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17756_ _17802_/S vssd1 vssd1 vccd1 vccd1 _17765_/S sky130_fd_sc_hd__clkbuf_4
X_14968_ _22499_/Q _14232_/A _14223_/X _14967_/X _15179_/A vssd1 vssd1 vccd1 vccd1
+ _14968_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_47_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16707_ _16804_/A vssd1 vssd1 vccd1 vccd1 _16723_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13919_ _13913_/A _13355_/A _13911_/X _13516_/B vssd1 vssd1 vccd1 vccd1 _13920_/B
+ sky130_fd_sc_hd__a31o_2
X_17687_ _22724_/Q _17582_/X _17693_/S vssd1 vssd1 vccd1 vccd1 _17688_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_310 _18856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14899_ _16168_/B vssd1 vssd1 vccd1 vccd1 _14988_/B sky130_fd_sc_hd__buf_2
XFILLER_262_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_321 _16107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_332 _17029_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19426_ _19426_/A vssd1 vssd1 vccd1 vccd1 _23370_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_343 _17165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16638_ _22467_/Q _16249_/X _16640_/S vssd1 vssd1 vccd1 vccd1 _16639_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_354 _22064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_365 _23472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_376 _23469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_387 input270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19357_ _23340_/Q _18795_/X _19361_/S vssd1 vssd1 vccd1 vccd1 _19358_/A sky130_fd_sc_hd__mux2_1
X_16569_ _16569_/A vssd1 vssd1 vccd1 vccd1 _22436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_398 _14090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18308_ _18316_/D vssd1 vssd1 vccd1 vccd1 _18314_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19288_ _19288_/A vssd1 vssd1 vccd1 vccd1 _23309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_337_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18239_ hold7/X _18229_/X _18238_/X _18232_/X vssd1 vssd1 vccd1 vccd1 _22907_/D sky130_fd_sc_hd__o211a_1
XFILLER_198_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_325_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21250_ _21258_/A _21250_/B vssd1 vssd1 vccd1 vccd1 _21251_/A sky130_fd_sc_hd__and2_1
XFILLER_8_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_317_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20201_ _20196_/X _20198_/X _20199_/Y _21437_/A _20200_/X vssd1 vssd1 vccd1 vccd1
+ _20585_/A sky130_fd_sc_hd__a32o_4
XFILLER_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21181_ _23875_/Q _21168_/X _21180_/X _21163_/X vssd1 vssd1 vccd1 vccd1 _23875_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_333_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20132_ _20137_/A _20132_/B _20136_/C vssd1 vssd1 vccd1 vccd1 _23650_/D sky130_fd_sc_hd__nor3_1
XFILLER_132_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_292_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20063_ _20066_/A _23627_/Q _20063_/C _20076_/D vssd1 vssd1 vccd1 vccd1 _20079_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_301_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_161_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23706_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_292_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_14 _17410_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_25 _17743_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_36 _19638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_47 _20966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_58 _21150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23822_ _23878_/CLK _23822_/D vssd1 vssd1 vccd1 vccd1 _23822_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_69 _21335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23753_ _23755_/CLK _23753_/D vssd1 vssd1 vccd1 vccd1 _23753_/Q sky130_fd_sc_hd__dfxtp_4
X_20965_ _23804_/Q _20953_/X _20962_/X _20964_/X vssd1 vssd1 vccd1 vccd1 _23804_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22704_ _23583_/CLK _22704_/D vssd1 vssd1 vccd1 vccd1 _22704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ _20970_/A vssd1 vssd1 vccd1 vccd1 _20926_/A sky130_fd_sc_hd__buf_2
X_23684_ _23684_/CLK _23684_/D vssd1 vssd1 vccd1 vccd1 _23684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22635_ _23578_/CLK _22635_/D vssd1 vssd1 vccd1 vccd1 _22635_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_241_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_356_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22566_ _22600_/CLK _22566_/D vssd1 vssd1 vccd1 vccd1 _22566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_328_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21517_ _21517_/A _21517_/B vssd1 vssd1 vccd1 vccd1 _21517_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_343_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22497_ _23704_/CLK _22497_/D vssd1 vssd1 vccd1 vccd1 _22497_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_103_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12250_ _11713_/A _12239_/Y _12241_/Y _12249_/X _11214_/A vssd1 vssd1 vccd1 vccd1
+ _12260_/B sky130_fd_sc_hd__o311a_1
X_21448_ _22012_/B _21448_/B vssd1 vssd1 vccd1 vccd1 _21485_/B sky130_fd_sc_hd__and2b_1
XFILLER_170_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11201_ _22324_/Q _23460_/Q _13254_/S vssd1 vssd1 vccd1 vccd1 _11202_/B sky130_fd_sc_hd__mux2_1
X_12181_ _12423_/A _12181_/B vssd1 vssd1 vccd1 vccd1 _12181_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_292_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21379_ _21379_/A vssd1 vssd1 vccd1 vccd1 _21379_/X sky130_fd_sc_hd__buf_2
XFILLER_312_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11132_ _11132_/A vssd1 vssd1 vccd1 vccd1 _11133_/A sky130_fd_sc_hd__buf_2
XFILLER_122_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23118_ _23502_/CLK _23118_/D vssd1 vssd1 vccd1 vccd1 _23118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_295_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_352_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15940_ _22087_/A _15940_/B vssd1 vssd1 vccd1 vccd1 _15941_/B sky130_fd_sc_hd__nor2_1
X_23049_ _23561_/CLK _23049_/D vssd1 vssd1 vccd1 vccd1 _23049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_295_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15871_ _15871_/A _15871_/B vssd1 vssd1 vccd1 vccd1 _15871_/Y sky130_fd_sc_hd__nand2_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17610_ _18836_/A vssd1 vssd1 vccd1 vccd1 _17610_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14822_ _14822_/A vssd1 vssd1 vccd1 vccd1 _14822_/X sky130_fd_sc_hd__clkbuf_2
X_18590_ _18590_/A vssd1 vssd1 vccd1 vccd1 _23028_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ _17541_/A vssd1 vssd1 vccd1 vccd1 _22676_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14753_ _14753_/A vssd1 vssd1 vccd1 vccd1 _14753_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ _11965_/A vssd1 vssd1 vccd1 vccd1 _12687_/A sky130_fd_sc_hd__buf_2
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ _13879_/B vssd1 vssd1 vccd1 vccd1 _15180_/A sky130_fd_sc_hd__buf_2
XFILLER_301_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17472_ _19091_/A _17804_/B vssd1 vssd1 vccd1 vccd1 _17529_/A sky130_fd_sc_hd__nor2_4
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14684_ _16180_/B vssd1 vssd1 vccd1 vccd1 _16131_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_233_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11896_ _12071_/A _11893_/X _11895_/X vssd1 vssd1 vccd1 vccd1 _11896_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19211_ _19210_/X _23283_/Q _19211_/S vssd1 vssd1 vccd1 vccd1 _19212_/A sky130_fd_sc_hd__mux2_1
X_16423_ _15625_/X _22373_/Q _16429_/S vssd1 vssd1 vccd1 vccd1 _16424_/A sky130_fd_sc_hd__mux2_1
XFILLER_301_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ _13967_/A _13972_/A vssd1 vssd1 vccd1 vccd1 _13636_/D sky130_fd_sc_hd__nor2_1
X_19142_ _23259_/Q _18843_/X _19146_/S vssd1 vssd1 vccd1 vccd1 _19143_/A sky130_fd_sc_hd__mux2_1
X_16354_ _16354_/A vssd1 vssd1 vccd1 vccd1 _22343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13566_ _13570_/A _13566_/B vssd1 vssd1 vccd1 vccd1 _13566_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15305_ _23759_/Q _15215_/X _15216_/X _15303_/X _15304_/X vssd1 vssd1 vccd1 vccd1
+ _15305_/X sky130_fd_sc_hd__a221o_1
X_19073_ _16892_/X _23229_/Q _19073_/S vssd1 vssd1 vccd1 vccd1 _19074_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12517_ _12506_/A _12516_/X _11678_/A vssd1 vssd1 vccd1 vccd1 _12517_/X sky130_fd_sc_hd__o21a_1
XFILLER_346_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16285_ _22317_/Q _16284_/X _16285_/S vssd1 vssd1 vccd1 vccd1 _16286_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13497_ _13497_/A vssd1 vssd1 vccd1 vccd1 _13497_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_346_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18024_ _18009_/B _18017_/X _18020_/X _22978_/Q _18023_/X vssd1 vssd1 vccd1 vccd1
+ _18024_/X sky130_fd_sc_hd__a221o_1
X_15236_ _22986_/Q _14138_/A _15164_/A input245/X vssd1 vssd1 vccd1 vccd1 _21591_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12448_ _12465_/A _12448_/B vssd1 vssd1 vccd1 vccd1 _12448_/Y sky130_fd_sc_hd__nor2_1
XFILLER_315_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_315_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_314_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15167_ _18795_/A vssd1 vssd1 vccd1 vccd1 _19188_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12379_ _23400_/Q _23016_/Q _23368_/Q _23336_/Q _11646_/A _11651_/A vssd1 vssd1 vccd1
+ vccd1 _12379_/X sky130_fd_sc_hd__mux4_1
XFILLER_315_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14118_ _14119_/B _14121_/C _14121_/D _14110_/B _17991_/A vssd1 vssd1 vccd1 vccd1
+ _17908_/A sky130_fd_sc_hd__o41a_2
XFILLER_326_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19975_ _23602_/Q _19975_/B _23598_/Q _19975_/D vssd1 vssd1 vccd1 vccd1 _19976_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_299_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15098_ _14570_/X _21217_/A _15097_/X _14521_/A vssd1 vssd1 vccd1 vccd1 _15099_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_141_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_302_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_286_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18926_ _18926_/A vssd1 vssd1 vccd1 vccd1 _23163_/D sky130_fd_sc_hd__clkbuf_1
X_14049_ _14049_/A vssd1 vssd1 vccd1 vccd1 _14049_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18857_ _23135_/Q _18856_/X _18866_/S vssd1 vssd1 vccd1 vccd1 _18858_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17808_ _17808_/A vssd1 vssd1 vccd1 vccd1 _22777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18788_ _18788_/A vssd1 vssd1 vccd1 vccd1 _18788_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_282_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17739_ _22747_/Q _17553_/X _17743_/S vssd1 vssd1 vccd1 vccd1 _17740_/A sky130_fd_sc_hd__mux2_1
XFILLER_270_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20750_ _21605_/A _20642_/A _20662_/X vssd1 vssd1 vccd1 vccd1 _20750_/X sky130_fd_sc_hd__a21o_1
XFILLER_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_140 _13022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_151 _14675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_162 _13974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19409_ _23364_/Q _18871_/X _19409_/S vssd1 vssd1 vccd1 vccd1 _19410_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_173 _17029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20681_ _17172_/A _20642_/X _20649_/X vssd1 vssd1 vccd1 vccd1 _20681_/Y sky130_fd_sc_hd__a21oi_2
XINSDIODE2_184 _14064_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_195 _13945_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22420_ _22666_/CLK _22420_/D vssd1 vssd1 vccd1 vccd1 _22420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_287_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22351_ _23551_/CLK _22351_/D vssd1 vssd1 vccd1 vccd1 _22351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_325_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21302_ _21300_/X _21301_/X _17390_/X vssd1 vssd1 vccd1 vccd1 _23911_/D sky130_fd_sc_hd__o21a_1
XFILLER_325_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22282_ _23546_/CLK _22282_/D vssd1 vssd1 vccd1 vccd1 _22282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_340_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21233_ _21233_/A _21240_/B vssd1 vssd1 vccd1 vccd1 _21233_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_305_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21164_ _23869_/Q _21139_/X _21162_/X _21163_/X vssd1 vssd1 vccd1 vccd1 _23869_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_320_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20115_ _23645_/Q _20119_/A _20101_/X vssd1 vssd1 vccd1 vccd1 _20115_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_277_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_293_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21095_ _21161_/A vssd1 vssd1 vccd1 vccd1 _21150_/A sky130_fd_sc_hd__buf_4
XFILLER_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_293_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20046_ _23625_/Q _20056_/C _23626_/Q vssd1 vssd1 vccd1 vccd1 _20049_/B sky130_fd_sc_hd__a21oi_1
XFILLER_320_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_286_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_292_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23805_ _23810_/CLK _23805_/D vssd1 vssd1 vccd1 vccd1 _23805_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ _22215_/A _21997_/B vssd1 vssd1 vccd1 vccd1 _21997_/Y sky130_fd_sc_hd__nand2_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11986_/A _11750_/B vssd1 vssd1 vccd1 vccd1 _11750_/Y sky130_fd_sc_hd__nor2_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23736_ _23866_/CLK _23736_/D vssd1 vssd1 vccd1 vccd1 _23736_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ _20948_/A vssd1 vssd1 vccd1 vccd1 _20948_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11681_/A vssd1 vssd1 vccd1 vccd1 _11681_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23667_ _23684_/CLK _23667_/D vssd1 vssd1 vccd1 vccd1 _23667_/Q sky130_fd_sc_hd__dfxtp_1
X_20879_ _20879_/A _20879_/B vssd1 vssd1 vccd1 vccd1 _20880_/A sky130_fd_sc_hd__and2_1
XFILLER_42_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13420_ _15080_/A _15081_/B vssd1 vssd1 vccd1 vccd1 _14760_/A sky130_fd_sc_hd__nor2_4
XFILLER_201_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22618_ _22618_/CLK _22618_/D vssd1 vssd1 vccd1 vccd1 _22618_/Q sky130_fd_sc_hd__dfxtp_1
X_23598_ _23600_/CLK _23598_/D vssd1 vssd1 vccd1 vccd1 _23598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_344_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13351_ _13351_/A _13351_/B vssd1 vssd1 vccd1 vccd1 _13386_/A sky130_fd_sc_hd__xnor2_2
XFILLER_328_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22549_ _23553_/CLK _22549_/D vssd1 vssd1 vccd1 vccd1 _22549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_344_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12302_ _23306_/Q _23274_/Q _23242_/Q _23530_/Q _11700_/A _11565_/A vssd1 vssd1 vccd1
+ vccd1 _12303_/B sky130_fd_sc_hd__mux4_1
X_16070_ _16070_/A _16070_/B vssd1 vssd1 vccd1 vccd1 _16070_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13282_ _13287_/A _13282_/B vssd1 vssd1 vccd1 vccd1 _13282_/Y sky130_fd_sc_hd__nor2_1
XFILLER_344_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15021_ _16054_/B vssd1 vssd1 vccd1 vccd1 _15996_/B sky130_fd_sc_hd__clkbuf_4
X_12233_ _12235_/A _12233_/B vssd1 vssd1 vccd1 vccd1 _12233_/X sky130_fd_sc_hd__or2_1
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_296_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_311_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12164_ _23924_/Q vssd1 vssd1 vccd1 vccd1 _21738_/A sky130_fd_sc_hd__buf_6
XFILLER_135_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_312_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11115_ _23900_/Q vssd1 vssd1 vccd1 vccd1 _11609_/A sky130_fd_sc_hd__buf_2
X_19760_ _19760_/A vssd1 vssd1 vccd1 vccd1 _23519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_300_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16972_ _17082_/A vssd1 vssd1 vccd1 vccd1 _17028_/A sky130_fd_sc_hd__clkbuf_4
X_12095_ _23314_/Q _23282_/Q _23250_/Q _23538_/Q _12094_/X _11755_/A vssd1 vssd1 vccd1
+ vccd1 _12095_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18711_ _16831_/X _23082_/Q _18719_/S vssd1 vssd1 vccd1 vccd1 _18712_/A sky130_fd_sc_hd__mux2_1
X_15923_ _15923_/A _15923_/B vssd1 vssd1 vccd1 vccd1 _15923_/X sky130_fd_sc_hd__or2_1
XFILLER_265_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19691_ _19255_/X _23489_/Q _19693_/S vssd1 vssd1 vccd1 vccd1 _19692_/A sky130_fd_sc_hd__mux2_1
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18642_ _18642_/A vssd1 vssd1 vccd1 vccd1 _23051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_264_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _16188_/A _15853_/Y _15673_/A vssd1 vssd1 vccd1 vccd1 _15854_/X sky130_fd_sc_hd__a21o_1
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14805_ _14804_/A _14714_/X _14804_/Y _14698_/X vssd1 vssd1 vccd1 vccd1 _14805_/X
+ sky130_fd_sc_hd__a211o_2
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _16841_/X _23021_/Q _18575_/S vssd1 vssd1 vccd1 vccd1 _18574_/A sky130_fd_sc_hd__mux2_1
X_15785_ _19229_/A vssd1 vssd1 vccd1 vccd1 _15785_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_264_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12997_ _23419_/Q _23035_/Q _23387_/Q _23355_/Q _12024_/X _12025_/X vssd1 vssd1 vccd1
+ vccd1 _12998_/B sky130_fd_sc_hd__mux4_2
XFILLER_18_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17524_ _17524_/A vssd1 vssd1 vccd1 vccd1 _22668_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14736_ _20161_/A _20989_/B vssd1 vssd1 vccd1 vccd1 _21084_/A sky130_fd_sc_hd__or2_1
XFILLER_189_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11948_ _11972_/A vssd1 vssd1 vccd1 vccd1 _12675_/A sky130_fd_sc_hd__buf_4
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17455_ _17455_/A vssd1 vssd1 vccd1 vccd1 _22638_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14667_ _14667_/A vssd1 vssd1 vccd1 vccd1 _14667_/Y sky130_fd_sc_hd__inv_2
X_11879_ _12586_/A _11879_/B vssd1 vssd1 vccd1 vccd1 _11879_/X sky130_fd_sc_hd__or2_1
XFILLER_220_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16406_ _16406_/A vssd1 vssd1 vccd1 vccd1 _22365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13618_ _13618_/A _13618_/B _13618_/C vssd1 vssd1 vccd1 vccd1 _13619_/B sky130_fd_sc_hd__and3_1
X_17386_ _17386_/A vssd1 vssd1 vccd1 vccd1 _22611_/D sky130_fd_sc_hd__clkbuf_1
X_14598_ _16102_/B vssd1 vssd1 vccd1 vccd1 _15353_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19125_ _19125_/A vssd1 vssd1 vccd1 vccd1 _23251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16337_ _16337_/A vssd1 vssd1 vccd1 vccd1 _22335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_307_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13549_ _13562_/A _13549_/B vssd1 vssd1 vccd1 vccd1 _13549_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19056_ _16867_/X _23221_/Q _19062_/S vssd1 vssd1 vccd1 vccd1 _19057_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16268_ _18833_/A vssd1 vssd1 vccd1 vccd1 _16268_/X sky130_fd_sc_hd__buf_2
XFILLER_195_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18007_ _22844_/Q _17932_/A _18006_/X _18000_/X vssd1 vssd1 vccd1 vccd1 _22844_/D
+ sky130_fd_sc_hd__o211a_1
Xoutput303 _23950_/X vssd1 vssd1 vccd1 vccd1 clk0 sky130_fd_sc_hd__clkbuf_1
X_15219_ _15219_/A vssd1 vssd1 vccd1 vccd1 _15219_/X sky130_fd_sc_hd__buf_2
Xoutput314 _13971_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[19] sky130_fd_sc_hd__buf_2
X_16199_ _16199_/A vssd1 vssd1 vccd1 vccd1 _22292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput325 _13908_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[4] sky130_fd_sc_hd__buf_2
Xoutput336 _13767_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[13] sky130_fd_sc_hd__buf_2
Xoutput347 _13828_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[23] sky130_fd_sc_hd__buf_2
Xoutput358 _13720_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[4] sky130_fd_sc_hd__buf_2
XFILLER_273_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput369 _11102_/X vssd1 vssd1 vccd1 vccd1 core_wb_we_o sky130_fd_sc_hd__buf_2
XFILLER_287_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19958_ _19975_/B _19959_/C _19957_/Y vssd1 vssd1 vccd1 vccd1 _23601_/D sky130_fd_sc_hd__o21a_1
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_330_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_287_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_353_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18909_ _18931_/A vssd1 vssd1 vccd1 vccd1 _18918_/S sky130_fd_sc_hd__buf_2
XFILLER_268_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19889_ _19900_/A vssd1 vssd1 vccd1 vccd1 _19898_/S sky130_fd_sc_hd__buf_2
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21920_ _21920_/A _22091_/B vssd1 vssd1 vccd1 vccd1 _21920_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21851_ _21849_/X _21848_/Y _21846_/Y _21844_/Y vssd1 vssd1 vccd1 vccd1 _21877_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_222_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20802_ _20613_/B _20791_/X _20792_/X _23756_/Q vssd1 vssd1 vccd1 vccd1 _20803_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21782_ _23796_/Q _21746_/X _21781_/Y _21660_/X vssd1 vssd1 vccd1 vccd1 _21782_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_230_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23521_ _23553_/CLK _23521_/D vssd1 vssd1 vccd1 vccd1 _23521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20733_ _20733_/A vssd1 vssd1 vccd1 vccd1 _20733_/X sky130_fd_sc_hd__buf_4
XFILLER_196_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23452_ _23576_/CLK _23452_/D vssd1 vssd1 vccd1 vccd1 _23452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20664_ _17133_/X _20632_/X _20663_/X vssd1 vssd1 vccd1 vccd1 _20665_/C sky130_fd_sc_hd__o21a_1
XFILLER_184_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22403_ _23441_/CLK _22403_/D vssd1 vssd1 vccd1 vccd1 _22403_/Q sky130_fd_sc_hd__dfxtp_1
X_23383_ _23446_/CLK _23383_/D vssd1 vssd1 vccd1 vccd1 _23383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20595_ _20595_/A vssd1 vssd1 vccd1 vccd1 _20597_/A sky130_fd_sc_hd__inv_2
XFILLER_13_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_353_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_326_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22334_ _23566_/CLK _22334_/D vssd1 vssd1 vccd1 vccd1 _22334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_326_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_352_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_317_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22265_ _23558_/CLK _22265_/D vssd1 vssd1 vccd1 vccd1 _22265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21216_ _21216_/A vssd1 vssd1 vccd1 vccd1 _23884_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22196_ _22195_/A _22195_/B _22195_/C vssd1 vssd1 vccd1 vccd1 _22196_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_160_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_330_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21147_ _21168_/A vssd1 vssd1 vccd1 vccd1 _21147_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_294_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21078_ _21078_/A _21078_/B _21078_/C _21078_/D vssd1 vssd1 vccd1 vccd1 _21079_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_47_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20029_ _23621_/Q _20042_/C _19962_/X vssd1 vssd1 vccd1 vccd1 _20029_/Y sky130_fd_sc_hd__a21oi_1
X_12920_ _12920_/A vssd1 vssd1 vccd1 vccd1 _12921_/S sky130_fd_sc_hd__buf_4
XFILLER_274_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _23420_/Q _23036_/Q _23388_/Q _23356_/Q _12733_/A _12710_/A vssd1 vssd1 vccd1
+ vccd1 _12852_/B sky130_fd_sc_hd__mux4_2
XFILLER_261_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11802_ _11926_/A _11802_/B vssd1 vssd1 vccd1 vccd1 _11802_/X sky130_fd_sc_hd__or2_1
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _19213_/A vssd1 vssd1 vccd1 vccd1 _15570_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12906_/A _12781_/X _11631_/X vssd1 vssd1 vccd1 vccd1 _12782_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _14521_/A _14521_/B _14521_/C vssd1 vssd1 vccd1 vccd1 _14521_/X sky130_fd_sc_hd__or3_1
XFILLER_349_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23719_ _23856_/CLK _23719_/D vssd1 vssd1 vccd1 vccd1 _23719_/Q sky130_fd_sc_hd__dfxtp_1
X_11733_ _11733_/A vssd1 vssd1 vccd1 vccd1 _11742_/A sky130_fd_sc_hd__buf_4
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _17324_/A vssd1 vssd1 vccd1 vccd1 _17240_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14500_/A _14510_/B _20770_/A vssd1 vssd1 vccd1 vccd1 _14733_/A sky130_fd_sc_hd__or3_4
XFILLER_159_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11676_/A vssd1 vssd1 vccd1 vccd1 _12793_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_175_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13403_ _13403_/A _13403_/B vssd1 vssd1 vccd1 vccd1 _13404_/B sky130_fd_sc_hd__xnor2_1
X_17171_ _14167_/X _15656_/Y _17172_/B _17170_/Y vssd1 vssd1 vccd1 vccd1 _17171_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_344_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14383_ _14762_/A vssd1 vssd1 vccd1 vccd1 _16057_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11595_ _11595_/A vssd1 vssd1 vccd1 vccd1 _11893_/S sky130_fd_sc_hd__buf_8
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16122_ _16117_/X _16119_/Y _22197_/A _15321_/X vssd1 vssd1 vccd1 vccd1 _18865_/A
+ sky130_fd_sc_hd__a2bb2o_4
X_13334_ _13510_/A _13510_/B _13334_/C _13334_/D vssd1 vssd1 vccd1 vccd1 _13334_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_328_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16053_ _13404_/B _13566_/B _16053_/S vssd1 vssd1 vccd1 vccd1 _16053_/X sky130_fd_sc_hd__mux2_1
X_13265_ _23425_/Q _23041_/Q _23393_/Q _23361_/Q _11492_/S _11200_/A vssd1 vssd1 vccd1
+ vccd1 _13265_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_331_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15004_ _14898_/X _14988_/X _14999_/X _15002_/X _15003_/X vssd1 vssd1 vccd1 vccd1
+ _15005_/B sky130_fd_sc_hd__o32a_4
X_12216_ _12216_/A vssd1 vssd1 vccd1 vccd1 _12216_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_331_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13196_ _22381_/Q _22413_/Q _22702_/Q _23069_/Q _13090_/S _13195_/X vssd1 vssd1 vccd1
+ vccd1 _13197_/B sky130_fd_sc_hd__mux4_1
XFILLER_296_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19812_ _19812_/A vssd1 vssd1 vccd1 vccd1 _23542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_285_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_307_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12147_ _23217_/Q _23185_/Q _23153_/Q _23121_/Q _11457_/C _12009_/A vssd1 vssd1 vccd1
+ vccd1 _12148_/B sky130_fd_sc_hd__mux4_1
XFILLER_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_296_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_312_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19743_ _19226_/X _23512_/Q _19743_/S vssd1 vssd1 vccd1 vccd1 _19744_/A sky130_fd_sc_hd__mux2_1
X_16955_ _16962_/A _20140_/B vssd1 vssd1 vccd1 vccd1 _17268_/A sky130_fd_sc_hd__nor2_2
X_12078_ _12082_/A _12078_/B vssd1 vssd1 vccd1 vccd1 _12078_/Y sky130_fd_sc_hd__nor2_1
XFILLER_256_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15906_ _23741_/Q _23871_/Q _16138_/S vssd1 vssd1 vccd1 vccd1 _15906_/X sky130_fd_sc_hd__mux2_1
X_16886_ _19236_/A vssd1 vssd1 vccd1 vccd1 _16886_/X sky130_fd_sc_hd__clkbuf_2
X_19674_ _19229_/X _23481_/Q _19682_/S vssd1 vssd1 vccd1 vccd1 _19675_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18625_ _19555_/B _18625_/B vssd1 vssd1 vccd1 vccd1 _18682_/A sky130_fd_sc_hd__nor2_8
X_15837_ _23675_/Q _15985_/B vssd1 vssd1 vccd1 vccd1 _15837_/X sky130_fd_sc_hd__or2_1
XFILLER_264_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15768_ _13395_/B _13633_/Y _16053_/S vssd1 vssd1 vccd1 vccd1 _15769_/B sky130_fd_sc_hd__mux2_1
X_18556_ _16813_/X _23013_/Q _18564_/S vssd1 vssd1 vccd1 vccd1 _18557_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14719_ input143/X input108/X _14719_/S vssd1 vssd1 vccd1 vccd1 _14719_/X sky130_fd_sc_hd__mux2_8
X_17507_ _17529_/A vssd1 vssd1 vccd1 vccd1 _17516_/S sky130_fd_sc_hd__buf_4
XFILLER_178_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18487_ _18480_/X _18486_/Y _18476_/X vssd1 vssd1 vccd1 vccd1 _22990_/D sky130_fd_sc_hd__a21oi_1
X_15699_ _15683_/X _15697_/Y _16188_/A vssd1 vssd1 vccd1 vccd1 _15699_/X sky130_fd_sc_hd__o21a_1
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_339_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17438_ _17438_/A vssd1 vssd1 vccd1 vccd1 _22630_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_354_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17369_ _22605_/Q input199/X _17369_/S vssd1 vssd1 vccd1 vccd1 _17370_/A sky130_fd_sc_hd__mux2_1
XFILLER_308_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_347_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19108_ _19108_/A vssd1 vssd1 vccd1 vccd1 _23243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_307_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20380_ _23680_/Q _20177_/A _20379_/Y _20360_/X vssd1 vssd1 vccd1 vccd1 _23680_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_308_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_335_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19039_ _19039_/A vssd1 vssd1 vccd1 vccd1 _23213_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_350_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_323_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_353_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22050_ _22100_/A _22051_/B vssd1 vssd1 vccd1 vccd1 _22052_/A sky130_fd_sc_hd__nand2_1
XFILLER_217_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21001_ _20570_/A _20988_/X _21000_/X _20997_/X vssd1 vssd1 vccd1 vccd1 _23815_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_287_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_68_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23575_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_269_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22952_ _23602_/CLK _22952_/D vssd1 vssd1 vccd1 vccd1 _22952_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_55_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21903_ _21849_/X _21898_/Y _21899_/Y _21902_/Y vssd1 vssd1 vccd1 vccd1 _21936_/C
+ sky130_fd_sc_hd__a211o_1
X_22883_ _23009_/CLK _22883_/D vssd1 vssd1 vccd1 vccd1 _22883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_358_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21834_ _23830_/Q _23764_/Q vssd1 vssd1 vccd1 vccd1 _21836_/A sky130_fd_sc_hd__and2_1
XFILLER_36_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21765_ _21765_/A _21765_/B vssd1 vssd1 vccd1 vccd1 _21765_/X sky130_fd_sc_hd__xor2_1
XFILLER_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23504_ _23504_/CLK _23504_/D vssd1 vssd1 vccd1 vccd1 _23504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20716_ _20727_/A _20716_/B _20716_/C vssd1 vssd1 vccd1 vccd1 _20716_/X sky130_fd_sc_hd__or3_1
XFILLER_197_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21696_ _21696_/A _21803_/A vssd1 vssd1 vccd1 vccd1 _21697_/B sky130_fd_sc_hd__or2_1
XFILLER_200_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_357_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23435_ _23467_/CLK _23435_/D vssd1 vssd1 vccd1 vccd1 _23435_/Q sky130_fd_sc_hd__dfxtp_1
X_20647_ _21025_/A _20669_/B vssd1 vssd1 vccd1 vccd1 _20652_/B sky130_fd_sc_hd__nor2_1
XFILLER_328_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11380_ _11288_/X _11367_/X _11369_/X _11373_/X _11483_/A vssd1 vssd1 vccd1 vccd1
+ _11380_/X sky130_fd_sc_hd__a311o_1
XFILLER_165_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20578_ _23719_/Q _20542_/X _20577_/X _20559_/X vssd1 vssd1 vccd1 vccd1 _23719_/D
+ sky130_fd_sc_hd__o211a_1
X_23366_ _23526_/CLK _23366_/D vssd1 vssd1 vccd1 vccd1 _23366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22317_ _23073_/CLK _22317_/D vssd1 vssd1 vccd1 vccd1 _22317_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_314_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_326_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23297_ _23453_/CLK _23297_/D vssd1 vssd1 vccd1 vccd1 _23297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_313_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13050_ _22288_/Q _23104_/Q _23520_/Q _22449_/Q _11432_/A _11435_/A vssd1 vssd1 vccd1
+ vccd1 _13051_/B sky130_fd_sc_hd__mux4_1
XFILLER_180_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22248_ _21191_/B _22247_/X _14556_/D vssd1 vssd1 vccd1 vccd1 _22257_/A sky130_fd_sc_hd__a21oi_1
XFILLER_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12001_ _11993_/X _11995_/X _11997_/X _12000_/X _11683_/X vssd1 vssd1 vccd1 vccd1
+ _12002_/C sky130_fd_sc_hd__a221o_1
XFILLER_79_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22179_ _22219_/A _22044_/X _22178_/X _22048_/X vssd1 vssd1 vccd1 vccd1 _22181_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_121_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_294_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_289_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16740_ _22500_/Q _16729_/X _16730_/X input14/X vssd1 vssd1 vccd1 vccd1 _16741_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13952_ _13918_/X _13948_/Y _13951_/Y _13924_/X vssd1 vssd1 vccd1 vccd1 _14099_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_247_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ _22282_/Q _23098_/Q _23514_/Q _22443_/Q _12776_/X _12777_/X vssd1 vssd1 vccd1
+ vccd1 _12904_/B sky130_fd_sc_hd__mux4_1
XFILLER_235_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16671_ _22482_/Q _16297_/X _16673_/S vssd1 vssd1 vccd1 vccd1 _16672_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13883_ _13892_/A _14074_/D vssd1 vssd1 vccd1 vccd1 _13883_/Y sky130_fd_sc_hd__nor2_8
XFILLER_262_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15622_ _22994_/Q _15780_/A _15781_/A input222/X vssd1 vssd1 vccd1 vccd1 _21829_/A
+ sky130_fd_sc_hd__a22o_4
X_18410_ _19923_/A _18410_/B _18412_/B vssd1 vssd1 vccd1 vccd1 _22964_/D sky130_fd_sc_hd__nor3_1
X_19390_ _23355_/Q _18843_/X _19394_/S vssd1 vssd1 vccd1 vccd1 _19391_/A sky130_fd_sc_hd__mux2_1
X_12834_ _12818_/A _12833_/X _12700_/X vssd1 vssd1 vccd1 vccd1 _12834_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _22939_/Q _22940_/Q _18341_/C vssd1 vssd1 vccd1 vccd1 _18343_/B sky130_fd_sc_hd__and3_1
XFILLER_250_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _23764_/Q _15215_/A _15216_/A _15551_/X _15552_/X vssd1 vssd1 vccd1 vccd1
+ _15553_/X sky130_fd_sc_hd__a221o_2
X_12765_ _12983_/A _12765_/B vssd1 vssd1 vccd1 vccd1 _12765_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14504_ _15835_/B vssd1 vssd1 vccd1 vccd1 _15360_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ _20067_/A vssd1 vssd1 vccd1 vccd1 _19932_/A sky130_fd_sc_hd__buf_2
XFILLER_188_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _11719_/A vssd1 vssd1 vccd1 vccd1 _12120_/S sky130_fd_sc_hd__buf_6
XFILLER_202_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15484_ _15484_/A _15484_/B vssd1 vssd1 vccd1 vccd1 _15484_/Y sky130_fd_sc_hd__nand2_2
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _22280_/Q _23096_/Q _23512_/Q _22441_/Q _12680_/X _12637_/X vssd1 vssd1 vccd1
+ vccd1 _12697_/B sky130_fd_sc_hd__mux4_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17223_ _17221_/X _17222_/Y _17318_/S vssd1 vssd1 vccd1 vccd1 _17223_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_336_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14435_ _14467_/C _14467_/B vssd1 vssd1 vccd1 vccd1 _20989_/C sky130_fd_sc_hd__or2b_2
XFILLER_187_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11647_ _11647_/A vssd1 vssd1 vccd1 vccd1 _11648_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_345_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 core_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17154_ _22568_/Q _17141_/X _17131_/X _17153_/X vssd1 vssd1 vccd1 vccd1 _22568_/D
+ sky130_fd_sc_hd__a211o_1
Xinput24 core_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_2
XFILLER_345_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput35 core_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
X_14366_ _15133_/A _14347_/X _14354_/X _14363_/Y _15249_/S vssd1 vssd1 vccd1 vccd1
+ _14366_/X sky130_fd_sc_hd__a221o_1
XFILLER_155_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11578_ _23901_/Q vssd1 vssd1 vccd1 vccd1 _12523_/A sky130_fd_sc_hd__clkbuf_4
Xinput46 dout0[12] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_2
Xinput57 dout0[22] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_2
Xinput68 dout0[32] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16105_ _23778_/Q _15595_/X _15596_/X _16103_/X _16104_/X vssd1 vssd1 vccd1 vccd1
+ _16105_/X sky130_fd_sc_hd__a221o_1
X_13317_ _13555_/A _13317_/B vssd1 vssd1 vccd1 vccd1 _13410_/B sky130_fd_sc_hd__xnor2_2
XFILLER_344_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17085_ _23470_/Q _17061_/X _17062_/X _17042_/X _15271_/X vssd1 vssd1 vccd1 vccd1
+ _17085_/X sky130_fd_sc_hd__a32o_1
Xinput79 dout0[42] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__clkbuf_1
X_14297_ _12171_/B _12636_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _14297_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_331_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16036_ _14682_/X _16031_/X _16035_/X _14801_/A vssd1 vssd1 vccd1 vccd1 _16036_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_304_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13248_ _14276_/B vssd1 vssd1 vccd1 vccd1 _13249_/B sky130_fd_sc_hd__inv_2
XFILLER_272_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13179_ _22802_/Q _22770_/Q _22671_/Q _22738_/Q _11543_/A _13127_/X vssd1 vssd1 vccd1
+ vccd1 _13180_/B sky130_fd_sc_hd__mux4_2
XFILLER_312_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_300_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_313_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17987_ input3/X input269/X _17987_/S vssd1 vssd1 vccd1 vccd1 _17987_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19726_ _19201_/X _23504_/Q _19732_/S vssd1 vssd1 vccd1 vccd1 _19727_/A sky130_fd_sc_hd__mux2_1
X_16938_ _16941_/A _16941_/B _16958_/B _16938_/D vssd1 vssd1 vccd1 vccd1 _17022_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_244_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19657_ _19657_/A vssd1 vssd1 vccd1 vccd1 _23473_/D sky130_fd_sc_hd__clkbuf_1
X_16869_ _16869_/A vssd1 vssd1 vccd1 vccd1 _22537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18608_ _16892_/X _23037_/Q _18608_/S vssd1 vssd1 vccd1 vccd1 _18609_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19588_ _23443_/Q _19210_/A _19588_/S vssd1 vssd1 vccd1 vccd1 _19589_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18539_ _22877_/Q _22876_/Q _22872_/Q vssd1 vssd1 vccd1 vccd1 _18539_/X sky130_fd_sc_hd__o21ba_1
XFILLER_252_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_186_wb_clk_i clkbuf_opt_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23907_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_339_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21550_ _21550_/A _21550_/B vssd1 vssd1 vccd1 vccd1 _21558_/A sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_115_wb_clk_i _22899_/CLK vssd1 vssd1 vccd1 vccd1 _23008_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_179_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20501_ _14195_/A _21336_/A _21482_/A vssd1 vssd1 vccd1 vccd1 _20502_/A sky130_fd_sc_hd__a21oi_2
XFILLER_339_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21481_ _22012_/B _21526_/A vssd1 vssd1 vccd1 vccd1 _21481_/X sky130_fd_sc_hd__or2b_1
XFILLER_355_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_336_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23220_ _23543_/CLK _23220_/D vssd1 vssd1 vccd1 vccd1 _23220_/Q sky130_fd_sc_hd__dfxtp_1
X_20432_ _21013_/A _20463_/B vssd1 vssd1 vccd1 vccd1 _20432_/Y sky130_fd_sc_hd__nand2_1
XFILLER_295_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23151_ _23535_/CLK _23151_/D vssd1 vssd1 vccd1 vccd1 _23151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20363_ _17258_/A _20261_/X _20364_/B vssd1 vssd1 vccd1 vccd1 _20363_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_335_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22102_ _22231_/A _22075_/B _22052_/A vssd1 vssd1 vccd1 vccd1 _22102_/Y sky130_fd_sc_hd__o21ai_1
XTAP_7019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23082_ _23530_/CLK _23082_/D vssd1 vssd1 vccd1 vccd1 _23082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_311_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20294_ _20307_/A vssd1 vssd1 vccd1 vccd1 _20294_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_304_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_350_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22033_ _21569_/X _22031_/Y _22032_/Y _21577_/X vssd1 vssd1 vccd1 vccd1 _22034_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_322_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22935_ _22947_/CLK _22935_/D vssd1 vssd1 vccd1 vccd1 _22935_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_113_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22866_ _23592_/CLK _22866_/D vssd1 vssd1 vccd1 vccd1 _22866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21817_ _23829_/Q _23763_/Q vssd1 vssd1 vccd1 vccd1 _21819_/A sky130_fd_sc_hd__nand2_1
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22797_ _23449_/CLK _22797_/D vssd1 vssd1 vccd1 vccd1 _22797_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12550_ _14313_/A _13502_/A vssd1 vssd1 vccd1 vccd1 _12550_/Y sky130_fd_sc_hd__nand2_1
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21748_ _20279_/A _21870_/A _15482_/Y _21842_/A vssd1 vssd1 vccd1 vccd1 _21748_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_358_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_339_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11501_ _23330_/Q _23298_/Q _23266_/Q _23554_/Q _11432_/X _11435_/X vssd1 vssd1 vccd1
+ vccd1 _11502_/B sky130_fd_sc_hd__mux4_2
XPHY_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12481_ _23398_/Q _23014_/Q _23366_/Q _23334_/Q _12475_/X _12329_/A vssd1 vssd1 vccd1
+ vccd1 _12481_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21679_ _21981_/A _21679_/B vssd1 vssd1 vccd1 vccd1 _21679_/Y sky130_fd_sc_hd__nand2_1
XFILLER_200_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14220_ _14220_/A _14224_/A _22611_/Q vssd1 vssd1 vccd1 vccd1 _14234_/A sky130_fd_sc_hd__or3b_1
XFILLER_138_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_327_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23418_ _23548_/CLK _23418_/D vssd1 vssd1 vccd1 vccd1 _23418_/Q sky130_fd_sc_hd__dfxtp_1
X_11432_ _11432_/A vssd1 vssd1 vccd1 vccd1 _11432_/X sky130_fd_sc_hd__buf_6
XFILLER_138_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_326_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_327_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14151_ _14161_/A vssd1 vssd1 vccd1 vccd1 _14151_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_342_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23349_ _23349_/CLK _23349_/D vssd1 vssd1 vccd1 vccd1 _23349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_299_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11363_ _13184_/A vssd1 vssd1 vccd1 vccd1 _20532_/B sky130_fd_sc_hd__buf_8
XFILLER_137_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13102_ _23423_/Q _23039_/Q _23391_/Q _23359_/Q _11205_/A _13085_/X vssd1 vssd1 vccd1
+ vccd1 _13102_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_341_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14082_ _14082_/A vssd1 vssd1 vccd1 vccd1 _14082_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_314_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11294_ _11914_/A vssd1 vssd1 vccd1 vccd1 _12028_/A sky130_fd_sc_hd__buf_4
XFILLER_301_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17910_ _22816_/Q _17891_/X _17909_/X _17657_/X vssd1 vssd1 vccd1 vccd1 _22816_/D
+ sky130_fd_sc_hd__o211a_1
X_13033_ _13089_/A vssd1 vssd1 vccd1 vccd1 _13034_/S sky130_fd_sc_hd__buf_6
X_18890_ _23147_/Q _18792_/X _18896_/S vssd1 vssd1 vccd1 vccd1 _18891_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17841_ _17841_/A vssd1 vssd1 vccd1 vccd1 _22792_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_294_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_294_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17772_ _22762_/Q _17601_/X _17776_/S vssd1 vssd1 vccd1 vccd1 _17773_/A sky130_fd_sc_hd__mux2_1
XFILLER_254_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14984_ _19178_/A vssd1 vssd1 vccd1 vccd1 _14984_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_266_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19511_ _19511_/A vssd1 vssd1 vccd1 vccd1 _23408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16723_ _16723_/A _16723_/B vssd1 vssd1 vccd1 vccd1 _16724_/A sky130_fd_sc_hd__or2_1
X_13935_ _13935_/A _13935_/B _13935_/C vssd1 vssd1 vccd1 vccd1 _13936_/B sky130_fd_sc_hd__and3_1
XFILLER_263_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16654_ _22474_/Q _16271_/X _16662_/S vssd1 vssd1 vccd1 vccd1 _16655_/A sky130_fd_sc_hd__mux2_1
X_19442_ _23378_/Q _18814_/X _19444_/S vssd1 vssd1 vccd1 vccd1 _19443_/A sky130_fd_sc_hd__mux2_1
XFILLER_262_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_503 _15054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13866_ _13863_/Y _13864_/Y _13865_/X vssd1 vssd1 vccd1 vccd1 _14066_/C sky130_fd_sc_hd__o21ai_4
XFILLER_90_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_514 _23471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_525 _14070_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_320_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15605_ _18314_/A _14868_/B _15604_/X _14898_/X vssd1 vssd1 vccd1 vccd1 _15605_/X
+ sky130_fd_sc_hd__a211o_1
XINSDIODE2_536 _23883_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_343_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12817_ _22800_/Q _22768_/Q _22669_/Q _22736_/Q _12692_/X _11594_/A vssd1 vssd1 vccd1
+ vccd1 _12818_/B sky130_fd_sc_hd__mux4_2
X_16585_ _16585_/A vssd1 vssd1 vccd1 vccd1 _22443_/D sky130_fd_sc_hd__clkbuf_1
X_19373_ _19373_/A vssd1 vssd1 vccd1 vccd1 _23347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_547 _21900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13797_ _13890_/B vssd1 vssd1 vccd1 vccd1 _14241_/A sky130_fd_sc_hd__buf_2
XINSDIODE2_558 _23943_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_304_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18324_ _18358_/A _18324_/B _18326_/B vssd1 vssd1 vccd1 vccd1 _22934_/D sky130_fd_sc_hd__nor3_1
XFILLER_31_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15536_ _15918_/S vssd1 vssd1 vccd1 vccd1 _16031_/S sky130_fd_sc_hd__clkbuf_2
X_12748_ _12985_/A _12748_/B vssd1 vssd1 vccd1 vccd1 _12748_/Y sky130_fd_sc_hd__nor2_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_337_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_309_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18255_ _22914_/Q vssd1 vssd1 vccd1 vccd1 _18263_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_188_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15467_ _15431_/X _15465_/X _16154_/A vssd1 vssd1 vccd1 vccd1 _15468_/B sky130_fd_sc_hd__mux2_1
XFILLER_337_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12679_ _12698_/A vssd1 vssd1 vccd1 vccd1 _12926_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_176_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17206_ _17169_/X _17205_/X _17195_/X _17127_/X vssd1 vssd1 vccd1 vccd1 _17206_/X
+ sky130_fd_sc_hd__a211o_1
X_14418_ _20161_/A _14500_/A vssd1 vssd1 vccd1 vccd1 _14510_/A sky130_fd_sc_hd__or2_1
X_18186_ _18195_/A _18186_/B vssd1 vssd1 vccd1 vccd1 _18186_/X sky130_fd_sc_hd__and2_1
XFILLER_129_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_345_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15398_ _23665_/Q _16170_/B vssd1 vssd1 vccd1 vccd1 _15398_/X sky130_fd_sc_hd__or2_1
XFILLER_200_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_329_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17137_ _17133_/X _17136_/X _17137_/S vssd1 vssd1 vccd1 vccd1 _17137_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_317_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14349_ _11555_/A _13364_/A _14358_/A vssd1 vssd1 vccd1 vccd1 _14349_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_289_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17068_ _22560_/Q _17038_/X _17028_/X _17067_/X vssd1 vssd1 vccd1 vccd1 _22560_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_116_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_332_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16019_ _22973_/Q _16070_/A vssd1 vssd1 vccd1 vccd1 _16019_/X sky130_fd_sc_hd__or2_1
XFILLER_170_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_298_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_297_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19709_ _19709_/A vssd1 vssd1 vccd1 vccd1 _23496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20981_ _23810_/Q _20969_/X _20980_/X _20978_/X vssd1 vssd1 vccd1 vccd1 _23810_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22720_ _23048_/CLK _22720_/D vssd1 vssd1 vccd1 vccd1 _22720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_281_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22651_ _23144_/CLK _22651_/D vssd1 vssd1 vccd1 vccd1 _22651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21602_ _21599_/Y _21601_/Y _16118_/A _21550_/B vssd1 vssd1 vccd1 vccd1 _21604_/A
+ sky130_fd_sc_hd__o211a_1
X_22582_ _23646_/CLK _22582_/D vssd1 vssd1 vccd1 vccd1 _22582_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_159_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21533_ _21533_/A _21533_/B vssd1 vssd1 vccd1 vccd1 _21535_/A sky130_fd_sc_hd__nand2_1
XFILLER_138_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_327_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21464_ _23818_/Q _21838_/A _21463_/Y _21377_/A vssd1 vssd1 vccd1 vccd1 _21464_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_308_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23203_ _23459_/CLK _23203_/D vssd1 vssd1 vccd1 vccd1 _23203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_308_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20415_ _20491_/B vssd1 vssd1 vccd1 vccd1 _20416_/B sky130_fd_sc_hd__buf_4
XFILLER_162_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21395_ _22129_/A vssd1 vssd1 vccd1 vccd1 _21395_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_335_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_324_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_323_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23134_ _23550_/CLK _23134_/D vssd1 vssd1 vccd1 vccd1 _23134_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_83_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23100_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_190_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20346_ _20333_/X _20713_/A _20345_/X _20324_/X vssd1 vssd1 vccd1 vccd1 _23675_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_12_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23565_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23065_ _23449_/CLK _23065_/D vssd1 vssd1 vccd1 vccd1 _23065_/Q sky130_fd_sc_hd__dfxtp_1
X_20277_ _23666_/Q _20277_/B vssd1 vssd1 vccd1 vccd1 _20277_/X sky130_fd_sc_hd__or2_1
XTAP_6126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22016_ _22231_/A _22041_/D vssd1 vssd1 vccd1 vccd1 _22037_/B sky130_fd_sc_hd__xnor2_1
Xinput203 localMemory_wb_adr_i[21] vssd1 vssd1 vccd1 vccd1 _14148_/A sky130_fd_sc_hd__buf_2
XTAP_6159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput214 localMemory_wb_cyc_i vssd1 vssd1 vccd1 vccd1 _17326_/A sky130_fd_sc_hd__clkbuf_2
Xinput225 localMemory_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 input225/X sky130_fd_sc_hd__buf_6
XTAP_5436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput236 localMemory_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 input236/X sky130_fd_sc_hd__buf_8
XTAP_5447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput247 localMemory_wb_sel_i[0] vssd1 vssd1 vccd1 vccd1 input247/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput258 manufacturerID[4] vssd1 vssd1 vccd1 vccd1 input258/X sky130_fd_sc_hd__buf_2
XTAP_5469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput269 partID[14] vssd1 vssd1 vccd1 vccd1 input269/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ _11543_/X _12913_/S _11401_/A _11980_/Y vssd1 vssd1 vccd1 vccd1 _12171_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13720_ _13720_/A vssd1 vssd1 vccd1 vccd1 _13720_/X sky130_fd_sc_hd__clkbuf_1
X_22918_ _22956_/CLK _22918_/D vssd1 vssd1 vccd1 vccd1 _22918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_354_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23898_ _23903_/CLK _23898_/D vssd1 vssd1 vccd1 vccd1 _23898_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_272_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13651_ _17385_/B _13651_/B vssd1 vssd1 vccd1 vccd1 _13651_/Y sky130_fd_sc_hd__nand2_1
XFILLER_216_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22849_ _23426_/CLK _22849_/D vssd1 vssd1 vccd1 vccd1 _22849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12602_ _12602_/A _14368_/A vssd1 vssd1 vccd1 vccd1 _12602_/X sky130_fd_sc_hd__or2b_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _16370_/A vssd1 vssd1 vccd1 vccd1 _22350_/D sky130_fd_sc_hd__clkbuf_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13582_ _13562_/A _17246_/A _13490_/X _13581_/Y vssd1 vssd1 vccd1 vccd1 _13979_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_358_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15321_ _15746_/A vssd1 vssd1 vccd1 vccd1 _15321_/X sky130_fd_sc_hd__buf_2
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12533_ _23205_/Q _23173_/Q _23141_/Q _23109_/Q _11146_/A _11701_/A vssd1 vssd1 vccd1
+ vccd1 _12534_/B sky130_fd_sc_hd__mux4_1
XFILLER_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_346_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18040_ _22851_/Q _18035_/X _18039_/X _18029_/X vssd1 vssd1 vccd1 vccd1 _22851_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15252_ _15252_/A vssd1 vssd1 vccd1 vccd1 _15252_/Y sky130_fd_sc_hd__inv_2
X_12464_ _23206_/Q _23174_/Q _23142_/Q _23110_/Q _12537_/S _12449_/X vssd1 vssd1 vccd1
+ vccd1 _12465_/B sky130_fd_sc_hd__mux4_2
XFILLER_8_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14203_ _22520_/Q _22519_/Q vssd1 vssd1 vccd1 vccd1 _16808_/A sky130_fd_sc_hd__nand2_8
X_11415_ _11894_/S vssd1 vssd1 vccd1 vccd1 _11972_/A sky130_fd_sc_hd__buf_6
XFILLER_327_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15183_ _15183_/A vssd1 vssd1 vccd1 vccd1 _15183_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12395_ _14313_/A _13502_/A vssd1 vssd1 vccd1 vccd1 _13903_/A sky130_fd_sc_hd__xnor2_4
XFILLER_4_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14134_ _14433_/S vssd1 vssd1 vccd1 vccd1 _14421_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11346_ _11346_/A vssd1 vssd1 vccd1 vccd1 _11347_/A sky130_fd_sc_hd__clkbuf_4
X_19991_ _23610_/Q _19994_/C vssd1 vssd1 vccd1 vccd1 _19992_/B sky130_fd_sc_hd__and2_1
XFILLER_299_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_298_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_314_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_286_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14065_ input235/X _14058_/X _14064_/X vssd1 vssd1 vccd1 vccd1 _14065_/X sky130_fd_sc_hd__a21bo_4
X_18942_ _23171_/Q _18868_/X _18944_/S vssd1 vssd1 vccd1 vccd1 _18943_/A sky130_fd_sc_hd__mux2_1
XTAP_7350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11277_ _11277_/A vssd1 vssd1 vccd1 vccd1 _11278_/A sky130_fd_sc_hd__clkbuf_8
XTAP_7361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13016_ _13492_/D vssd1 vssd1 vccd1 vccd1 _13601_/A sky130_fd_sc_hd__buf_4
XTAP_7383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18873_ _18873_/A vssd1 vssd1 vccd1 vccd1 _23140_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_315_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17824_ _22785_/Q _17572_/X _17826_/S vssd1 vssd1 vccd1 vccd1 _17825_/A sky130_fd_sc_hd__mux2_1
XFILLER_294_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_67_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14967_ input145/X input110/X _14967_/S vssd1 vssd1 vccd1 vccd1 _14967_/X sky130_fd_sc_hd__mux2_8
XFILLER_208_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17755_ _17755_/A vssd1 vssd1 vccd1 vccd1 _22754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_254_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_331_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16706_ _16779_/A vssd1 vssd1 vccd1 vccd1 _16804_/A sky130_fd_sc_hd__buf_4
XFILLER_331_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13918_ _13951_/A vssd1 vssd1 vccd1 vccd1 _13918_/X sky130_fd_sc_hd__clkbuf_2
X_14898_ _14898_/A vssd1 vssd1 vccd1 vccd1 _14898_/X sky130_fd_sc_hd__buf_2
XFILLER_208_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17686_ _17686_/A vssd1 vssd1 vccd1 vccd1 _22723_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_300 _15990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_311 _18856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19425_ _23370_/Q _18788_/X _19433_/S vssd1 vssd1 vccd1 vccd1 _19426_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_322 _16107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16637_ _16637_/A vssd1 vssd1 vccd1 vccd1 _22466_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_333 _17041_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13849_ _13846_/Y _13847_/Y _13848_/X vssd1 vssd1 vccd1 vccd1 _14061_/C sky130_fd_sc_hd__o21ai_4
XINSDIODE2_344 _17179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_355 _22116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_366 _23472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_377 _23470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19356_ _19356_/A vssd1 vssd1 vccd1 vccd1 _23339_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_388 input280/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16568_ _15523_/X _22436_/Q _16568_/S vssd1 vssd1 vccd1 vccd1 _16569_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_399 _14094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_337_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18307_ _22927_/Q _22928_/Q _22929_/Q _18307_/D vssd1 vssd1 vccd1 vccd1 _18316_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_176_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15519_ _15519_/A vssd1 vssd1 vccd1 vccd1 _16195_/S sky130_fd_sc_hd__buf_2
XFILLER_349_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16499_ _16499_/A vssd1 vssd1 vccd1 vccd1 _22406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19287_ _19191_/X _23309_/Q _19289_/S vssd1 vssd1 vccd1 vccd1 _19288_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18238_ _22907_/Q _18240_/B vssd1 vssd1 vccd1 vccd1 _18238_/X sky130_fd_sc_hd__or2_1
XFILLER_136_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18169_ _18178_/B _18187_/B _18144_/B _18142_/A _18181_/A vssd1 vssd1 vccd1 vccd1
+ _18169_/X sky130_fd_sc_hd__o221a_1
XFILLER_191_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_317_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20200_ _20307_/A vssd1 vssd1 vccd1 vccd1 _20200_/X sky130_fd_sc_hd__clkbuf_2
X_21180_ _21083_/A _20509_/A _21140_/X _20749_/A _21161_/X vssd1 vssd1 vccd1 vccd1
+ _21180_/X sky130_fd_sc_hd__a221o_1
XFILLER_172_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_289_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_320_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20131_ _23650_/Q _23649_/Q _23648_/Q _20131_/D vssd1 vssd1 vccd1 vccd1 _20136_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_144_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_321_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20062_ _23630_/Q _23629_/Q vssd1 vssd1 vccd1 vccd1 _20076_/D sky130_fd_sc_hd__and2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_15 _17483_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_300_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_26 _17743_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_37 _19638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_48 _20966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23821_ _23832_/CLK _23821_/D vssd1 vssd1 vccd1 vccd1 _23821_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_245_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_59 _21150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23752_ _23911_/CLK _23752_/D vssd1 vssd1 vccd1 vccd1 _23752_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_130_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _22956_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_214_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20964_ _21023_/A vssd1 vssd1 vccd1 vccd1 _20964_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22703_ _23070_/CLK _22703_/D vssd1 vssd1 vccd1 vccd1 _22703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23683_ _23706_/CLK _23683_/D vssd1 vssd1 vccd1 vccd1 _23683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20895_ _20895_/A _20895_/B vssd1 vssd1 vccd1 vccd1 _20970_/A sky130_fd_sc_hd__nor2_4
XFILLER_198_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22634_ _23577_/CLK _22634_/D vssd1 vssd1 vccd1 vccd1 _22634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22565_ _22600_/CLK _22565_/D vssd1 vssd1 vccd1 vccd1 _22565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_326_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_356_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21516_ _21515_/B _21514_/Y _21515_/Y _21327_/X vssd1 vssd1 vccd1 vccd1 _21516_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_357_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22496_ _23714_/CLK _22496_/D vssd1 vssd1 vccd1 vccd1 _22496_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_194_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_343_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21447_ _21480_/S vssd1 vssd1 vccd1 vccd1 _22012_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_336_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11200_ _11200_/A vssd1 vssd1 vccd1 vccd1 _14393_/A sky130_fd_sc_hd__buf_4
XFILLER_107_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12180_ _22461_/Q _22621_/Q _12349_/S vssd1 vssd1 vccd1 vccd1 _12181_/B sky130_fd_sc_hd__mux2_1
X_21378_ _23816_/Q _21418_/A _21374_/Y _21377_/X vssd1 vssd1 vccd1 vccd1 _21378_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_253_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11131_ _11131_/A vssd1 vssd1 vccd1 vccd1 _11132_/A sky130_fd_sc_hd__buf_2
XFILLER_253_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23117_ _23407_/CLK _23117_/D vssd1 vssd1 vccd1 vccd1 _23117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20329_ _20355_/A _20329_/B vssd1 vssd1 vccd1 vccd1 _20329_/Y sky130_fd_sc_hd__nand2_1
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_295_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23048_ _23048_/CLK _23048_/D vssd1 vssd1 vccd1 vccd1 _23048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_292_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15870_ _14839_/A _15195_/X _15194_/X _15338_/A vssd1 vssd1 vccd1 vccd1 _15871_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_103_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14821_ _15698_/A _14821_/B vssd1 vssd1 vccd1 vccd1 _14822_/A sky130_fd_sc_hd__nor2_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _14752_/A vssd1 vssd1 vccd1 vccd1 _14752_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_233_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17540_ _22676_/Q _16303_/X _17542_/S vssd1 vssd1 vccd1 vccd1 _17541_/A sky130_fd_sc_hd__mux2_1
X_11964_ _22372_/Q _22404_/Q _22693_/Q _23060_/Q _12825_/A _12756_/A vssd1 vssd1 vccd1
+ vccd1 _11964_/X sky130_fd_sc_hd__mux4_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _13728_/B vssd1 vssd1 vccd1 vccd1 _13786_/A sky130_fd_sc_hd__clkbuf_1
X_17471_ _17471_/A _17471_/B _19090_/A vssd1 vssd1 vccd1 vccd1 _17804_/B sky130_fd_sc_hd__nand3_4
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14683_ _14385_/B _14371_/Y _14175_/Y vssd1 vssd1 vccd1 vccd1 _16180_/B sky130_fd_sc_hd__o21a_2
XFILLER_232_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11895_ _11621_/X _11894_/X _11853_/A vssd1 vssd1 vccd1 vccd1 _11895_/X sky130_fd_sc_hd__a21o_1
XFILLER_17_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19210_ _19210_/A vssd1 vssd1 vccd1 vccd1 _19210_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16422_ _16422_/A vssd1 vssd1 vccd1 vccd1 _22372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13634_ _21950_/A _13588_/A _13633_/Y _13594_/A vssd1 vssd1 vccd1 vccd1 _13972_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_232_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19141_ _19141_/A vssd1 vssd1 vccd1 vccd1 _23258_/D sky130_fd_sc_hd__clkbuf_1
X_16353_ _15710_/X _22343_/Q _16355_/S vssd1 vssd1 vccd1 vccd1 _16354_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13565_ _13565_/A _13565_/B vssd1 vssd1 vccd1 vccd1 _13566_/B sky130_fd_sc_hd__xnor2_4
XFILLER_301_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15304_ _23791_/Q _15219_/X _14606_/X vssd1 vssd1 vccd1 vccd1 _15304_/X sky130_fd_sc_hd__a21o_1
X_19072_ _19072_/A vssd1 vssd1 vccd1 vccd1 _23228_/D sky130_fd_sc_hd__clkbuf_1
X_12516_ _22454_/Q _22614_/Q _22293_/Q _23429_/Q _12501_/X _12502_/X vssd1 vssd1 vccd1
+ vccd1 _12516_/X sky130_fd_sc_hd__mux4_2
X_16284_ _18849_/A vssd1 vssd1 vccd1 vccd1 _16284_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13496_ _12868_/A _13015_/B _13494_/X _13495_/Y vssd1 vssd1 vccd1 vccd1 _13540_/A
+ sky130_fd_sc_hd__o31a_2
X_18023_ _18054_/A vssd1 vssd1 vccd1 vccd1 _18023_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15235_ _14819_/X _15232_/X _15234_/Y _15162_/X vssd1 vssd1 vccd1 vccd1 _15235_/X
+ sky130_fd_sc_hd__a211o_1
X_12447_ _23462_/Q _23558_/Q _22522_/Q _22326_/Q _11411_/A _11189_/A vssd1 vssd1 vccd1
+ vccd1 _12448_/B sky130_fd_sc_hd__mux4_1
XFILLER_346_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15166_ _12230_/X _15048_/X _15163_/X _21515_/A _15041_/X vssd1 vssd1 vccd1 vccd1
+ _18795_/A sky130_fd_sc_hd__a32o_4
X_12378_ _12378_/A _12378_/B vssd1 vssd1 vccd1 vccd1 _12378_/X sky130_fd_sc_hd__or2_1
XFILLER_330_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_342_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14117_ _14119_/A _22888_/Q _22887_/Q _14119_/D vssd1 vssd1 vccd1 vccd1 _17991_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_315_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11329_ _12489_/A vssd1 vssd1 vccd1 vccd1 _11330_/A sky130_fd_sc_hd__buf_2
X_19974_ _23606_/Q _19980_/C vssd1 vssd1 vccd1 vccd1 _19979_/B sky130_fd_sc_hd__nor2_1
XFILLER_125_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15097_ _17052_/A _15096_/X _15097_/S vssd1 vssd1 vccd1 vccd1 _15097_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18925_ _23163_/Q _18843_/X _18929_/S vssd1 vssd1 vccd1 vccd1 _18926_/A sky130_fd_sc_hd__mux2_1
X_14048_ _14023_/X _13812_/B _14041_/X input227/X vssd1 vssd1 vccd1 vccd1 _14048_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_7180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18856_ _18856_/A vssd1 vssd1 vccd1 vccd1 _18856_/X sky130_fd_sc_hd__clkbuf_2
XTAP_6490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17807_ _22777_/Q _17544_/X _17815_/S vssd1 vssd1 vccd1 vccd1 _17808_/A sky130_fd_sc_hd__mux2_1
XFILLER_342_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18787_ _18787_/A vssd1 vssd1 vccd1 vccd1 _23113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15999_ _16097_/A _15013_/X _15998_/X _15636_/X vssd1 vssd1 vccd1 vccd1 _15999_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_208_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17738_ _17738_/A vssd1 vssd1 vccd1 vccd1 _22746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_130 _13695_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17669_ _22716_/Q _17556_/X _17671_/S vssd1 vssd1 vccd1 vccd1 _17670_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_141 _20340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19408_ _19408_/A vssd1 vssd1 vccd1 vccd1 _23363_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_152 _15080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_357_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_163 _13974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_174 _17029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20680_ _20680_/A _21301_/C vssd1 vssd1 vccd1 vccd1 _20683_/B sky130_fd_sc_hd__and2_2
XFILLER_126_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_185 _13889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_196 _13945_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19339_ _19555_/B _19483_/B vssd1 vssd1 vccd1 vccd1 _19396_/A sky130_fd_sc_hd__nor2_8
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22350_ _23070_/CLK _22350_/D vssd1 vssd1 vccd1 vccd1 _22350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_338_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21301_ _23781_/Q _21301_/B _21301_/C _21301_/D vssd1 vssd1 vccd1 vccd1 _21301_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22281_ _23515_/CLK _22281_/D vssd1 vssd1 vccd1 vccd1 _22281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_276_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21232_ _14538_/X _21229_/X _21231_/Y _21218_/X vssd1 vssd1 vccd1 vccd1 _23889_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21163_ _21163_/A vssd1 vssd1 vccd1 vccd1 _21163_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_278_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20114_ _20120_/A _20114_/B _20119_/A vssd1 vssd1 vccd1 vccd1 _23644_/D sky130_fd_sc_hd__nor3_1
XFILLER_259_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21094_ _21097_/A _20890_/B _21158_/A vssd1 vssd1 vccd1 vccd1 _21161_/A sky130_fd_sc_hd__o21a_2
XFILLER_302_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20045_ _20121_/A vssd1 vssd1 vccd1 vccd1 _20086_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_274_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_286_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1_2_wb_clk_i clkbuf_1_1_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23804_ _23804_/CLK _23804_/D vssd1 vssd1 vccd1 vccd1 _23804_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21996_ _23835_/Q _21995_/Y _22214_/S vssd1 vssd1 vccd1 vccd1 _21997_/B sky130_fd_sc_hd__mux2_1
XFILLER_54_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23735_ _23918_/CLK _23735_/D vssd1 vssd1 vccd1 vccd1 _23735_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20947_ _17180_/X _20936_/X _20689_/B _20940_/X vssd1 vssd1 vccd1 vccd1 _20947_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_324_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11680_/A vssd1 vssd1 vccd1 vccd1 _11681_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23666_ _23684_/CLK _23666_/D vssd1 vssd1 vccd1 vccd1 _23666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20878_ _20752_/B _20864_/X _20865_/X _23777_/Q vssd1 vssd1 vccd1 vccd1 _20879_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_328_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22617_ _23368_/CLK _22617_/D vssd1 vssd1 vccd1 vccd1 _22617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23597_ _23600_/CLK _23597_/D vssd1 vssd1 vccd1 vccd1 _23597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13350_ _13350_/A _13350_/B vssd1 vssd1 vccd1 vccd1 _15580_/A sky130_fd_sc_hd__nor2_1
X_22548_ _23264_/CLK _22548_/D vssd1 vssd1 vccd1 vccd1 _22548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12301_ _12291_/Y _12294_/Y _12298_/Y _12300_/Y _11214_/A vssd1 vssd1 vccd1 vccd1
+ _12311_/B sky130_fd_sc_hd__o221a_1
XFILLER_344_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13281_ _23489_/Q _23585_/Q _22549_/Q _22353_/Q _13275_/X _13276_/X vssd1 vssd1 vccd1
+ vccd1 _13282_/B sky130_fd_sc_hd__mux4_1
X_22479_ _23070_/CLK _22479_/D vssd1 vssd1 vccd1 vccd1 _22479_/Q sky130_fd_sc_hd__dfxtp_1
X_15020_ _15293_/A _15019_/X _15020_/S vssd1 vssd1 vccd1 vccd1 _15995_/B sky130_fd_sc_hd__mux2_1
X_12232_ _12235_/B vssd1 vssd1 vccd1 vccd1 _12233_/B sky130_fd_sc_hd__clkinv_2
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12163_ _12163_/A vssd1 vssd1 vccd1 vccd1 _12163_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_351_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_296_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_351_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_311_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11114_ _23901_/Q vssd1 vssd1 vccd1 vccd1 _12465_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_312_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16971_ _17382_/A _16971_/B vssd1 vssd1 vccd1 vccd1 _17082_/A sky130_fd_sc_hd__or2_1
X_12094_ _12094_/A vssd1 vssd1 vccd1 vccd1 _12094_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_111_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18710_ _18767_/S vssd1 vssd1 vccd1 vccd1 _18719_/S sky130_fd_sc_hd__buf_6
XFILLER_277_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15922_ _14215_/A _21267_/A _15921_/X _11099_/A vssd1 vssd1 vccd1 vccd1 _15923_/B
+ sky130_fd_sc_hd__o22a_1
X_19690_ _19690_/A vssd1 vssd1 vccd1 vccd1 _23488_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18641_ _23051_/Q _17566_/X _18647_/S vssd1 vssd1 vccd1 vccd1 _18642_/A sky130_fd_sc_hd__mux2_1
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15853_ _15964_/A _15846_/Y _15852_/X vssd1 vssd1 vccd1 vccd1 _15853_/Y sky130_fd_sc_hd__o21ai_1
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14804_ _14804_/A _14804_/B vssd1 vssd1 vccd1 vccd1 _14804_/Y sky130_fd_sc_hd__nor2_1
XFILLER_292_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18572_ _18572_/A vssd1 vssd1 vccd1 vccd1 _23020_/D sky130_fd_sc_hd__clkbuf_1
X_15784_ _18836_/A vssd1 vssd1 vccd1 vccd1 _19229_/A sky130_fd_sc_hd__buf_4
X_12996_ _23323_/Q _23291_/Q _23259_/Q _23547_/Q _12733_/X _12734_/X vssd1 vssd1 vccd1
+ vccd1 _12996_/X sky130_fd_sc_hd__mux4_2
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17523_ _22668_/Q _16278_/X _17527_/S vssd1 vssd1 vccd1 vccd1 _17524_/A sky130_fd_sc_hd__mux2_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14735_ _23591_/Q _14732_/X _14734_/X _23623_/Q vssd1 vssd1 vccd1 vccd1 _14735_/X
+ sky130_fd_sc_hd__o22a_2
X_11947_ _11957_/A vssd1 vssd1 vccd1 vccd1 _12754_/A sky130_fd_sc_hd__buf_2
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ _22638_/Q _16284_/X _17454_/S vssd1 vssd1 vccd1 vccd1 _17455_/A sky130_fd_sc_hd__mux2_1
X_14666_ _14662_/X _15017_/A _15132_/S vssd1 vssd1 vccd1 vccd1 _14667_/A sky130_fd_sc_hd__mux2_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11878_ _22463_/Q _22623_/Q _22302_/Q _23438_/Q _11799_/A _12269_/A vssd1 vssd1 vccd1
+ vccd1 _11879_/B sky130_fd_sc_hd__mux4_1
XFILLER_205_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13617_ _13594_/A _13615_/Y _13603_/A _21790_/A vssd1 vssd1 vccd1 vccd1 _13964_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_16405_ _15240_/X _22365_/Q _16407_/S vssd1 vssd1 vccd1 vccd1 _16406_/A sky130_fd_sc_hd__mux2_1
X_17385_ _18159_/A _17385_/B vssd1 vssd1 vccd1 vccd1 _17386_/A sky130_fd_sc_hd__and2_1
XFILLER_220_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14597_ _16137_/B vssd1 vssd1 vccd1 vccd1 _16102_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_186_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_347_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19124_ _23251_/Q _18817_/X _19124_/S vssd1 vssd1 vccd1 vccd1 _19125_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16336_ _15324_/X _22335_/Q _16344_/S vssd1 vssd1 vccd1 vccd1 _16337_/A sky130_fd_sc_hd__mux2_1
X_13548_ _13548_/A _13548_/B vssd1 vssd1 vccd1 vccd1 _13549_/B sky130_fd_sc_hd__xnor2_4
XFILLER_346_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_319_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_307_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19055_ _19055_/A vssd1 vssd1 vccd1 vccd1 _23220_/D sky130_fd_sc_hd__clkbuf_1
X_16267_ _16267_/A vssd1 vssd1 vccd1 vccd1 _22311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_346_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13479_ _11106_/A _13884_/B _13831_/B _13890_/A vssd1 vssd1 vccd1 vccd1 _13479_/X
+ sky130_fd_sc_hd__a31o_2
X_18006_ _22843_/Q _17990_/X _17986_/A _18005_/X _17933_/A vssd1 vssd1 vccd1 vccd1
+ _18006_/X sky130_fd_sc_hd__a221o_1
X_15218_ _23725_/Q _23855_/Q _16022_/S vssd1 vssd1 vccd1 vccd1 _15218_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput304 _23951_/X vssd1 vssd1 vccd1 vccd1 clk1 sky130_fd_sc_hd__clkbuf_1
X_16198_ _16197_/X _22292_/Q _16198_/S vssd1 vssd1 vccd1 vccd1 _16199_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput315 _13973_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[20] sky130_fd_sc_hd__buf_2
Xoutput326 _13917_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[5] sky130_fd_sc_hd__buf_2
Xoutput337 _13770_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[14] sky130_fd_sc_hd__buf_2
XFILLER_113_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ _15652_/A vssd1 vssd1 vccd1 vccd1 _15150_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput348 _13838_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[24] sky130_fd_sc_hd__buf_2
XFILLER_303_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput359 _13723_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19957_ _19981_/A _19957_/B vssd1 vssd1 vccd1 vccd1 _19957_/Y sky130_fd_sc_hd__nor2_1
XFILLER_287_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18908_ _18908_/A vssd1 vssd1 vccd1 vccd1 _23155_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19888_ _19888_/A vssd1 vssd1 vccd1 vccd1 _23576_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18839_ _18839_/A vssd1 vssd1 vccd1 vccd1 _23129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21850_ _21844_/Y _21846_/Y _21848_/Y _21849_/X vssd1 vssd1 vccd1 vccd1 _21876_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_271_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20801_ _20801_/A vssd1 vssd1 vccd1 vccd1 _23755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21781_ _21801_/D _21781_/B vssd1 vssd1 vccd1 vccd1 _21781_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_63_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23520_ _23552_/CLK _23520_/D vssd1 vssd1 vccd1 vccd1 _23520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_282_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20732_ _20732_/A vssd1 vssd1 vccd1 vccd1 _20732_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_51_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_357_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23451_ _23451_/CLK _23451_/D vssd1 vssd1 vccd1 vccd1 _23451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20663_ _13775_/A _20617_/X _20662_/X vssd1 vssd1 vccd1 vccd1 _20663_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22402_ _23570_/CLK _22402_/D vssd1 vssd1 vccd1 vccd1 _22402_/Q sky130_fd_sc_hd__dfxtp_1
X_23382_ _23414_/CLK _23382_/D vssd1 vssd1 vccd1 vccd1 _23382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_353_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20594_ _20768_/A vssd1 vssd1 vccd1 vccd1 _20626_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_164_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_326_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22333_ _23565_/CLK _22333_/D vssd1 vssd1 vccd1 vccd1 _22333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22264_ _23528_/CLK _22264_/D vssd1 vssd1 vccd1 vccd1 _22264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_353_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21215_ _21215_/A _21215_/B vssd1 vssd1 vccd1 vccd1 _21216_/A sky130_fd_sc_hd__and2_1
XFILLER_117_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22195_ _22195_/A _22195_/B _22195_/C vssd1 vssd1 vccd1 vccd1 _22195_/X sky130_fd_sc_hd__or3_1
XFILLER_333_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21146_ _23864_/Q _21139_/X _21145_/X _21073_/X vssd1 vssd1 vccd1 vccd1 _23864_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_330_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21077_ _21077_/A _21077_/B _21077_/C _21077_/D vssd1 vssd1 vccd1 vccd1 _21078_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_101_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20028_ _23620_/Q _20025_/C _20027_/Y vssd1 vssd1 vccd1 vccd1 _23620_/D sky130_fd_sc_hd__o21a_1
XFILLER_258_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12850_ _23324_/Q _23292_/Q _23260_/Q _23548_/Q _12843_/X _12844_/X vssd1 vssd1 vccd1
+ vccd1 _12850_/X sky130_fd_sc_hd__mux4_2
XFILLER_262_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _22367_/Q _22399_/Q _22688_/Q _23055_/Q _11799_/X _11800_/X vssd1 vssd1 vccd1
+ vccd1 _11802_/B sky130_fd_sc_hd__mux4_1
XFILLER_262_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _23479_/Q _23575_/Q _22539_/Q _22343_/Q _11308_/A _11320_/A vssd1 vssd1 vccd1
+ vccd1 _12781_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21979_ _21979_/A _22032_/B vssd1 vssd1 vccd1 vccd1 _21979_/Y sky130_fd_sc_hd__nor2_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14520_/A _14520_/B vssd1 vssd1 vccd1 vccd1 _14521_/C sky130_fd_sc_hd__nor2_1
XFILLER_242_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23718_ _23851_/CLK _23718_/D vssd1 vssd1 vccd1 vccd1 _23718_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _12269_/A vssd1 vssd1 vccd1 vccd1 _11733_/A sky130_fd_sc_hd__buf_4
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14465_/B _14451_/B _14465_/A vssd1 vssd1 vccd1 vccd1 _14510_/B sky130_fd_sc_hd__or3b_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23649_ _23649_/CLK _23649_/D vssd1 vssd1 vccd1 vccd1 _23649_/Q sky130_fd_sc_hd__dfxtp_1
X_11663_ _12141_/A vssd1 vssd1 vccd1 vccd1 _12909_/A sky130_fd_sc_hd__buf_2
XFILLER_168_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_357_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13402_ _13402_/A _13402_/B vssd1 vssd1 vccd1 vccd1 _13404_/A sky130_fd_sc_hd__xnor2_1
XFILLER_328_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17170_ _23478_/Q _17170_/B vssd1 vssd1 vccd1 vccd1 _17170_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14382_ _15387_/S _14380_/Y _15253_/A vssd1 vssd1 vccd1 vccd1 _14382_/X sky130_fd_sc_hd__a21o_1
XFILLER_328_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11594_ _11594_/A _11594_/B vssd1 vssd1 vccd1 vccd1 _11594_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16121_ _22219_/B vssd1 vssd1 vccd1 vccd1 _22197_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_128_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13333_ _13510_/A _13333_/B vssd1 vssd1 vccd1 vccd1 _13371_/B sky130_fd_sc_hd__or2_1
XFILLER_343_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_332_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16052_ _15633_/X _15380_/Y _15942_/A vssd1 vssd1 vccd1 vccd1 _21276_/A sky130_fd_sc_hd__a21oi_4
X_13264_ _13268_/A _13264_/B vssd1 vssd1 vccd1 vccd1 _13264_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15003_ _15003_/A vssd1 vssd1 vccd1 vccd1 _15003_/X sky130_fd_sc_hd__buf_4
XFILLER_331_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_307_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12215_ _12475_/A vssd1 vssd1 vccd1 vccd1 _12215_/X sky130_fd_sc_hd__buf_4
XFILLER_343_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13195_ _13195_/A vssd1 vssd1 vccd1 vccd1 _13195_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19811_ _23542_/Q _19220_/A _19815_/S vssd1 vssd1 vccd1 vccd1 _19812_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12146_ _11285_/A _12139_/X _12141_/X _12145_/X _11657_/A vssd1 vssd1 vccd1 vccd1
+ _12156_/B sky130_fd_sc_hd__a311o_1
XFILLER_155_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_312_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_296_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19742_ _19742_/A vssd1 vssd1 vccd1 vccd1 _23511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_284_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16954_ _17145_/B vssd1 vssd1 vccd1 vccd1 _17231_/A sky130_fd_sc_hd__buf_2
X_12077_ _23314_/Q _23282_/Q _23250_/Q _23538_/Q _11700_/X _11839_/A vssd1 vssd1 vccd1
+ vccd1 _12078_/B sky130_fd_sc_hd__mux4_1
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15905_ _23677_/Q _15905_/B vssd1 vssd1 vccd1 vccd1 _15905_/X sky130_fd_sc_hd__or2_1
X_19673_ _19684_/A vssd1 vssd1 vccd1 vccd1 _19682_/S sky130_fd_sc_hd__buf_2
XFILLER_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16885_ _16885_/A vssd1 vssd1 vccd1 vccd1 _22542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18624_ _18624_/A vssd1 vssd1 vccd1 vccd1 _23044_/D sky130_fd_sc_hd__clkbuf_1
X_15836_ _23611_/Q _15589_/X _15590_/X _23643_/Q vssd1 vssd1 vccd1 vccd1 _15836_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_266_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18555_ _18623_/S vssd1 vssd1 vccd1 vccd1 _18564_/S sky130_fd_sc_hd__buf_6
X_12979_ _11587_/A _12978_/X _12759_/A vssd1 vssd1 vccd1 vccd1 _12979_/X sky130_fd_sc_hd__a21o_1
X_15767_ _15558_/X _15755_/X _15764_/X _15766_/X _14755_/A vssd1 vssd1 vccd1 vccd1
+ _15767_/X sky130_fd_sc_hd__o32a_4
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17506_ _17506_/A vssd1 vssd1 vccd1 vccd1 _22660_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14718_ _22505_/Q _13691_/A _13888_/B _14717_/X vssd1 vssd1 vccd1 vccd1 _15286_/A
+ sky130_fd_sc_hd__o211ai_2
X_18486_ _22990_/Q _18492_/B vssd1 vssd1 vccd1 vccd1 _18486_/Y sky130_fd_sc_hd__nand2_1
XFILLER_205_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15698_ _15698_/A vssd1 vssd1 vccd1 vccd1 _16188_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_339_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17437_ _22630_/Q _16259_/X _17443_/S vssd1 vssd1 vccd1 vccd1 _17438_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14649_ _14645_/X _14648_/X _15085_/S vssd1 vssd1 vccd1 vccd1 _14649_/X sky130_fd_sc_hd__mux2_2
XFILLER_268_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_348_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17368_ _17368_/A vssd1 vssd1 vccd1 vccd1 _22604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19107_ _23243_/Q _18792_/X _19113_/S vssd1 vssd1 vccd1 vccd1 _19108_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16319_ _16319_/A vssd1 vssd1 vccd1 vccd1 _22327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_347_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17299_ _23490_/Q _17016_/X _17017_/X _17268_/X _17298_/Y vssd1 vssd1 vccd1 vccd1
+ _17299_/X sky130_fd_sc_hd__a32o_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_307_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19038_ _16841_/X _23213_/Q _19040_/S vssd1 vssd1 vccd1 vccd1 _19039_/A sky130_fd_sc_hd__mux2_1
XFILLER_322_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_316_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21000_ _23815_/Q _21009_/B vssd1 vssd1 vccd1 vccd1 _21000_/X sky130_fd_sc_hd__or2_1
XFILLER_303_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_331_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22951_ _23602_/CLK _22951_/D vssd1 vssd1 vccd1 vccd1 _22951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_290_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21902_ _21900_/X _21901_/X _22048_/A vssd1 vssd1 vccd1 vccd1 _21902_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22882_ _23327_/CLK _22882_/D vssd1 vssd1 vccd1 vccd1 _22882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21833_ _21821_/A _21821_/B _21819_/A vssd1 vssd1 vccd1 vccd1 _21837_/A sky130_fd_sc_hd__o21ai_1
XFILLER_37_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_37_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23450_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_243_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21764_ _21740_/A _21739_/B _21739_/A vssd1 vssd1 vccd1 vccd1 _21765_/B sky130_fd_sc_hd__a21bo_1
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23503_ _23503_/CLK _23503_/D vssd1 vssd1 vccd1 vccd1 _23503_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20715_ _17224_/A _20701_/X _20714_/Y vssd1 vssd1 vccd1 vccd1 _20716_/C sky130_fd_sc_hd__a21oi_2
XFILLER_357_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21695_ _21693_/X _21690_/C _21694_/Y _21689_/C vssd1 vssd1 vccd1 vccd1 _21803_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_12_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23434_ _23530_/CLK _23434_/D vssd1 vssd1 vccd1 vccd1 _23434_/Q sky130_fd_sc_hd__dfxtp_1
X_20646_ _23728_/Q _20628_/X _20645_/X _20637_/X vssd1 vssd1 vccd1 vccd1 _23728_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_326_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_326_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_325_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23365_ _23525_/CLK _23365_/D vssd1 vssd1 vccd1 vccd1 _23365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_326_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20577_ _20591_/A _20577_/B _20577_/C vssd1 vssd1 vccd1 vccd1 _20577_/X sky130_fd_sc_hd__or3_1
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_353_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22316_ _23580_/CLK _22316_/D vssd1 vssd1 vccd1 vccd1 _22316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23296_ _23552_/CLK _23296_/D vssd1 vssd1 vccd1 vccd1 _23296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_340_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_298_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22247_ _16936_/C _21321_/A _21295_/B _22712_/Q vssd1 vssd1 vccd1 vccd1 _22247_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_340_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_344_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12000_ _12900_/A _11999_/X _11681_/X vssd1 vssd1 vccd1 vccd1 _12000_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_322_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22178_ _20387_/A _22045_/X _16115_/B _21842_/X vssd1 vssd1 vccd1 vccd1 _22178_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_79_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21129_ _23859_/Q _21123_/X _21124_/X _21025_/A vssd1 vssd1 vccd1 vccd1 _21130_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_238_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_294_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13951_ _13951_/A _13951_/B vssd1 vssd1 vccd1 vccd1 _13951_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12902_ _12707_/X _12895_/X _12897_/X _12901_/X vssd1 vssd1 vccd1 vccd1 _12902_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_247_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16670_ _16670_/A vssd1 vssd1 vccd1 vccd1 _22481_/D sky130_fd_sc_hd__clkbuf_1
X_13882_ _13882_/A _15112_/A vssd1 vssd1 vccd1 vccd1 _14074_/D sky130_fd_sc_hd__or2_4
XFILLER_46_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12833_ _23484_/Q _23580_/Q _22544_/Q _22348_/Q _12692_/X _12041_/X vssd1 vssd1 vccd1
+ vccd1 _12833_/X sky130_fd_sc_hd__mux4_1
X_15621_ _15621_/A vssd1 vssd1 vccd1 vccd1 _15781_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _15950_/X _18341_/C _22940_/Q vssd1 vssd1 vccd1 vccd1 _18342_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _23319_/Q _23287_/Q _23255_/Q _23543_/Q _12922_/S _12746_/X vssd1 vssd1 vccd1
+ vccd1 _12765_/B sky130_fd_sc_hd__mux4_2
XFILLER_226_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _23796_/Q _15219_/A _14606_/A vssd1 vssd1 vccd1 vccd1 _15552_/X sky130_fd_sc_hd__a21o_1
XFILLER_187_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14503_ _15501_/B vssd1 vssd1 vccd1 vccd1 _15835_/B sky130_fd_sc_hd__clkbuf_2
X_11715_ _11698_/Y _11707_/Y _11711_/Y _11714_/Y _11215_/A vssd1 vssd1 vccd1 vccd1
+ _11727_/B sky130_fd_sc_hd__o221a_1
XFILLER_188_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18271_ _18275_/A _18275_/C _18270_/Y vssd1 vssd1 vccd1 vccd1 _22918_/D sky130_fd_sc_hd__o21a_1
X_15483_ _15483_/A _15483_/B vssd1 vssd1 vccd1 vccd1 _15483_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_348_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12695_ _12983_/A vssd1 vssd1 vccd1 vccd1 _12968_/A sky130_fd_sc_hd__buf_2
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17222_ _21077_/B _17222_/B vssd1 vssd1 vccd1 vccd1 _17222_/Y sky130_fd_sc_hd__nor2_1
X_14434_ _14465_/A _14434_/B vssd1 vssd1 vccd1 vccd1 _14506_/B sky130_fd_sc_hd__or2_1
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11646_ _11646_/A vssd1 vssd1 vccd1 vccd1 _11647_/A sky130_fd_sc_hd__buf_6
XFILLER_187_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 core_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_2
X_17153_ _17070_/A _17143_/X _17152_/X _17109_/X vssd1 vssd1 vccd1 vccd1 _17153_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput25 core_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_2
X_14365_ _15385_/S vssd1 vssd1 vccd1 vccd1 _15249_/S sky130_fd_sc_hd__clkbuf_2
X_11577_ _12983_/A _11576_/X _11232_/A vssd1 vssd1 vccd1 vccd1 _11577_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput36 core_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_345_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput47 dout0[13] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_2
XFILLER_318_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16104_ _23810_/Q _14742_/X _15067_/X vssd1 vssd1 vccd1 vccd1 _16104_/X sky130_fd_sc_hd__a21o_1
X_13316_ _13316_/A _13316_/B vssd1 vssd1 vccd1 vccd1 _13317_/B sky130_fd_sc_hd__nand2_1
Xinput58 dout0[23] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_2
XFILLER_183_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17084_ input78/X input106/X _17084_/S vssd1 vssd1 vccd1 vccd1 _17084_/X sky130_fd_sc_hd__mux2_8
Xinput69 dout0[33] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_1
XFILLER_305_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14296_ _14280_/X _14293_/X _15129_/S vssd1 vssd1 vccd1 vccd1 _14296_/X sky130_fd_sc_hd__mux2_2
XFILLER_289_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_304_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13247_ _13402_/A _13244_/X _13246_/Y vssd1 vssd1 vccd1 vccd1 _13247_/Y sky130_fd_sc_hd__a21oi_1
X_16035_ _15338_/A _14956_/X _16033_/Y _16034_/X vssd1 vssd1 vccd1 vccd1 _16035_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_331_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_331_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_297_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13178_ _13117_/A _13177_/X _12745_/X vssd1 vssd1 vccd1 vccd1 _13178_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_313_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12129_ _22273_/Q _23089_/Q _23505_/Q _22434_/Q _11561_/A _11568_/A vssd1 vssd1 vccd1
+ vccd1 _12130_/B sky130_fd_sc_hd__mux4_1
XFILLER_111_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17986_ _17986_/A vssd1 vssd1 vccd1 vccd1 _17986_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19725_ _19725_/A vssd1 vssd1 vccd1 vccd1 _23503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_300_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16937_ _16937_/A _22246_/A _16942_/C _21320_/A vssd1 vssd1 vccd1 vccd1 _16938_/D
+ sky130_fd_sc_hd__or4b_1
XFILLER_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_300_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19656_ _19204_/X _23473_/Q _19660_/S vssd1 vssd1 vccd1 vccd1 _19657_/A sky130_fd_sc_hd__mux2_1
X_16868_ _16867_/X _22537_/Q _16877_/S vssd1 vssd1 vccd1 vccd1 _16869_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18607_ _18607_/A vssd1 vssd1 vccd1 vccd1 _23036_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15819_ _15480_/X _13605_/Y _15663_/X vssd1 vssd1 vccd1 vccd1 _15819_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_350_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19587_ _19587_/A vssd1 vssd1 vccd1 vccd1 _23442_/D sky130_fd_sc_hd__clkbuf_1
X_16799_ _16799_/A vssd1 vssd1 vccd1 vccd1 _22516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18538_ _14700_/C _18537_/Y _18203_/B vssd1 vssd1 vccd1 vccd1 _18538_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_234_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18469_ _22983_/Q _18478_/B vssd1 vssd1 vccd1 vccd1 _18469_/Y sky130_fd_sc_hd__nand2_1
XFILLER_178_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20500_ _20500_/A _20500_/B vssd1 vssd1 vccd1 vccd1 _21313_/B sky130_fd_sc_hd__xor2_2
XFILLER_327_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21480_ _21526_/A _15051_/Y _21480_/S vssd1 vssd1 vccd1 vccd1 _21480_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_348_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20431_ _20491_/B vssd1 vssd1 vccd1 vccd1 _20463_/B sky130_fd_sc_hd__buf_2
XFILLER_335_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_155_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23824_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_295_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23150_ _23502_/CLK _23150_/D vssd1 vssd1 vccd1 vccd1 _23150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20362_ _20362_/A _20387_/B vssd1 vssd1 vccd1 vccd1 _20364_/B sky130_fd_sc_hd__or2_1
XFILLER_335_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22101_ _22101_/A _22101_/B vssd1 vssd1 vccd1 vccd1 _22155_/C sky130_fd_sc_hd__nor2_1
XTAP_7009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23081_ _23560_/CLK _23081_/D vssd1 vssd1 vccd1 vccd1 _23081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20293_ _23668_/Q _20165_/X _20292_/Y _20285_/X vssd1 vssd1 vccd1 vccd1 _23668_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_6308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_288_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22032_ _22032_/A _22032_/B vssd1 vssd1 vccd1 vccd1 _22032_/Y sky130_fd_sc_hd__nor2_1
XFILLER_310_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_304_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_303_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_291_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22934_ _22947_/CLK _22934_/D vssd1 vssd1 vccd1 vccd1 _22934_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_272_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22865_ _23599_/CLK _22865_/D vssd1 vssd1 vccd1 vccd1 _22865_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_243_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21816_ _21816_/A vssd1 vssd1 vccd1 vccd1 _22242_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_271_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22796_ _23450_/CLK _22796_/D vssd1 vssd1 vccd1 vccd1 _22796_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21747_ _14675_/A _21556_/X _21849_/A vssd1 vssd1 vccd1 vccd1 _21779_/A sky130_fd_sc_hd__o21a_2
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11500_ _11236_/A _11491_/Y _11495_/Y _11497_/Y _11499_/Y vssd1 vssd1 vccd1 vccd1
+ _11500_/X sky130_fd_sc_hd__o32a_1
XPHY_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12480_ _12485_/A _12480_/B vssd1 vssd1 vccd1 vccd1 _12480_/X sky130_fd_sc_hd__or2_1
XFILLER_184_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21678_ _22197_/B _21675_/Y _21676_/Y _21677_/X vssd1 vssd1 vccd1 vccd1 _21679_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_339_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23417_ _23419_/CLK _23417_/D vssd1 vssd1 vccd1 vccd1 _23417_/Q sky130_fd_sc_hd__dfxtp_1
X_11431_ _11431_/A vssd1 vssd1 vccd1 vccd1 _11432_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20629_ _20768_/A vssd1 vssd1 vccd1 vccd1 _20665_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_295_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14150_ _14159_/A _16917_/A vssd1 vssd1 vccd1 vccd1 _14161_/A sky130_fd_sc_hd__nor2_1
X_23348_ _23414_/CLK _23348_/D vssd1 vssd1 vccd1 vccd1 _23348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_299_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11362_ _12864_/A vssd1 vssd1 vccd1 vccd1 _13184_/A sky130_fd_sc_hd__buf_6
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13101_ _13107_/A _13101_/B vssd1 vssd1 vccd1 vccd1 _13101_/Y sky130_fd_sc_hd__nor2_1
XFILLER_299_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14081_ _14081_/A vssd1 vssd1 vccd1 vccd1 _14081_/X sky130_fd_sc_hd__buf_2
XFILLER_164_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23279_ _23535_/CLK _23279_/D vssd1 vssd1 vccd1 vccd1 _23279_/Q sky130_fd_sc_hd__dfxtp_1
X_11293_ _12316_/A vssd1 vssd1 vccd1 vccd1 _11914_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_342_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13032_ _22481_/Q _22641_/Q _13032_/S vssd1 vssd1 vccd1 vccd1 _13032_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_313_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17840_ _22792_/Q _17594_/X _17848_/S vssd1 vssd1 vccd1 vccd1 _17841_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17771_ _17771_/A vssd1 vssd1 vccd1 vccd1 _22761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14983_ _18785_/A vssd1 vssd1 vccd1 vccd1 _19178_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_281_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_304_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19510_ _19201_/X _23408_/Q _19516_/S vssd1 vssd1 vccd1 vccd1 _19511_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16722_ _22495_/Q _16711_/X _16712_/X input40/X vssd1 vssd1 vccd1 vccd1 _16723_/B
+ sky130_fd_sc_hd__o22a_1
X_13934_ _13934_/A vssd1 vssd1 vccd1 vccd1 _16679_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_281_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19441_ _19441_/A vssd1 vssd1 vccd1 vccd1 _23377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16653_ _16664_/A vssd1 vssd1 vccd1 vccd1 _16662_/S sky130_fd_sc_hd__buf_2
X_13865_ _11511_/B _13798_/B _13709_/A vssd1 vssd1 vccd1 vccd1 _13865_/X sky130_fd_sc_hd__a21o_1
XFILLER_62_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_504 _18792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_515 _23464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15604_ _22962_/Q _15603_/X _16109_/A vssd1 vssd1 vccd1 vccd1 _15604_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_526 _14017_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12816_ _12816_/A vssd1 vssd1 vccd1 vccd1 _12816_/X sky130_fd_sc_hd__buf_4
X_19372_ _23347_/Q _18817_/X _19372_/S vssd1 vssd1 vccd1 vccd1 _19373_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_537 _23911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_343_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16584_ _15823_/X _22443_/Q _16590_/S vssd1 vssd1 vccd1 vccd1 _16585_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_548 _20305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13796_ _13969_/A vssd1 vssd1 vccd1 vccd1 _13855_/A sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_559 _23879_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18323_ _22933_/Q _22934_/Q _18323_/C vssd1 vssd1 vccd1 vccd1 _18326_/B sky130_fd_sc_hd__and3_1
XFILLER_16_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15535_ _15113_/B _15181_/X _15183_/X _15534_/Y vssd1 vssd1 vccd1 vccd1 _21244_/A
+ sky130_fd_sc_hd__a22o_4
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_349_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12747_ _22795_/Q _22763_/Q _22664_/Q _22731_/Q _12920_/A _12746_/X vssd1 vssd1 vccd1
+ vccd1 _12748_/B sky130_fd_sc_hd__mux4_1
XFILLER_249_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ _22865_/Q _18242_/X _18253_/X _18245_/X vssd1 vssd1 vccd1 vccd1 _22913_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_337_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12678_ _13195_/A _12674_/X _12677_/X vssd1 vssd1 vccd1 vccd1 _12678_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_230_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15466_ _20493_/B vssd1 vssd1 vccd1 vccd1 _16154_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_187_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17205_ _21949_/A _17204_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17205_/X sky130_fd_sc_hd__mux2_1
X_14417_ _14447_/A vssd1 vssd1 vccd1 vccd1 _14500_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11629_ _23928_/Q vssd1 vssd1 vccd1 vccd1 _21846_/A sky130_fd_sc_hd__clkinv_8
X_18185_ _18188_/A _18163_/A _18171_/X _18166_/B vssd1 vssd1 vccd1 vccd1 _18186_/B
+ sky130_fd_sc_hd__a31o_1
X_15397_ _19975_/B _14731_/A _14733_/A _23633_/Q vssd1 vssd1 vccd1 vccd1 _15397_/X
+ sky130_fd_sc_hd__o22a_4
X_17136_ _13775_/A _17135_/X _17234_/S vssd1 vssd1 vccd1 vccd1 _17136_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_305_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14348_ _14348_/A vssd1 vssd1 vccd1 vccd1 _14358_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_289_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17067_ _17000_/A _17060_/X _17066_/X _17057_/X vssd1 vssd1 vccd1 vccd1 _17067_/X
+ sky130_fd_sc_hd__o211a_4
X_14279_ _14292_/A vssd1 vssd1 vccd1 vccd1 _14639_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_304_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_289_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16018_ _22941_/Q _15000_/X _15001_/X _22973_/Q vssd1 vssd1 vccd1 vccd1 _16018_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_171_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_313_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_297_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17969_ _22833_/Q _17956_/X _17959_/X input279/X _17966_/X vssd1 vssd1 vccd1 vccd1
+ _17969_/X sky130_fd_sc_hd__a221o_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19708_ _19175_/X _23496_/Q _19710_/S vssd1 vssd1 vccd1 vccd1 _19709_/A sky130_fd_sc_hd__mux2_1
X_20980_ _22193_/A _21085_/A _20757_/B _20970_/X vssd1 vssd1 vccd1 vccd1 _20980_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_168_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19639_ _19639_/A vssd1 vssd1 vccd1 vccd1 _23465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22650_ _23054_/CLK _22650_/D vssd1 vssd1 vccd1 vccd1 _22650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21601_ _21601_/A _21845_/A vssd1 vssd1 vccd1 vccd1 _21601_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22581_ _23643_/CLK _22581_/D vssd1 vssd1 vccd1 vccd1 _22581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21532_ _23820_/Q _23754_/Q vssd1 vssd1 vccd1 vccd1 _21533_/B sky130_fd_sc_hd__nand2_1
XFILLER_167_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21463_ _22025_/A _21463_/B vssd1 vssd1 vccd1 vccd1 _21463_/Y sky130_fd_sc_hd__nand2_1
XFILLER_355_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_324_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23202_ _23489_/CLK _23202_/D vssd1 vssd1 vccd1 vccd1 _23202_/Q sky130_fd_sc_hd__dfxtp_1
X_20414_ _20470_/A vssd1 vssd1 vccd1 vccd1 _20491_/B sky130_fd_sc_hd__buf_4
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21394_ _21613_/A vssd1 vssd1 vccd1 vccd1 _22129_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_335_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23133_ _23549_/CLK _23133_/D vssd1 vssd1 vccd1 vccd1 _23133_/Q sky130_fd_sc_hd__dfxtp_1
X_20345_ _23675_/Q _20391_/B vssd1 vssd1 vccd1 vccd1 _20345_/X sky130_fd_sc_hd__or2_1
XFILLER_108_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_350_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_324_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_350_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23064_ _23450_/CLK _23064_/D vssd1 vssd1 vccd1 vccd1 _23064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20276_ _20187_/X _20274_/Y _20275_/X _21741_/A _20192_/X vssd1 vssd1 vccd1 vccd1
+ _20654_/A sky130_fd_sc_hd__a32o_4
XFILLER_350_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_288_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22015_ _12841_/Y _21867_/X _22014_/X _21865_/X vssd1 vssd1 vccd1 vccd1 _22041_/D
+ sky130_fd_sc_hd__a22oi_4
XFILLER_310_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput204 localMemory_wb_adr_i[22] vssd1 vssd1 vccd1 vccd1 _14148_/C sky130_fd_sc_hd__buf_2
XFILLER_276_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput215 localMemory_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input215/X sky130_fd_sc_hd__buf_4
XTAP_5437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput226 localMemory_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input226/X sky130_fd_sc_hd__buf_4
XTAP_5448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput237 localMemory_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input237/X sky130_fd_sc_hd__buf_4
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23441_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput248 localMemory_wb_sel_i[1] vssd1 vssd1 vccd1 vccd1 input248/X sky130_fd_sc_hd__clkbuf_1
Xinput259 manufacturerID[5] vssd1 vssd1 vccd1 vccd1 input259/X sky130_fd_sc_hd__buf_2
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ _12661_/A _13875_/A vssd1 vssd1 vccd1 vccd1 _11980_/Y sky130_fd_sc_hd__nand2_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22917_ _23599_/CLK _22917_/D vssd1 vssd1 vccd1 vccd1 _22917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23897_ _23903_/CLK _23897_/D vssd1 vssd1 vccd1 vccd1 _23897_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_260_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13650_ _13650_/A vssd1 vssd1 vccd1 vccd1 _13651_/B sky130_fd_sc_hd__clkbuf_16
X_22848_ _23426_/CLK _22848_/D vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XFILLER_231_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _13334_/D vssd1 vssd1 vccd1 vccd1 _13355_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13581_ _13581_/A _13581_/B vssd1 vssd1 vccd1 vccd1 _13581_/Y sky130_fd_sc_hd__nand2_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22779_ _22779_/CLK _22779_/D vssd1 vssd1 vccd1 vccd1 _22779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15320_ _22988_/Q _15416_/A _15417_/A input216/X vssd1 vssd1 vccd1 vccd1 _21641_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_212_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12532_ _12532_/A _12532_/B vssd1 vssd1 vccd1 vccd1 _12532_/Y sky130_fd_sc_hd__nor2_1
XFILLER_240_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_319_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15251_ _15091_/Y _15250_/Y _15341_/S vssd1 vssd1 vccd1 vccd1 _15251_/X sky130_fd_sc_hd__mux2_1
X_12463_ _12463_/A _12463_/B vssd1 vssd1 vccd1 vccd1 _12463_/Y sky130_fd_sc_hd__nor2_1
XFILLER_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14202_ _16530_/A _20533_/C _14202_/C _21289_/B vssd1 vssd1 vccd1 vccd1 _14526_/A
+ sky130_fd_sc_hd__or4_2
X_11414_ _11414_/A vssd1 vssd1 vccd1 vccd1 _11894_/S sky130_fd_sc_hd__buf_6
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15182_ _14725_/A _15901_/B _15180_/A vssd1 vssd1 vccd1 vccd1 _15183_/A sky130_fd_sc_hd__o21a_1
XFILLER_314_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12394_ _12596_/B _21386_/A _12393_/Y vssd1 vssd1 vccd1 vccd1 _13502_/A sky130_fd_sc_hd__o21a_4
XFILLER_327_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_299_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_354_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14133_ _20191_/A _14133_/B _20532_/D vssd1 vssd1 vccd1 vccd1 _14133_/X sky130_fd_sc_hd__or3_2
XFILLER_326_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_315_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11345_ _11678_/A vssd1 vssd1 vccd1 vccd1 _11346_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19990_ _23609_/Q _20003_/C _19989_/Y vssd1 vssd1 vccd1 vccd1 _23609_/D sky130_fd_sc_hd__o21a_1
XFILLER_315_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_298_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_330_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18941_ _18941_/A vssd1 vssd1 vccd1 vccd1 _23170_/D sky130_fd_sc_hd__clkbuf_1
X_14064_ _14064_/A _14066_/B _14064_/C vssd1 vssd1 vccd1 vccd1 _14064_/X sky130_fd_sc_hd__or3_1
XFILLER_140_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11276_ _11276_/A vssd1 vssd1 vccd1 vccd1 _11277_/A sky130_fd_sc_hd__buf_8
XFILLER_125_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_315_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13015_ _13015_/A _13015_/B vssd1 vssd1 vccd1 vccd1 _13492_/D sky130_fd_sc_hd__nor2_1
XFILLER_3_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18872_ _23140_/Q _18871_/X _18872_/S vssd1 vssd1 vccd1 vccd1 _18873_/A sky130_fd_sc_hd__mux2_1
XTAP_7395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17823_ _17823_/A vssd1 vssd1 vccd1 vccd1 _22784_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_310_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_295_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_239_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17754_ _22754_/Q _17575_/X _17754_/S vssd1 vssd1 vccd1 vccd1 _17755_/A sky130_fd_sc_hd__mux2_1
XTAP_5993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14966_ _22507_/Q _14231_/A _13887_/A _14965_/X vssd1 vssd1 vccd1 vccd1 _15381_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_82_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16705_ _16705_/A vssd1 vssd1 vccd1 vccd1 _22490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13917_ _13917_/A vssd1 vssd1 vccd1 vccd1 _13917_/X sky130_fd_sc_hd__clkbuf_1
X_17685_ _22723_/Q _17578_/X _17693_/S vssd1 vssd1 vccd1 vccd1 _17686_/A sky130_fd_sc_hd__mux2_1
X_14897_ _14897_/A vssd1 vssd1 vccd1 vccd1 _14898_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_301 _15990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_312 _16045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19424_ _19481_/S vssd1 vssd1 vccd1 vccd1 _19433_/S sky130_fd_sc_hd__buf_4
XFILLER_235_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_323 _16107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16636_ _22466_/Q _16246_/X _16640_/S vssd1 vssd1 vccd1 vccd1 _16637_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_334 _17067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13848_ _13110_/B _13808_/X _13781_/X vssd1 vssd1 vccd1 vccd1 _13848_/X sky130_fd_sc_hd__a21o_1
XFILLER_90_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_345 _21949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_356 _22116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_367 _23475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19355_ _23339_/Q _18792_/X _19361_/S vssd1 vssd1 vccd1 vccd1 _19356_/A sky130_fd_sc_hd__mux2_1
XFILLER_250_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_378 _22487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16567_ _16567_/A vssd1 vssd1 vccd1 vccd1 _22435_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13779_ _13779_/A _13890_/A _19969_/D vssd1 vssd1 vccd1 vccd1 _13808_/A sky130_fd_sc_hd__and3_1
XFILLER_149_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_389 _16530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18306_ _18315_/A _18306_/B _18306_/C vssd1 vssd1 vccd1 vccd1 _22928_/D sky130_fd_sc_hd__nor3_1
XFILLER_31_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15518_ _15480_/X _15517_/X _14529_/A vssd1 vssd1 vccd1 vccd1 _15518_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_188_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19286_ _19286_/A vssd1 vssd1 vccd1 vccd1 _23308_/D sky130_fd_sc_hd__clkbuf_1
X_16498_ _15668_/X _22406_/Q _16502_/S vssd1 vssd1 vccd1 vccd1 _16499_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18237_ hold8/X _18229_/X _18236_/X _18232_/X vssd1 vssd1 vccd1 vccd1 _22906_/D sky130_fd_sc_hd__o211a_1
X_15449_ _15440_/X _15441_/X _15448_/Y _15150_/A vssd1 vssd1 vccd1 vccd1 _15450_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18168_ _18163_/B _18144_/B _18167_/X _18162_/X vssd1 vssd1 vccd1 vccd1 _18168_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_345_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17119_ _17070_/X _17112_/X _17118_/X _17109_/X vssd1 vssd1 vccd1 vccd1 _17119_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_289_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18099_ _18099_/A vssd1 vssd1 vccd1 vccd1 _18099_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_306_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_332_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_292_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_321_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20130_ _23649_/Q _20127_/C _23650_/Q vssd1 vssd1 vccd1 vccd1 _20132_/B sky130_fd_sc_hd__a21oi_1
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20061_ _23629_/Q _20076_/C _23630_/Q vssd1 vssd1 vccd1 vccd1 _20064_/B sky130_fd_sc_hd__a21oi_1
XFILLER_301_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_297_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_16 _17483_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_27 _17743_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_38 _20058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_300_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23820_ _23824_/CLK _23820_/D vssd1 vssd1 vccd1 vccd1 _23820_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_49 _20966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23751_ _23862_/CLK _23751_/D vssd1 vssd1 vccd1 vccd1 _23751_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_260_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20963_ _20963_/A vssd1 vssd1 vccd1 vccd1 _21023_/A sky130_fd_sc_hd__buf_4
XFILLER_53_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22702_ _23073_/CLK _22702_/D vssd1 vssd1 vccd1 vccd1 _22702_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23682_ _23706_/CLK _23682_/D vssd1 vssd1 vccd1 vccd1 _23682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20894_ _20966_/A vssd1 vssd1 vccd1 vccd1 _20894_/X sky130_fd_sc_hd__buf_2
XFILLER_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22633_ _23448_/CLK _22633_/D vssd1 vssd1 vccd1 vccd1 _22633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_170_wb_clk_i _23917_/CLK vssd1 vssd1 vccd1 vccd1 _23841_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_213_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22564_ _22600_/CLK _22564_/D vssd1 vssd1 vccd1 vccd1 _22564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21515_ _21515_/A _21515_/B vssd1 vssd1 vccd1 vccd1 _21515_/Y sky130_fd_sc_hd__nor2_1
XFILLER_221_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_355_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22495_ _23714_/CLK _22495_/D vssd1 vssd1 vccd1 vccd1 _22495_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_319_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_343_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21446_ _11084_/A _21518_/A _14564_/A vssd1 vssd1 vccd1 vccd1 _21480_/S sky130_fd_sc_hd__a21oi_1
XFILLER_119_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_292_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21377_ _21377_/A vssd1 vssd1 vccd1 vccd1 _21377_/X sky130_fd_sc_hd__buf_4
XFILLER_312_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11130_ _12371_/A vssd1 vssd1 vccd1 vccd1 _11131_/A sky130_fd_sc_hd__clkbuf_4
X_23116_ _23950_/A _23116_/D vssd1 vssd1 vccd1 vccd1 _23116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_296_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20328_ _15767_/X _20169_/X _20329_/B vssd1 vssd1 vccd1 vccd1 _20328_/X sky130_fd_sc_hd__a21o_1
XFILLER_123_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_312_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23047_ _23047_/CLK _23047_/D vssd1 vssd1 vccd1 vccd1 _23047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_311_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20259_ _23664_/Q _20277_/B vssd1 vssd1 vccd1 vccd1 _20259_/X sky130_fd_sc_hd__or2_1
XFILLER_352_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_295_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_297_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_291_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14820_ _14820_/A vssd1 vssd1 vccd1 vccd1 _15698_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14751_ _14729_/X _14749_/X _16109_/A vssd1 vssd1 vccd1 vccd1 _14751_/X sky130_fd_sc_hd__mux2_1
XFILLER_218_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11963_ _12073_/A vssd1 vssd1 vccd1 vccd1 _12756_/A sky130_fd_sc_hd__buf_4
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _13969_/A vssd1 vssd1 vccd1 vccd1 _13728_/B sky130_fd_sc_hd__buf_2
XFILLER_233_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17470_ _17470_/A vssd1 vssd1 vccd1 vccd1 _22645_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _14682_/A vssd1 vssd1 vccd1 vccd1 _14682_/X sky130_fd_sc_hd__clkbuf_4
X_11894_ _22301_/Q _23437_/Q _11894_/S vssd1 vssd1 vccd1 vccd1 _11894_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16421_ _15570_/X _22372_/Q _16429_/S vssd1 vssd1 vccd1 vccd1 _16422_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13633_ _13633_/A _13633_/B vssd1 vssd1 vccd1 vccd1 _13633_/Y sky130_fd_sc_hd__nor2_4
XFILLER_232_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19140_ _23258_/Q _18840_/X _19146_/S vssd1 vssd1 vccd1 vccd1 _19141_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16352_ _16352_/A vssd1 vssd1 vccd1 vccd1 _22342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13564_ _13570_/A vssd1 vssd1 vccd1 vccd1 _13581_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15303_ _23727_/Q _23857_/Q _16022_/S vssd1 vssd1 vccd1 vccd1 _15303_/X sky130_fd_sc_hd__mux2_1
X_19071_ _16889_/X _23228_/Q _19073_/S vssd1 vssd1 vccd1 vccd1 _19072_/A sky130_fd_sc_hd__mux2_1
X_12515_ _23896_/Q _12515_/B vssd1 vssd1 vccd1 vccd1 _12515_/X sky130_fd_sc_hd__or2_2
XFILLER_319_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16283_ _16283_/A vssd1 vssd1 vccd1 vccd1 _22316_/D sky130_fd_sc_hd__clkbuf_1
X_13495_ _13495_/A vssd1 vssd1 vccd1 vccd1 _13495_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18022_ _18099_/A vssd1 vssd1 vccd1 vccd1 _18054_/A sky130_fd_sc_hd__buf_2
XFILLER_306_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12446_ _12463_/A _12446_/B vssd1 vssd1 vccd1 vccd1 _12446_/Y sky130_fd_sc_hd__nor2_1
X_15234_ _15318_/A _15234_/B vssd1 vssd1 vccd1 vccd1 _15234_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_315_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15165_ _22985_/Q _14138_/A _15417_/A input244/X vssd1 vssd1 vccd1 vccd1 _21515_/A
+ sky130_fd_sc_hd__a22o_4
X_12377_ _23304_/Q _23272_/Q _23240_/Q _23528_/Q _12215_/X _12216_/X vssd1 vssd1 vccd1
+ vccd1 _12378_/B sky130_fd_sc_hd__mux4_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_330_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14116_ _22887_/Q vssd1 vssd1 vccd1 vccd1 _14121_/C sky130_fd_sc_hd__inv_2
XFILLER_153_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ _11659_/A vssd1 vssd1 vccd1 vccd1 _12489_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19973_ _23605_/Q _19985_/C _19972_/Y vssd1 vssd1 vccd1 vccd1 _23605_/D sky130_fd_sc_hd__o21a_1
X_15096_ _20138_/B _15078_/X _15079_/Y _15095_/X vssd1 vssd1 vccd1 vccd1 _15096_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_314_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18924_ _18924_/A vssd1 vssd1 vccd1 vccd1 _23162_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_330_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14047_ input225/X _14038_/X _14046_/X vssd1 vssd1 vccd1 vccd1 _14047_/X sky130_fd_sc_hd__a21bo_4
XFILLER_69_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11259_ _12345_/B _14132_/D _11382_/B vssd1 vssd1 vccd1 vccd1 _14371_/A sky130_fd_sc_hd__nand3_2
XFILLER_141_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18855_ _18855_/A vssd1 vssd1 vccd1 vccd1 _23134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_311_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17806_ _17874_/S vssd1 vssd1 vccd1 vccd1 _17815_/S sky130_fd_sc_hd__buf_6
XFILLER_94_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18786_ _23113_/Q _18785_/X _18786_/S vssd1 vssd1 vccd1 vccd1 _18787_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15998_ _13404_/A _13570_/B _16053_/S vssd1 vssd1 vccd1 vccd1 _15998_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17737_ _22746_/Q _17550_/X _17743_/S vssd1 vssd1 vccd1 vccd1 _17738_/A sky130_fd_sc_hd__mux2_1
X_14949_ _14311_/X _14280_/X _14949_/S vssd1 vssd1 vccd1 vccd1 _14949_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17668_ _17668_/A vssd1 vssd1 vccd1 vccd1 _22715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_120 _21444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_131 _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19407_ _23363_/Q _18868_/X _19409_/S vssd1 vssd1 vccd1 vccd1 _19408_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_142 _20374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_153 _13433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16619_ _16619_/A vssd1 vssd1 vccd1 vccd1 _22458_/D sky130_fd_sc_hd__clkbuf_1
X_17599_ _22694_/Q _17598_/X _17608_/S vssd1 vssd1 vccd1 vccd1 _17600_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_164 _21790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_175 _14204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_186 _13889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_356_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19338_ _19338_/A vssd1 vssd1 vccd1 vccd1 _23332_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_197 _13948_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19269_ _19337_/S vssd1 vssd1 vccd1 vccd1 _19278_/S sky130_fd_sc_hd__buf_6
XFILLER_353_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21300_ _21479_/A _21300_/B vssd1 vssd1 vccd1 vccd1 _21300_/X sky130_fd_sc_hd__and2b_1
XFILLER_352_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22280_ _23480_/CLK _22280_/D vssd1 vssd1 vccd1 vccd1 _22280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21231_ _21231_/A _21240_/B vssd1 vssd1 vccd1 vccd1 _21231_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_4_3_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_191_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21162_ _21083_/A _20520_/D _21140_/X _20713_/A _21161_/X vssd1 vssd1 vccd1 vccd1
+ _21162_/X sky130_fd_sc_hd__a221o_1
XFILLER_117_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_305_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20113_ _20126_/C vssd1 vssd1 vccd1 vccd1 _20119_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_236_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21093_ _21093_/A vssd1 vssd1 vccd1 vccd1 _21158_/A sky130_fd_sc_hd__buf_2
XFILLER_132_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20044_ _23625_/Q _20051_/A _20043_/Y vssd1 vssd1 vccd1 vccd1 _23625_/D sky130_fd_sc_hd__o21a_1
XFILLER_219_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_302_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23803_ _23942_/CLK _23803_/D vssd1 vssd1 vccd1 vccd1 _23803_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ _21995_/A _21995_/B vssd1 vssd1 vccd1 vccd1 _21995_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20946_ _23798_/Q _20939_/X _20945_/X _20934_/X vssd1 vssd1 vccd1 vccd1 _23798_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23734_ _23918_/CLK _23734_/D vssd1 vssd1 vccd1 vccd1 _23734_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20877_ _20877_/A vssd1 vssd1 vccd1 vccd1 _23776_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23665_ _23704_/CLK _23665_/D vssd1 vssd1 vccd1 vccd1 _23665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22616_ _23527_/CLK _22616_/D vssd1 vssd1 vccd1 vccd1 _22616_/Q sky130_fd_sc_hd__dfxtp_1
X_23596_ _23637_/CLK _23596_/D vssd1 vssd1 vccd1 vccd1 _23596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22547_ _23582_/CLK _22547_/D vssd1 vssd1 vccd1 vccd1 _22547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_329_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ _12565_/A _12299_/X _11844_/X vssd1 vssd1 vccd1 vccd1 _12300_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_316_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13280_ _13287_/A _13279_/X _11353_/A vssd1 vssd1 vccd1 vccd1 _13280_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_155_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_300_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22478_ _23581_/CLK _22478_/D vssd1 vssd1 vccd1 vccd1 _22478_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_344_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_343_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12231_ _12596_/B _21517_/A _12230_/X vssd1 vssd1 vccd1 vccd1 _12235_/B sky130_fd_sc_hd__o21a_4
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21429_ _22129_/A vssd1 vssd1 vccd1 vccd1 _21813_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_163_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12162_ _13623_/A vssd1 vssd1 vccd1 vccd1 _12162_/Y sky130_fd_sc_hd__inv_2
XFILLER_352_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_297_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11113_ _11113_/A vssd1 vssd1 vccd1 vccd1 _11595_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_312_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16970_ _17000_/A _16926_/X _17109_/A _16969_/X vssd1 vssd1 vccd1 vccd1 _16970_/X
+ sky130_fd_sc_hd__o211a_2
X_12093_ _12105_/A _12093_/B vssd1 vssd1 vccd1 vccd1 _12093_/X sky130_fd_sc_hd__or2_1
XFILLER_110_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15921_ _15815_/A _15914_/X _15920_/X _14690_/X vssd1 vssd1 vccd1 vccd1 _15921_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_104_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18640_ _18640_/A vssd1 vssd1 vccd1 vccd1 _23050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_276_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15852_ _15848_/Y _15849_/X _15851_/X _14801_/A vssd1 vssd1 vccd1 vccd1 _15852_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_77_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14803_ _14215_/X _21206_/A _14802_/X _14521_/A vssd1 vssd1 vccd1 vccd1 _14804_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ _16838_/X _23020_/Q _18575_/S vssd1 vssd1 vccd1 vccd1 _18572_/A sky130_fd_sc_hd__mux2_1
X_15783_ _15779_/X _21954_/A _16047_/S vssd1 vssd1 vccd1 vccd1 _18836_/A sky130_fd_sc_hd__mux2_8
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12995_ _12995_/A _12995_/B vssd1 vssd1 vccd1 vccd1 _12995_/X sky130_fd_sc_hd__or2_1
XFILLER_252_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _17522_/A vssd1 vssd1 vccd1 vccd1 _22667_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14734_ _14902_/A vssd1 vssd1 vccd1 vccd1 _14734_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ _13343_/B _11943_/Y _11945_/X vssd1 vssd1 vccd1 vccd1 _11946_/X sky130_fd_sc_hd__o21a_2
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ _17453_/A vssd1 vssd1 vccd1 vccd1 _22637_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14665_ _14663_/X _14664_/X _14665_/S vssd1 vssd1 vccd1 vccd1 _15017_/A sky130_fd_sc_hd__mux2_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11877_ _12321_/A vssd1 vssd1 vccd1 vccd1 _12586_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_338_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16404_ _16404_/A vssd1 vssd1 vccd1 vccd1 _22364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13616_ _13616_/A vssd1 vssd1 vccd1 vccd1 _21790_/A sky130_fd_sc_hd__buf_8
X_17384_ _20790_/A vssd1 vssd1 vccd1 vccd1 _18159_/A sky130_fd_sc_hd__clkbuf_2
X_14596_ _16170_/B vssd1 vssd1 vccd1 vccd1 _16137_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_220_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19123_ _19123_/A vssd1 vssd1 vccd1 vccd1 _23250_/D sky130_fd_sc_hd__clkbuf_1
X_16335_ _16381_/S vssd1 vssd1 vccd1 vccd1 _16344_/S sky130_fd_sc_hd__buf_4
XFILLER_125_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13547_ _13403_/B _13565_/B _16054_/A vssd1 vssd1 vccd1 vccd1 _13548_/B sky130_fd_sc_hd__a21oi_2
XFILLER_347_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_346_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_346_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19054_ _16863_/X _23220_/Q _19062_/S vssd1 vssd1 vccd1 vccd1 _19055_/A sky130_fd_sc_hd__mux2_1
XFILLER_307_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16266_ _22311_/Q _16265_/X _16269_/S vssd1 vssd1 vccd1 vccd1 _16267_/A sky130_fd_sc_hd__mux2_1
X_13478_ _13367_/C _13467_/A _13474_/A _23911_/Q vssd1 vssd1 vccd1 vccd1 _13831_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18005_ input8/X input283/X _18005_/S vssd1 vssd1 vccd1 vccd1 _18005_/X sky130_fd_sc_hd__mux2_1
XFILLER_346_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15217_ _15806_/S vssd1 vssd1 vccd1 vccd1 _16022_/S sky130_fd_sc_hd__buf_4
X_12429_ _11844_/A _12419_/Y _12421_/Y _12428_/X _11240_/A vssd1 vssd1 vccd1 vccd1
+ _12439_/B sky130_fd_sc_hd__o311a_1
X_16197_ _19264_/A vssd1 vssd1 vccd1 vccd1 _16197_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput305 _13953_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[10] sky130_fd_sc_hd__buf_2
XFILLER_127_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput316 _13974_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[21] sky130_fd_sc_hd__buf_2
XFILLER_315_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput327 _13926_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[6] sky130_fd_sc_hd__buf_2
X_15148_ _15148_/A _15148_/B vssd1 vssd1 vccd1 vccd1 _15652_/A sky130_fd_sc_hd__nand2_2
XFILLER_154_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput338 _13773_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[15] sky130_fd_sc_hd__buf_2
XFILLER_126_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput349 _13845_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[25] sky130_fd_sc_hd__buf_2
XFILLER_259_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_303_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19956_ _19975_/B _19959_/C vssd1 vssd1 vccd1 vccd1 _19957_/B sky130_fd_sc_hd__and2_1
X_15079_ _15079_/A _15079_/B vssd1 vssd1 vccd1 vccd1 _15079_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18907_ _23155_/Q _18817_/X _18907_/S vssd1 vssd1 vccd1 vccd1 _18908_/A sky130_fd_sc_hd__mux2_1
XFILLER_296_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19887_ _16268_/X _23576_/Q _19887_/S vssd1 vssd1 vccd1 vccd1 _19888_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18838_ _23129_/Q _18836_/X _18850_/S vssd1 vssd1 vccd1 vccd1 _18839_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_109_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _22822_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_67_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_347_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18769_ _18769_/A vssd1 vssd1 vccd1 vccd1 _18769_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_282_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20800_ _20806_/A _20800_/B vssd1 vssd1 vccd1 vccd1 _20801_/A sky130_fd_sc_hd__and2_1
X_21780_ _21801_/C _21752_/B _21799_/A vssd1 vssd1 vccd1 vccd1 _21781_/B sky130_fd_sc_hd__a21bo_1
XFILLER_298_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20731_ _20731_/A _20731_/B vssd1 vssd1 vccd1 vccd1 _20736_/B sky130_fd_sc_hd__and2_1
XFILLER_169_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23450_ _23450_/CLK _23450_/D vssd1 vssd1 vccd1 vccd1 _23450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_357_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20662_ _20662_/A vssd1 vssd1 vccd1 vccd1 _20662_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22401_ _23571_/CLK _22401_/D vssd1 vssd1 vccd1 vccd1 _22401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_338_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23381_ _23573_/CLK _23381_/D vssd1 vssd1 vccd1 vccd1 _23381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20593_ _20628_/A vssd1 vssd1 vccd1 vccd1 _20593_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22332_ _23564_/CLK _22332_/D vssd1 vssd1 vccd1 vccd1 _22332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_353_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_337_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_353_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22263_ _23555_/CLK _22263_/D vssd1 vssd1 vccd1 vccd1 _22263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21214_ _13440_/B _15035_/X _21214_/S vssd1 vssd1 vccd1 vccd1 _21215_/B sky130_fd_sc_hd__mux2_8
XFILLER_2_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22194_ _22167_/A _22170_/B _22166_/Y vssd1 vssd1 vccd1 vccd1 _22195_/C sky130_fd_sc_hd__o21ai_1
XFILLER_117_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21145_ _20680_/A _21140_/X _21142_/X _20525_/C _21135_/X vssd1 vssd1 vccd1 vccd1
+ _21145_/X sky130_fd_sc_hd__a221o_1
XFILLER_105_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_330_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21076_ _21076_/A _21550_/A vssd1 vssd1 vccd1 vccd1 _21078_/C sky130_fd_sc_hd__nand2_1
XFILLER_101_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_293_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20027_ _20027_/A _20042_/C vssd1 vssd1 vccd1 vccd1 _20027_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _11800_/A vssd1 vssd1 vccd1 vccd1 _11800_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _12780_/A vssd1 vssd1 vccd1 vccd1 _12906_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21978_ _21978_/A _21978_/B vssd1 vssd1 vccd1 vccd1 _21978_/X sky130_fd_sc_hd__xor2_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23717_ _23851_/CLK _23717_/D vssd1 vssd1 vccd1 vccd1 _23717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _12216_/A vssd1 vssd1 vccd1 vccd1 _12269_/A sky130_fd_sc_hd__buf_2
XFILLER_70_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20929_ _15329_/A _20922_/X _20645_/B _20926_/X vssd1 vssd1 vccd1 vccd1 _20929_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_242_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14450_ _14450_/A vssd1 vssd1 vccd1 vccd1 _14450_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_329_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23648_ _23649_/CLK _23648_/D vssd1 vssd1 vccd1 vccd1 _23648_/Q sky130_fd_sc_hd__dfxtp_1
X_11662_ _12144_/A vssd1 vssd1 vccd1 vccd1 _12141_/A sky130_fd_sc_hd__buf_2
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_329_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_329_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13401_ _13399_/A _13239_/C _13244_/X vssd1 vssd1 vccd1 vccd1 _13402_/B sky130_fd_sc_hd__a21o_1
X_11593_ _22310_/Q _23446_/Q _12042_/S vssd1 vssd1 vccd1 vccd1 _11594_/B sky130_fd_sc_hd__mux2_1
X_14381_ _14848_/A _14381_/B vssd1 vssd1 vccd1 vccd1 _15253_/A sky130_fd_sc_hd__nor2_1
X_23579_ _23581_/CLK _23579_/D vssd1 vssd1 vccd1 vccd1 _23579_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_317_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16120_ _23007_/Q _16944_/A _16085_/X input236/X vssd1 vssd1 vccd1 vccd1 _22219_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_10_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13332_ _13510_/B _12603_/X _13353_/B vssd1 vssd1 vccd1 vccd1 _13333_/B sky130_fd_sc_hd__o21a_1
XFILLER_6_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_328_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16051_ _16051_/A vssd1 vssd1 vccd1 vccd1 _22288_/D sky130_fd_sc_hd__clkbuf_1
X_13263_ _23329_/Q _23297_/Q _23265_/Q _23553_/Q _11206_/X _11208_/X vssd1 vssd1 vccd1
+ vccd1 _13264_/B sky130_fd_sc_hd__mux4_1
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15002_ _22919_/Q _15000_/X _15001_/X _14989_/X vssd1 vssd1 vccd1 vccd1 _15002_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_157_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12214_ _12383_/A _12214_/B vssd1 vssd1 vccd1 vccd1 _12214_/X sky130_fd_sc_hd__or2_1
XFILLER_312_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13194_ _13095_/A _13189_/X _13193_/X _11134_/A vssd1 vssd1 vccd1 vccd1 _13194_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_307_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19810_ _19810_/A vssd1 vssd1 vccd1 vccd1 _23541_/D sky130_fd_sc_hd__clkbuf_1
X_12145_ _12007_/A _12142_/X _12144_/X _12797_/A vssd1 vssd1 vccd1 vccd1 _12145_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_7_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23561_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_269_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19741_ _19223_/X _23511_/Q _19743_/S vssd1 vssd1 vccd1 vccd1 _19742_/A sky130_fd_sc_hd__mux2_1
X_16953_ _16962_/A _16953_/B vssd1 vssd1 vccd1 vccd1 _17145_/B sky130_fd_sc_hd__nor2_1
X_12076_ _11774_/A _12071_/Y _12073_/Y _12075_/Y vssd1 vssd1 vccd1 vccd1 _12076_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_278_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15904_ _23613_/Q _14450_/A _14455_/A _23645_/Q vssd1 vssd1 vccd1 vccd1 _15904_/X
+ sky130_fd_sc_hd__o22a_2
X_19672_ _19672_/A vssd1 vssd1 vccd1 vccd1 _23480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16884_ _16883_/X _22542_/Q _16893_/S vssd1 vssd1 vccd1 vccd1 _16885_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_202_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23144_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18623_ _16914_/X _23044_/Q _18623_/S vssd1 vssd1 vccd1 vccd1 _18624_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15835_ _22968_/Q _15835_/B vssd1 vssd1 vccd1 vccd1 _15835_/X sky130_fd_sc_hd__or2_1
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18554_ _18610_/A vssd1 vssd1 vccd1 vccd1 _18623_/S sky130_fd_sc_hd__buf_6
X_15766_ _22934_/Q _14752_/A _14753_/A _18418_/A vssd1 vssd1 vccd1 vccd1 _15766_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_307_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12978_ _22476_/Q _22636_/Q _12978_/S vssd1 vssd1 vccd1 vccd1 _12978_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _22660_/Q _16252_/X _17505_/S vssd1 vssd1 vccd1 vccd1 _17506_/A sky130_fd_sc_hd__mux2_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14717_ input152/X _13651_/B _14719_/S input116/X _14235_/X vssd1 vssd1 vccd1 vccd1
+ _14717_/X sky130_fd_sc_hd__a221o_4
XFILLER_233_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18485_ _18480_/X _18484_/Y _18476_/X vssd1 vssd1 vccd1 vccd1 _22989_/D sky130_fd_sc_hd__a21oi_1
XFILLER_261_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11929_ _23309_/Q _23277_/Q _23245_/Q _23533_/Q _11799_/X _11800_/X vssd1 vssd1 vccd1
+ vccd1 _11929_/X sky130_fd_sc_hd__mux4_1
XFILLER_307_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15697_ _15697_/A _17182_/A vssd1 vssd1 vccd1 vccd1 _15697_/Y sky130_fd_sc_hd__nor2_1
XFILLER_220_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17436_ _17436_/A vssd1 vssd1 vccd1 vccd1 _22629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14648_ _14646_/X _14647_/X _14665_/S vssd1 vssd1 vccd1 vccd1 _14648_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17367_ _22604_/Q input198/X _17369_/S vssd1 vssd1 vccd1 vccd1 _17368_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14579_ input142/X input170/X _14719_/S vssd1 vssd1 vccd1 vccd1 _14579_/X sky130_fd_sc_hd__mux2_8
XFILLER_146_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19106_ _19106_/A vssd1 vssd1 vccd1 vccd1 _23242_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16318_ _14811_/X _22327_/Q _16322_/S vssd1 vssd1 vccd1 vccd1 _16319_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_348_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_308_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17298_ _17298_/A vssd1 vssd1 vccd1 vccd1 _17298_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_307_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19037_ _19037_/A vssd1 vssd1 vccd1 vccd1 _23212_/D sky130_fd_sc_hd__clkbuf_1
X_16249_ _18814_/A vssd1 vssd1 vccd1 vccd1 _16249_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_322_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_350_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_303_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_288_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19939_ _13640_/A _19969_/B _19968_/A _19969_/D vssd1 vssd1 vccd1 vccd1 _19978_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_275_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22950_ _23602_/CLK _22950_/D vssd1 vssd1 vccd1 vccd1 _22950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21901_ _13432_/A _13432_/B _22045_/A _15716_/X vssd1 vssd1 vccd1 vccd1 _21901_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_228_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22881_ _23327_/CLK _22881_/D vssd1 vssd1 vccd1 vccd1 _22881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21832_ _17163_/A _21479_/X _21815_/Y _21831_/X _21681_/X vssd1 vssd1 vccd1 vccd1
+ _23927_/D sky130_fd_sc_hd__o221a_1
XFILLER_24_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21763_ _21763_/A _21763_/B vssd1 vssd1 vccd1 vccd1 _21765_/A sky130_fd_sc_hd__nand2_1
XPHY_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23502_ _23502_/CLK _23502_/D vssd1 vssd1 vccd1 vccd1 _23502_/Q sky130_fd_sc_hd__dfxtp_1
X_20714_ _21077_/B _20692_/X _20702_/X vssd1 vssd1 vccd1 vccd1 _20714_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_178_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_77_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23070_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_211_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21694_ _21694_/A _21694_/B vssd1 vssd1 vccd1 vccd1 _21694_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_357_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23433_ _23558_/CLK _23433_/D vssd1 vssd1 vccd1 vccd1 _23433_/Q sky130_fd_sc_hd__dfxtp_1
X_20645_ _20665_/A _20645_/B _20645_/C vssd1 vssd1 vccd1 vccd1 _20645_/X sky130_fd_sc_hd__or3_1
XFILLER_338_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_326_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23364_ _23578_/CLK _23364_/D vssd1 vssd1 vccd1 vccd1 _23364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20576_ _21351_/A _20572_/X _20575_/Y vssd1 vssd1 vccd1 vccd1 _20577_/C sky130_fd_sc_hd__a21oi_2
XFILLER_258_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_326_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22315_ _22801_/CLK _22315_/D vssd1 vssd1 vccd1 vccd1 _22315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23295_ _23423_/CLK _23295_/D vssd1 vssd1 vccd1 vccd1 _23295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_353_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22246_ _22246_/A vssd1 vssd1 vccd1 vccd1 _22246_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_344_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_322_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22177_ _22177_/A _22177_/B vssd1 vssd1 vccd1 vccd1 _22183_/A sky130_fd_sc_hd__nand2_2
XFILLER_106_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21128_ _21134_/A _21128_/B vssd1 vssd1 vccd1 vccd1 _23858_/D sky130_fd_sc_hd__nor2_1
XFILLER_321_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_289_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13950_ _21636_/A vssd1 vssd1 vccd1 vccd1 _13951_/B sky130_fd_sc_hd__buf_8
XFILLER_47_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21059_ _20731_/A _21047_/X _21058_/X _21049_/X vssd1 vssd1 vccd1 vccd1 _23838_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_275_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12901_ _12897_/A _12898_/X _12900_/X _12797_/X vssd1 vssd1 vccd1 vccd1 _12901_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13881_ _14250_/A _13603_/X _14216_/B _13879_/A vssd1 vssd1 vccd1 vccd1 _15112_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_47_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15620_ _15620_/A vssd1 vssd1 vccd1 vccd1 _15780_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _12818_/A _12831_/X _11132_/A vssd1 vssd1 vccd1 vccd1 _12832_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _23732_/Q _23862_/Q _15806_/S vssd1 vssd1 vccd1 vccd1 _15551_/X sky130_fd_sc_hd__mux2_1
X_12763_ _12700_/X _12748_/Y _12753_/Y _12758_/Y _12762_/Y vssd1 vssd1 vccd1 vccd1
+ _12763_/X sky130_fd_sc_hd__o32a_2
XFILLER_261_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _15735_/A vssd1 vssd1 vccd1 vccd1 _15501_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_159_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _18275_/A _18275_/C _18175_/X vssd1 vssd1 vccd1 vccd1 _18270_/Y sky130_fd_sc_hd__a21oi_1
X_11714_ _11698_/A _11712_/X _11713_/X vssd1 vssd1 vccd1 vccd1 _11714_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_349_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15482_ _21762_/A _15529_/C vssd1 vssd1 vccd1 vccd1 _15482_/Y sky130_fd_sc_hd__xnor2_4
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12818_/A _12693_/X _11132_/A vssd1 vssd1 vccd1 vccd1 _12694_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_348_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17221_ _14167_/X _15846_/Y _17222_/B _17220_/Y vssd1 vssd1 vccd1 vccd1 _17221_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_203_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _16016_/A _14550_/C _14433_/S vssd1 vssd1 vccd1 vccd1 _14465_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11645_ _11919_/A vssd1 vssd1 vccd1 vccd1 _11646_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_329_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17152_ _17073_/X _17150_/Y _17151_/Y _17024_/X vssd1 vssd1 vccd1 vccd1 _17152_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_168_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14364_ _12344_/X _12368_/X _12370_/Y _12371_/X _15565_/A vssd1 vssd1 vccd1 vccd1
+ _15385_/S sky130_fd_sc_hd__o311a_4
Xinput15 core_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_2
XFILLER_345_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11576_ _22374_/Q _22406_/Q _22695_/Q _23062_/Q _12978_/S _12685_/A vssd1 vssd1 vccd1
+ vccd1 _11576_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput26 core_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput37 core_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_1
X_16103_ _23746_/Q _23876_/Q _16103_/S vssd1 vssd1 vccd1 vccd1 _16103_/X sky130_fd_sc_hd__mux2_1
Xinput48 dout0[14] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__buf_2
X_13315_ _13554_/A _11489_/Y _13309_/X _13427_/B vssd1 vssd1 vccd1 vccd1 _13410_/A
+ sky130_fd_sc_hd__a31oi_4
Xinput59 dout0[24] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_2
XFILLER_345_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17083_ _17324_/A vssd1 vssd1 vccd1 vccd1 _17083_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_318_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14295_ _14952_/S vssd1 vssd1 vccd1 vccd1 _15129_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_109_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16034_ _16034_/A _16034_/B vssd1 vssd1 vccd1 vccd1 _16034_/X sky130_fd_sc_hd__or2_1
X_13246_ _13246_/A _14274_/B vssd1 vssd1 vccd1 vccd1 _13246_/Y sky130_fd_sc_hd__nor2_1
XFILLER_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_313_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13177_ _22382_/Q _22414_/Q _22703_/Q _23070_/Q _11543_/A _13127_/X vssd1 vssd1 vccd1
+ vccd1 _13177_/X sky130_fd_sc_hd__mux4_2
XFILLER_272_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_297_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12128_ _12117_/A _12127_/X _11131_/A vssd1 vssd1 vccd1 vccd1 _12128_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_229_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17985_ _22838_/Q _17981_/X _17984_/X _17979_/X vssd1 vssd1 vccd1 vccd1 _22838_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12059_ _12052_/Y _12054_/Y _12056_/Y _12058_/Y _11559_/A vssd1 vssd1 vccd1 vccd1
+ _12059_/X sky130_fd_sc_hd__o221a_1
X_16936_ _22249_/D _16936_/B _16936_/C vssd1 vssd1 vccd1 vccd1 _16942_/C sky130_fd_sc_hd__or3_1
X_19724_ _19197_/X _23503_/Q _19732_/S vssd1 vssd1 vccd1 vccd1 _19725_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16867_ _19217_/A vssd1 vssd1 vccd1 vccd1 _16867_/X sky130_fd_sc_hd__clkbuf_2
X_19655_ _19655_/A vssd1 vssd1 vccd1 vccd1 _23472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18606_ _16889_/X _23036_/Q _18608_/S vssd1 vssd1 vccd1 vccd1 _18607_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15818_ _15818_/A _15818_/B _15818_/C vssd1 vssd1 vccd1 vccd1 _15818_/X sky130_fd_sc_hd__and3_1
XFILLER_280_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19586_ _23442_/Q _19207_/A _19588_/S vssd1 vssd1 vccd1 vccd1 _19587_/A sky130_fd_sc_hd__mux2_1
X_16798_ _16804_/A _16798_/B vssd1 vssd1 vccd1 vccd1 _16799_/A sky130_fd_sc_hd__or2_1
XFILLER_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18537_ _18549_/B _18537_/B vssd1 vssd1 vccd1 vccd1 _18537_/Y sky130_fd_sc_hd__nor2_1
X_15749_ _19226_/A vssd1 vssd1 vccd1 vccd1 _15749_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18468_ _18534_/B vssd1 vssd1 vccd1 vccd1 _18478_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_339_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17419_ _22622_/Q _16233_/X _17421_/S vssd1 vssd1 vccd1 vccd1 _17420_/A sky130_fd_sc_hd__mux2_1
X_18399_ _15501_/A _18400_/C _22961_/Q vssd1 vssd1 vccd1 vccd1 _18401_/B sky130_fd_sc_hd__a21oi_1
XFILLER_193_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_308_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20430_ _20604_/A _20428_/X _20429_/X _20420_/X vssd1 vssd1 vccd1 vccd1 _23691_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_348_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_295_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_335_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20361_ _20333_/X _20723_/A _20357_/X _20360_/X vssd1 vssd1 vccd1 vccd1 _23677_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22100_ _22100_/A _22100_/B vssd1 vssd1 vccd1 vccd1 _22101_/B sky130_fd_sc_hd__nor2_1
X_23080_ _23528_/CLK _23080_/D vssd1 vssd1 vccd1 vccd1 _23080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20292_ _20323_/A _21033_/A vssd1 vssd1 vccd1 vccd1 _20292_/Y sky130_fd_sc_hd__nand2_1
XFILLER_316_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_350_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_195_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23558_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22031_ _22031_/A _22031_/B vssd1 vssd1 vccd1 vccd1 _22031_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_322_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_124_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23652_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_303_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_291_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22933_ _23602_/CLK _22933_/D vssd1 vssd1 vccd1 vccd1 _22933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22864_ _23599_/CLK _22864_/D vssd1 vssd1 vccd1 vccd1 _22864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_272_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21815_ _21813_/X _21814_/Y _22234_/A vssd1 vssd1 vccd1 vccd1 _21815_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22795_ _23575_/CLK _22795_/D vssd1 vssd1 vccd1 vccd1 _22795_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_349_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21746_ _22130_/B vssd1 vssd1 vccd1 vccd1 _21746_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21677_ _21677_/A vssd1 vssd1 vccd1 vccd1 _21677_/X sky130_fd_sc_hd__buf_2
XFILLER_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11430_ _13089_/A vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__buf_4
X_23416_ _23546_/CLK _23416_/D vssd1 vssd1 vccd1 vccd1 _23416_/Q sky130_fd_sc_hd__dfxtp_1
X_20628_ _20628_/A vssd1 vssd1 vccd1 vccd1 _20628_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_326_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_295_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11361_ _12156_/A vssd1 vssd1 vccd1 vccd1 _12864_/A sky130_fd_sc_hd__buf_4
XFILLER_138_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23347_ _23507_/CLK _23347_/D vssd1 vssd1 vccd1 vccd1 _23347_/Q sky130_fd_sc_hd__dfxtp_1
X_20559_ _20602_/A vssd1 vssd1 vccd1 vccd1 _20559_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_295_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_342_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13100_ _23327_/Q _23295_/Q _23263_/Q _23551_/Q _13034_/S _13096_/X vssd1 vssd1 vccd1
+ vccd1 _13101_/B sky130_fd_sc_hd__mux4_1
XFILLER_153_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_298_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14080_ _14080_/A vssd1 vssd1 vccd1 vccd1 _14081_/A sky130_fd_sc_hd__clkbuf_2
X_11292_ _12321_/A vssd1 vssd1 vccd1 vccd1 _12316_/A sky130_fd_sc_hd__buf_4
XFILLER_152_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23278_ _23534_/CLK _23278_/D vssd1 vssd1 vccd1 vccd1 _23278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_341_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_298_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13031_ _13329_/A _13018_/X _13030_/Y vssd1 vssd1 vccd1 vccd1 _13399_/A sky130_fd_sc_hd__a21o_4
X_22229_ _20400_/A _21900_/B _16165_/Y _21842_/X vssd1 vssd1 vccd1 vccd1 _22229_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_6810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17770_ _22761_/Q _17598_/X _17776_/S vssd1 vssd1 vccd1 vccd1 _17771_/A sky130_fd_sc_hd__mux2_1
XTAP_6898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_304_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14982_ _12596_/Y _14530_/X _14979_/X _21437_/A _14703_/X vssd1 vssd1 vccd1 vccd1
+ _18785_/A sky130_fd_sc_hd__a32o_4
XFILLER_219_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16721_ _16721_/A vssd1 vssd1 vccd1 vccd1 _22494_/D sky130_fd_sc_hd__clkbuf_1
X_13933_ _13933_/A _14093_/A vssd1 vssd1 vccd1 vccd1 _13933_/Y sky130_fd_sc_hd__nor2_2
XFILLER_247_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19440_ _23377_/Q _18811_/X _19444_/S vssd1 vssd1 vccd1 vccd1 _19441_/A sky130_fd_sc_hd__mux2_1
X_16652_ _16652_/A vssd1 vssd1 vccd1 vccd1 _22473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13864_ _13864_/A _13864_/B vssd1 vssd1 vccd1 vccd1 _13864_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_505 _15377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15603_ _14730_/X _15591_/X _15602_/X _14748_/X vssd1 vssd1 vccd1 vccd1 _15603_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_222_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_516 _22488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19371_ _19371_/A vssd1 vssd1 vccd1 vccd1 _23346_/D sky130_fd_sc_hd__clkbuf_1
X_12815_ _13608_/A _13350_/A _12806_/Y _12814_/X vssd1 vssd1 vccd1 vccd1 _13329_/A
+ sky130_fd_sc_hd__a31o_2
XINSDIODE2_527 _14018_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16583_ _16583_/A vssd1 vssd1 vccd1 vccd1 _22442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_538 _23912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13795_ _13807_/A _14043_/C vssd1 vssd1 vccd1 vccd1 _13795_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_549 _13615_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18322_ _15724_/X _18323_/C _22934_/Q vssd1 vssd1 vccd1 vccd1 _18324_/B sky130_fd_sc_hd__a21oi_1
XFILLER_215_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15534_ _13738_/A _15865_/B _15533_/Y _13834_/A vssd1 vssd1 vccd1 vccd1 _15534_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _12746_/A vssd1 vssd1 vccd1 vccd1 _12746_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_349_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _22913_/Q _18253_/B vssd1 vssd1 vccd1 vccd1 _18253_/X sky130_fd_sc_hd__or2_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15465_ _15676_/A _21238_/A _15464_/X _15775_/A vssd1 vssd1 vccd1 vccd1 _15465_/X
+ sky130_fd_sc_hd__o22a_1
X_12677_ _11195_/A _12676_/X _12683_/A vssd1 vssd1 vccd1 vccd1 _12677_/X sky130_fd_sc_hd__a21o_1
XFILLER_176_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17204_ _13454_/A _17009_/S _17203_/X vssd1 vssd1 vccd1 vccd1 _17204_/X sky130_fd_sc_hd__o21a_1
XFILLER_31_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14416_ _14416_/A _14416_/B _14458_/B _14458_/A vssd1 vssd1 vccd1 vccd1 _14447_/A
+ sky130_fd_sc_hd__or4bb_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18184_ _18118_/X _18162_/A _18135_/X _18183_/X vssd1 vssd1 vccd1 vccd1 _22891_/D
+ sky130_fd_sc_hd__o211a_1
X_11628_ _13225_/A _12801_/A _11401_/A _11627_/Y vssd1 vssd1 vccd1 vccd1 _13536_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15396_ _23601_/Q vssd1 vssd1 vccd1 vccd1 _19975_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17135_ _23475_/Q _17113_/X _17114_/X _17094_/X _17134_/Y vssd1 vssd1 vccd1 vccd1
+ _17135_/X sky130_fd_sc_hd__a32o_1
X_14347_ _14341_/X _14345_/X _14841_/S vssd1 vssd1 vccd1 vccd1 _14347_/X sky130_fd_sc_hd__mux2_1
X_11559_ _11559_/A vssd1 vssd1 vccd1 vccd1 _11559_/X sky130_fd_sc_hd__buf_2
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17066_ _16951_/X _17065_/X _17078_/A _16968_/X vssd1 vssd1 vccd1 vccd1 _17066_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14278_ _14275_/X _14277_/Y _14310_/S vssd1 vssd1 vccd1 vccd1 _14278_/X sky130_fd_sc_hd__mux2_1
X_16017_ _15865_/A _15332_/Y _15942_/X vssd1 vssd1 vccd1 vccd1 _21274_/A sky130_fd_sc_hd__a21oi_4
X_13229_ _13229_/A _13229_/B vssd1 vssd1 vccd1 vccd1 _13229_/X sky130_fd_sc_hd__or2_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17968_ _22833_/Q _17965_/X _17967_/X _17963_/X vssd1 vssd1 vccd1 vccd1 _22833_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19707_ _19707_/A vssd1 vssd1 vccd1 vccd1 _23495_/D sky130_fd_sc_hd__clkbuf_1
X_16919_ _14001_/A _13671_/Y _16918_/X vssd1 vssd1 vccd1 vccd1 _16927_/B sky130_fd_sc_hd__a21o_4
XFILLER_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17899_ _17933_/A vssd1 vssd1 vccd1 vccd1 _17899_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19638_ _19178_/X _23465_/Q _19638_/S vssd1 vssd1 vccd1 vccd1 _19639_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19569_ _23434_/Q _19181_/A _19577_/S vssd1 vssd1 vccd1 vccd1 _19570_/A sky130_fd_sc_hd__mux2_1
XFILLER_209_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21600_ _21600_/A vssd1 vssd1 vccd1 vccd1 _21845_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22580_ _23643_/CLK _22580_/D vssd1 vssd1 vccd1 vccd1 _22580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21531_ _23820_/Q _23754_/Q vssd1 vssd1 vccd1 vccd1 _21533_/A sky130_fd_sc_hd__or2_1
XFILLER_355_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21462_ _21462_/A _21462_/B vssd1 vssd1 vccd1 vccd1 _21463_/B sky130_fd_sc_hd__xnor2_1
XFILLER_119_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23201_ _23451_/CLK _23201_/D vssd1 vssd1 vccd1 vccd1 _23201_/Q sky130_fd_sc_hd__dfxtp_1
X_20413_ _20482_/B vssd1 vssd1 vccd1 vccd1 _20413_/X sky130_fd_sc_hd__buf_2
XFILLER_309_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21393_ _21393_/A _21393_/B vssd1 vssd1 vccd1 vccd1 _21393_/X sky130_fd_sc_hd__xor2_2
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_324_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23132_ _23420_/CLK _23132_/D vssd1 vssd1 vccd1 vccd1 _23132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20344_ _20344_/A vssd1 vssd1 vccd1 vccd1 _20391_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_350_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23063_ _23446_/CLK _23063_/D vssd1 vssd1 vccd1 vccd1 _23063_/Q sky130_fd_sc_hd__dfxtp_1
X_20275_ _20275_/A _20275_/B vssd1 vssd1 vccd1 vccd1 _20275_/X sky130_fd_sc_hd__or2_1
XTAP_6106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_289_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22014_ _20347_/A _22045_/A _15891_/B _22046_/A vssd1 vssd1 vccd1 vccd1 _22014_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_350_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_304_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_303_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput205 localMemory_wb_adr_i[23] vssd1 vssd1 vccd1 vccd1 _13662_/B sky130_fd_sc_hd__buf_6
XTAP_5416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput216 localMemory_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input216/X sky130_fd_sc_hd__buf_6
XTAP_5427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput227 localMemory_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 input227/X sky130_fd_sc_hd__buf_8
XTAP_5438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput238 localMemory_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 input238/X sky130_fd_sc_hd__buf_8
XTAP_5449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput249 localMemory_wb_sel_i[2] vssd1 vssd1 vccd1 vccd1 input249/X sky130_fd_sc_hd__clkbuf_1
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22916_ _23599_/CLK _22916_/D vssd1 vssd1 vccd1 vccd1 _22916_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_245_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_92_wb_clk_i clkbuf_opt_4_1_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23888_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23896_ _23896_/CLK _23896_/D vssd1 vssd1 vccd1 vccd1 _23896_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_244_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22847_ _23426_/CLK _22847_/D vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dfxtp_1
XFILLER_232_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_21_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23527_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_232_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12600_ _12600_/A _12600_/B vssd1 vssd1 vccd1 vccd1 _13334_/D sky130_fd_sc_hd__nor2_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13580_/A _13580_/B vssd1 vssd1 vccd1 vccd1 _13581_/B sky130_fd_sc_hd__nand2_4
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22778_ _23496_/CLK _22778_/D vssd1 vssd1 vccd1 vccd1 _22778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _22357_/Q _22389_/Q _22678_/Q _23045_/Q _12535_/S _11609_/A vssd1 vssd1 vccd1
+ vccd1 _12532_/B sky130_fd_sc_hd__mux4_2
XFILLER_197_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21729_ _21942_/A _21729_/B vssd1 vssd1 vccd1 vccd1 _21729_/Y sky130_fd_sc_hd__nor2_1
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_303_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _15250_/A vssd1 vssd1 vccd1 vccd1 _15250_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12462_ _22358_/Q _22390_/Q _22679_/Q _23046_/Q _11411_/A _12449_/X vssd1 vssd1 vccd1
+ vccd1 _12463_/B sky130_fd_sc_hd__mux4_2
XFILLER_32_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14201_ _20530_/B _14200_/Y _22711_/Q vssd1 vssd1 vccd1 vccd1 _21289_/B sky130_fd_sc_hd__a21oi_2
X_11413_ _11413_/A vssd1 vssd1 vccd1 vccd1 _11414_/A sky130_fd_sc_hd__buf_4
XFILLER_126_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15181_ _15181_/A vssd1 vssd1 vccd1 vccd1 _15181_/X sky130_fd_sc_hd__clkbuf_2
X_12393_ _13901_/A _12596_/B vssd1 vssd1 vccd1 vccd1 _12393_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_326_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14132_ _14132_/A _14172_/B _14172_/C _14132_/D vssd1 vssd1 vccd1 vccd1 _20532_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_341_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11344_ _23897_/Q vssd1 vssd1 vccd1 vccd1 _11678_/A sky130_fd_sc_hd__buf_2
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_330_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_314_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18940_ _23170_/Q _18865_/X _18940_/S vssd1 vssd1 vccd1 vccd1 _18941_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14063_ _14049_/X _13855_/B _14009_/X input234/X vssd1 vssd1 vccd1 vccd1 _14063_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_7330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11275_ _11275_/A vssd1 vssd1 vccd1 vccd1 _11276_/A sky130_fd_sc_hd__buf_6
XFILLER_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13014_ _13026_/A _14307_/B vssd1 vssd1 vccd1 vccd1 _13015_/B sky130_fd_sc_hd__nor2_1
XFILLER_295_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_315_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18871_ _18871_/A vssd1 vssd1 vccd1 vccd1 _18871_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_7385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17822_ _22784_/Q _17569_/X _17826_/S vssd1 vssd1 vccd1 vccd1 _17823_/A sky130_fd_sc_hd__mux2_1
XTAP_6684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_310_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_310_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14965_ input154/X _13650_/A _15057_/S input119/X _14235_/A vssd1 vssd1 vccd1 vccd1
+ _14965_/X sky130_fd_sc_hd__a221o_4
XFILLER_248_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17753_ _17753_/A vssd1 vssd1 vccd1 vccd1 _22753_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16704_ _16704_/A _16704_/B vssd1 vssd1 vccd1 vccd1 _16705_/A sky130_fd_sc_hd__or2_1
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13916_ _13967_/B _13991_/B vssd1 vssd1 vccd1 vccd1 _13917_/A sky130_fd_sc_hd__and2_2
X_17684_ _17730_/S vssd1 vssd1 vccd1 vccd1 _17693_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_208_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14896_ _14896_/A vssd1 vssd1 vccd1 vccd1 _15097_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_251_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_302 _15990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_331_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16635_ _16635_/A vssd1 vssd1 vccd1 vccd1 _22465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19423_ _19423_/A vssd1 vssd1 vccd1 vccd1 _23369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13847_ _13847_/A _13864_/B vssd1 vssd1 vccd1 vccd1 _13847_/Y sky130_fd_sc_hd__nor2_1
XINSDIODE2_313 _22139_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_324 _16107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_335 _17071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_346 _17207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_357 _17264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16566_ _15474_/X _22435_/Q _16568_/S vssd1 vssd1 vccd1 vccd1 _16567_/A sky130_fd_sc_hd__mux2_1
X_19354_ _19354_/A vssd1 vssd1 vccd1 vccd1 _23338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_349_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_368 _23476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13778_ _13778_/A _13875_/B vssd1 vssd1 vccd1 vccd1 _13835_/A sky130_fd_sc_hd__and2_1
XINSDIODE2_379 _22498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18305_ _18305_/A _22928_/Q _18305_/C vssd1 vssd1 vccd1 vccd1 _18306_/C sky130_fd_sc_hd__and3_1
X_15517_ _15482_/Y _15516_/X _16079_/A vssd1 vssd1 vccd1 vccd1 _15517_/X sky130_fd_sc_hd__mux2_1
X_12729_ _22376_/Q _22408_/Q _22697_/Q _23064_/Q _12727_/X _12728_/X vssd1 vssd1 vccd1
+ vccd1 _12729_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19285_ _19188_/X _23308_/Q _19289_/S vssd1 vssd1 vccd1 vccd1 _19286_/A sky130_fd_sc_hd__mux2_1
XFILLER_337_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16497_ _16497_/A vssd1 vssd1 vccd1 vccd1 _22405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18236_ _22906_/Q _18240_/B vssd1 vssd1 vccd1 vccd1 _18236_/X sky130_fd_sc_hd__or2_1
X_15448_ _23698_/Q _15210_/A _15447_/X vssd1 vssd1 vccd1 vccd1 _15448_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_129_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18167_ _18167_/A vssd1 vssd1 vccd1 vccd1 _18167_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15379_ _15430_/B _15379_/B vssd1 vssd1 vccd1 vccd1 _15379_/Y sky130_fd_sc_hd__nor2_4
XFILLER_306_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17118_ _17073_/A _17117_/X _17107_/X _17078_/X vssd1 vssd1 vccd1 vccd1 _17118_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_144_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_332_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18098_ _18098_/A vssd1 vssd1 vccd1 vccd1 _18098_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_356_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_289_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17049_ _17000_/X _17041_/X _17048_/X _17012_/X vssd1 vssd1 vccd1 vccd1 _17049_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_292_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_289_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20060_ _23629_/Q _20076_/C _20059_/X vssd1 vssd1 vccd1 vccd1 _23629_/D sky130_fd_sc_hd__o21ba_1
XFILLER_225_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_17 _17483_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_28 _17743_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_39 _20101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23750_ _23911_/CLK _23750_/D vssd1 vssd1 vccd1 vccd1 _23750_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20962_ _22029_/A _20950_/X _20721_/B _20954_/X vssd1 vssd1 vccd1 vccd1 _20962_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_66_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22701_ _23068_/CLK _22701_/D vssd1 vssd1 vccd1 vccd1 _22701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23681_ _23714_/CLK _23681_/D vssd1 vssd1 vccd1 vccd1 _23681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20893_ _20925_/A vssd1 vssd1 vccd1 vccd1 _20893_/X sky130_fd_sc_hd__clkbuf_2
X_22632_ _22632_/CLK _22632_/D vssd1 vssd1 vccd1 vccd1 _22632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22563_ _22600_/CLK _22563_/D vssd1 vssd1 vccd1 vccd1 _22563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_356_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_355_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21514_ _21514_/A _21514_/B vssd1 vssd1 vccd1 vccd1 _21514_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_356_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22494_ _23714_/CLK _22494_/D vssd1 vssd1 vccd1 vccd1 _22494_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_182_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21445_ _15037_/A _21619_/B _21442_/Y _20502_/A _21444_/Y vssd1 vssd1 vccd1 vccd1
+ _21485_/A sky130_fd_sc_hd__a221o_1
XFILLER_308_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21376_ _21634_/A vssd1 vssd1 vccd1 vccd1 _21377_/A sky130_fd_sc_hd__buf_2
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_323_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23115_ _23531_/CLK _23115_/D vssd1 vssd1 vccd1 vccd1 _23115_/Q sky130_fd_sc_hd__dfxtp_1
X_20327_ _20327_/A _20400_/B vssd1 vssd1 vccd1 vccd1 _20329_/B sky130_fd_sc_hd__nor2_1
XFILLER_296_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_311_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23046_ _23494_/CLK _23046_/D vssd1 vssd1 vccd1 vccd1 _23046_/Q sky130_fd_sc_hd__dfxtp_1
X_20258_ _20192_/X _21676_/A _20256_/Y _20257_/X vssd1 vssd1 vccd1 vccd1 _20639_/A
+ sky130_fd_sc_hd__a22o_4
XTAP_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20189_ _14879_/X _20169_/A _20190_/B vssd1 vssd1 vccd1 vccd1 _20189_/X sky130_fd_sc_hd__a21o_1
XFILLER_292_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14750_ _15501_/B vssd1 vssd1 vccd1 vccd1 _16109_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11962_ _12119_/S vssd1 vssd1 vccd1 vccd1 _12825_/A sky130_fd_sc_hd__buf_4
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _13701_/A vssd1 vssd1 vccd1 vccd1 _13701_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_233_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14681_ _15090_/A _14671_/X _14677_/X _13505_/X _20138_/B vssd1 vssd1 vccd1 vccd1
+ _14681_/X sky130_fd_sc_hd__a221o_1
XFILLER_205_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23879_ _23910_/CLK _23879_/D vssd1 vssd1 vccd1 vccd1 _23879_/Q sky130_fd_sc_hd__dfxtp_4
X_11893_ _22462_/Q _22622_/Q _11893_/S vssd1 vssd1 vccd1 vccd1 _11893_/X sky130_fd_sc_hd__mux2_1
XFILLER_301_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16420_ _16442_/A vssd1 vssd1 vccd1 vccd1 _16429_/S sky130_fd_sc_hd__buf_6
XFILLER_233_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13632_ _13632_/A _13632_/B _13632_/C vssd1 vssd1 vccd1 vccd1 _13633_/B sky130_fd_sc_hd__nor3_1
XFILLER_60_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_260_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16351_ _15668_/X _22342_/Q _16355_/S vssd1 vssd1 vccd1 vccd1 _16352_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13563_ _13647_/A _23938_/Q _13490_/X _13562_/Y vssd1 vssd1 vccd1 vccd1 _13985_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_358_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15302_ _23663_/Q _16021_/B vssd1 vssd1 vccd1 vccd1 _15302_/X sky130_fd_sc_hd__or2_1
X_19070_ _19070_/A vssd1 vssd1 vccd1 vccd1 _23227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12514_ _22777_/Q _22745_/Q _22646_/Q _22713_/Q _23894_/Q _23895_/Q vssd1 vssd1 vccd1
+ vccd1 _12515_/B sky130_fd_sc_hd__mux4_1
X_16282_ _22316_/Q _16281_/X _16285_/S vssd1 vssd1 vccd1 vccd1 _16283_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_358_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13494_ _12916_/B _12965_/A _13013_/A _13493_/Y vssd1 vssd1 vccd1 vccd1 _13494_/X
+ sky130_fd_sc_hd__o211a_1
X_18021_ _18198_/B _18021_/B vssd1 vssd1 vccd1 vccd1 _18099_/A sky130_fd_sc_hd__or2_2
XFILLER_9_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15233_ _21570_/A _15274_/C vssd1 vssd1 vccd1 vccd1 _15234_/B sky130_fd_sc_hd__xnor2_4
XFILLER_157_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12445_ _22262_/Q _23078_/Q _23494_/Q _22423_/Q _11411_/A _11189_/A vssd1 vssd1 vccd1
+ vccd1 _12446_/B sky130_fd_sc_hd__mux4_2
XFILLER_154_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15164_ _15164_/A vssd1 vssd1 vccd1 vccd1 _15417_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12376_ _11330_/A _12375_/X _11819_/A vssd1 vssd1 vccd1 vccd1 _12376_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14115_ _14119_/A _14119_/B _14119_/C _14119_/D vssd1 vssd1 vccd1 vccd1 _14115_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11327_ _23896_/Q vssd1 vssd1 vccd1 vccd1 _11659_/A sky130_fd_sc_hd__buf_2
XFILLER_326_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19972_ _19981_/A _19980_/C vssd1 vssd1 vccd1 vccd1 _19972_/Y sky130_fd_sc_hd__nor2_1
XFILLER_314_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15095_ _12287_/B _15082_/X _15090_/Y _15094_/X vssd1 vssd1 vccd1 vccd1 _15095_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_330_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18923_ _23162_/Q _18840_/X _18929_/S vssd1 vssd1 vccd1 vccd1 _18924_/A sky130_fd_sc_hd__mux2_1
X_14046_ _14046_/A _14052_/B _14046_/C vssd1 vssd1 vccd1 vccd1 _14046_/X sky130_fd_sc_hd__or3_1
XFILLER_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_326_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11258_ _12544_/B vssd1 vssd1 vccd1 vccd1 _11404_/A sky130_fd_sc_hd__inv_2
XTAP_7171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18854_ _23134_/Q _18852_/X _18866_/S vssd1 vssd1 vccd1 vccd1 _18855_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11189_ _11189_/A vssd1 vssd1 vccd1 vccd1 _12536_/A sky130_fd_sc_hd__clkinv_2
XTAP_6481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_295_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17805_ _17861_/A vssd1 vssd1 vccd1 vccd1 _17874_/S sky130_fd_sc_hd__buf_6
XFILLER_255_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15997_ _13491_/A _15583_/X _14942_/X _13402_/A _15996_/Y vssd1 vssd1 vccd1 vccd1
+ _15997_/X sky130_fd_sc_hd__o221a_1
XFILLER_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18785_ _18785_/A vssd1 vssd1 vccd1 vccd1 _18785_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14948_ _15089_/S _14947_/Y _14860_/X vssd1 vssd1 vccd1 vccd1 _16034_/B sky130_fd_sc_hd__a21o_1
X_17736_ _17736_/A vssd1 vssd1 vccd1 vccd1 _22745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_270_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14879_ _14431_/X _14868_/X _14877_/X _14878_/X _14518_/X vssd1 vssd1 vccd1 vccd1
+ _14879_/X sky130_fd_sc_hd__o32a_4
XINSDIODE2_110 _13875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17667_ _22715_/Q _17553_/X _17671_/S vssd1 vssd1 vccd1 vccd1 _17668_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_121 _13714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19406_ _19406_/A vssd1 vssd1 vccd1 vccd1 _23362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_132 _21900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16618_ _22458_/Q _16220_/X _16618_/S vssd1 vssd1 vccd1 vccd1 _16619_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_143 _20368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17598_ _18824_/A vssd1 vssd1 vccd1 vccd1 _17598_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_250_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_154 _21077_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_165 _13967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_176 _14204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_187 _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19337_ _19264_/X _23332_/Q _19337_/S vssd1 vssd1 vccd1 vccd1 _19338_/A sky130_fd_sc_hd__mux2_1
X_16549_ _15044_/X _22427_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _16550_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_198 _13951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_337_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19268_ _19324_/A vssd1 vssd1 vccd1 vccd1 _19337_/S sky130_fd_sc_hd__buf_8
XFILLER_337_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18219_ _18245_/A vssd1 vssd1 vccd1 vccd1 _18219_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19199_ _19197_/X _23279_/Q _19211_/S vssd1 vssd1 vccd1 vccd1 _19200_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_346_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21230_ _21243_/A vssd1 vssd1 vccd1 vccd1 _21240_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21161_ _21161_/A vssd1 vssd1 vccd1 vccd1 _21161_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_321_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20112_ _23644_/Q _23643_/Q _20112_/C _20112_/D vssd1 vssd1 vccd1 vccd1 _20126_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_259_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21092_ _21122_/A vssd1 vssd1 vccd1 vccd1 _21108_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20043_ _23625_/Q _20051_/A _18268_/A vssd1 vssd1 vccd1 vccd1 _20043_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_259_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23802_ _23942_/CLK _23802_/D vssd1 vssd1 vccd1 vccd1 _23802_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21994_ _21972_/A _21971_/B _21971_/A vssd1 vssd1 vccd1 vccd1 _21995_/B sky130_fd_sc_hd__o21ba_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23733_ _23918_/CLK _23733_/D vssd1 vssd1 vccd1 vccd1 _23733_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20945_ _21856_/A _20936_/X _20683_/B _20940_/X vssd1 vssd1 vccd1 vccd1 _20945_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23664_ _23700_/CLK _23664_/D vssd1 vssd1 vccd1 vccd1 _23664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20876_ _20879_/A _20876_/B vssd1 vssd1 vccd1 vccd1 _20877_/A sky130_fd_sc_hd__and2_1
XFILLER_81_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_329_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22615_ _23558_/CLK _22615_/D vssd1 vssd1 vccd1 vccd1 _22615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23595_ _23637_/CLK _23595_/D vssd1 vssd1 vccd1 vccd1 _23595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22546_ _23582_/CLK _22546_/D vssd1 vssd1 vccd1 vccd1 _22546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_347_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_356_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22477_ _22666_/CLK _22477_/D vssd1 vssd1 vccd1 vccd1 _22477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12230_ _23918_/Q _12283_/B vssd1 vssd1 vccd1 vccd1 _12230_/X sky130_fd_sc_hd__or2_1
XFILLER_107_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21428_ _21543_/B _21428_/B vssd1 vssd1 vccd1 vccd1 _21428_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_170_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12161_ _13615_/A _13351_/A _13623_/A _13342_/A vssd1 vssd1 vccd1 vccd1 _12161_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_136_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21359_ _21456_/A vssd1 vssd1 vccd1 vccd1 _21816_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11112_ _11112_/A vssd1 vssd1 vccd1 vccd1 _11113_/A sky130_fd_sc_hd__buf_6
XFILLER_151_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12092_ _23474_/Q _23570_/Q _22534_/Q _22338_/Q _11637_/A _11755_/A vssd1 vssd1 vccd1
+ vccd1 _12093_/B sky130_fd_sc_hd__mux4_1
XFILLER_268_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23029_ _23349_/CLK _23029_/D vssd1 vssd1 vccd1 vccd1 _23029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_311_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15920_ _15920_/A _15920_/B _15920_/C vssd1 vssd1 vccd1 vccd1 _15920_/X sky130_fd_sc_hd__and3_1
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15851_ _13018_/D _14942_/X _15251_/X _15801_/A _15850_/X vssd1 vssd1 vccd1 vccd1
+ _15851_/X sky130_fd_sc_hd__o221a_1
XFILLER_76_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _15815_/A _14756_/X _14799_/X _15345_/A vssd1 vssd1 vccd1 vccd1 _14802_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15782_ _22998_/Q _15931_/A _15932_/A input227/X vssd1 vssd1 vccd1 vccd1 _21954_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_218_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18570_ _18570_/A vssd1 vssd1 vccd1 vccd1 _23019_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_291_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12994_ _23483_/Q _23579_/Q _22543_/Q _22347_/Q _12727_/X _12728_/X vssd1 vssd1 vccd1
+ vccd1 _12995_/B sky130_fd_sc_hd__mux4_1
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14733_ _14733_/A vssd1 vssd1 vccd1 vccd1 _14902_/A sky130_fd_sc_hd__clkbuf_2
X_17521_ _22667_/Q _16275_/X _17527_/S vssd1 vssd1 vccd1 vccd1 _17522_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11945_ _13521_/A _13521_/B vssd1 vssd1 vccd1 vccd1 _11945_/X sky130_fd_sc_hd__or2b_1
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _22637_/Q _16281_/X _17454_/S vssd1 vssd1 vccd1 vccd1 _17453_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14664_ _14343_/X _14316_/X _14664_/S vssd1 vssd1 vccd1 vccd1 _14664_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11876_ _22786_/Q _22754_/Q _22655_/Q _22722_/Q _12094_/A _11754_/A vssd1 vssd1 vccd1
+ vccd1 _11876_/X sky130_fd_sc_hd__mux4_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16403_ _15168_/X _22364_/Q _16407_/S vssd1 vssd1 vccd1 vccd1 _16404_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13615_ _13615_/A _13615_/B vssd1 vssd1 vccd1 vccd1 _13615_/Y sky130_fd_sc_hd__xnor2_4
X_17383_ _20808_/A vssd1 vssd1 vccd1 vccd1 _20790_/A sky130_fd_sc_hd__buf_8
XFILLER_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14595_ _20161_/A _14595_/B vssd1 vssd1 vccd1 vccd1 _16170_/B sky130_fd_sc_hd__or2_2
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19122_ _23250_/Q _18814_/X _19124_/S vssd1 vssd1 vccd1 vccd1 _19123_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16334_ _16334_/A vssd1 vssd1 vccd1 vccd1 _22334_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_319_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13546_ _13574_/A _13083_/A _13569_/A _13573_/B _13545_/X vssd1 vssd1 vccd1 vccd1
+ _13565_/B sky130_fd_sc_hd__a41o_4
XFILLER_201_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_347_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19053_ _19075_/A vssd1 vssd1 vccd1 vccd1 _19062_/S sky130_fd_sc_hd__buf_4
X_16265_ _18830_/A vssd1 vssd1 vccd1 vccd1 _16265_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_335_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13477_ _16980_/A _13474_/A _13476_/Y _13593_/A vssd1 vssd1 vccd1 vccd1 _13882_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18004_ _22843_/Q _17932_/A _18003_/X _18000_/X vssd1 vssd1 vccd1 vccd1 _22843_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15216_ _15216_/A vssd1 vssd1 vccd1 vccd1 _15216_/X sky130_fd_sc_hd__clkbuf_4
X_23947__506 vssd1 vssd1 vccd1 vccd1 _23947__506/HI core_wb_adr_o[0] sky130_fd_sc_hd__conb_1
X_12428_ _12534_/A _12423_/Y _12425_/Y _12427_/Y vssd1 vssd1 vccd1 vccd1 _12428_/X
+ sky130_fd_sc_hd__a31o_1
X_16196_ _18871_/A vssd1 vssd1 vccd1 vccd1 _19264_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput306 _13955_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[11] sky130_fd_sc_hd__buf_2
XFILLER_299_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput317 _13976_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[22] sky130_fd_sc_hd__buf_2
X_15147_ _23692_/Q _14494_/S _15146_/X vssd1 vssd1 vccd1 vccd1 _15147_/Y sky130_fd_sc_hd__o21ai_4
Xoutput328 _13933_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[7] sky130_fd_sc_hd__buf_2
XFILLER_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_342_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12359_ _12365_/A _12359_/B vssd1 vssd1 vccd1 vccd1 _12359_/Y sky130_fd_sc_hd__nor2_1
XFILLER_330_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_315_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput339 _13787_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[16] sky130_fd_sc_hd__buf_2
XFILLER_236_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_330_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19955_ _23600_/Q _19950_/B _19954_/Y vssd1 vssd1 vccd1 vccd1 _23600_/D sky130_fd_sc_hd__o21a_1
X_15078_ _15078_/A _15256_/B vssd1 vssd1 vccd1 vccd1 _15078_/X sky130_fd_sc_hd__or2_1
XFILLER_303_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18906_ _18906_/A vssd1 vssd1 vccd1 vccd1 _23154_/D sky130_fd_sc_hd__clkbuf_1
X_14029_ input216/X _14027_/X _14028_/X vssd1 vssd1 vccd1 vccd1 _14029_/X sky130_fd_sc_hd__a21o_4
X_19886_ _19886_/A vssd1 vssd1 vccd1 vccd1 _23575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_311_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_353_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_296_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18837_ _18853_/A vssd1 vssd1 vccd1 vccd1 _18850_/S sky130_fd_sc_hd__buf_2
XFILLER_68_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18768_ _18768_/A vssd1 vssd1 vccd1 vccd1 _23108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_270_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17719_ _17719_/A vssd1 vssd1 vccd1 vccd1 _22738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_282_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18699_ _18767_/S vssd1 vssd1 vccd1 vccd1 _18708_/S sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_149_wb_clk_i _23945_/CLK vssd1 vssd1 vccd1 vccd1 _23946_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_212_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20730_ _20730_/A vssd1 vssd1 vccd1 vccd1 _20757_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_169_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_323_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20661_ _20661_/A _20669_/B vssd1 vssd1 vccd1 vccd1 _20665_/B sky130_fd_sc_hd__nor2_8
XFILLER_323_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22400_ _23440_/CLK _22400_/D vssd1 vssd1 vccd1 vccd1 _22400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_337_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23380_ _23414_/CLK _23380_/D vssd1 vssd1 vccd1 vccd1 _23380_/Q sky130_fd_sc_hd__dfxtp_1
X_20592_ _23721_/Q _20542_/X _20591_/X _20559_/X vssd1 vssd1 vccd1 vccd1 _23721_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22331_ _23563_/CLK _22331_/D vssd1 vssd1 vccd1 vccd1 _22331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_353_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22262_ _23494_/CLK _22262_/D vssd1 vssd1 vccd1 vccd1 _22262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_353_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21213_ _21213_/A vssd1 vssd1 vccd1 vccd1 _23883_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_321_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22193_ _22193_/A _22197_/A vssd1 vssd1 vccd1 vccd1 _22195_/B sky130_fd_sc_hd__and2_1
XFILLER_132_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21144_ _23863_/Q _21139_/X _21143_/X _21073_/X vssd1 vssd1 vccd1 vccd1 _23863_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21075_ _23846_/Q vssd1 vssd1 vccd1 vccd1 _21075_/Y sky130_fd_sc_hd__inv_2
XFILLER_247_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20026_ _23620_/Q _20034_/B _20026_/C _20031_/D vssd1 vssd1 vccd1 vccd1 _20042_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_330_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21977_ _21977_/A _21977_/B vssd1 vssd1 vccd1 vccd1 _21978_/B sky130_fd_sc_hd__nand2_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _11914_/A vssd1 vssd1 vccd1 vccd1 _12139_/A sky130_fd_sc_hd__buf_2
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23716_ _23871_/CLK _23716_/D vssd1 vssd1 vccd1 vccd1 _23716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20928_ _23791_/Q _20925_/X _20927_/X _20920_/X vssd1 vssd1 vccd1 vccd1 _23791_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23647_ _23652_/CLK _23647_/D vssd1 vssd1 vccd1 vccd1 _23647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _12406_/A vssd1 vssd1 vccd1 vccd1 _12144_/A sky130_fd_sc_hd__buf_4
XFILLER_202_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20859_ _20859_/A vssd1 vssd1 vccd1 vccd1 _23771_/D sky130_fd_sc_hd__clkbuf_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13400_ _13400_/A _13400_/B _13400_/C _13399_/Y vssd1 vssd1 vccd1 vccd1 _13409_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_186_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_357_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14380_ _14380_/A vssd1 vssd1 vccd1 vccd1 _14380_/Y sky130_fd_sc_hd__inv_2
XFILLER_322_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11592_ _12041_/A vssd1 vssd1 vccd1 vccd1 _11594_/A sky130_fd_sc_hd__buf_4
X_23578_ _23578_/CLK _23578_/D vssd1 vssd1 vccd1 vccd1 _23578_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ _13351_/A vssd1 vssd1 vccd1 vccd1 _13618_/A sky130_fd_sc_hd__inv_2
XFILLER_328_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22529_ _23565_/CLK _22529_/D vssd1 vssd1 vccd1 vccd1 _22529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_317_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16050_ _16049_/X _22288_/Q _16125_/S vssd1 vssd1 vccd1 vccd1 _16051_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13262_ _11236_/X _13253_/Y _13257_/Y _13259_/Y _13261_/Y vssd1 vssd1 vccd1 vccd1
+ _13262_/X sky130_fd_sc_hd__o32a_1
XFILLER_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15001_ _15001_/A vssd1 vssd1 vccd1 vccd1 _15001_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12213_ _23308_/Q _23276_/Q _23244_/Q _23532_/Q _12209_/X _12210_/X vssd1 vssd1 vccd1
+ vccd1 _12214_/B sky130_fd_sc_hd__mux4_2
XFILLER_194_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_324_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13193_ _11435_/A _13190_/X _13192_/X vssd1 vssd1 vccd1 vccd1 _13193_/X sky130_fd_sc_hd__a21o_1
XFILLER_136_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_312_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12144_ _12144_/A _12144_/B vssd1 vssd1 vccd1 vccd1 _12144_/X sky130_fd_sc_hd__or2_1
XFILLER_297_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19740_ _19740_/A vssd1 vssd1 vccd1 vccd1 _23510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16952_ _17145_/A vssd1 vssd1 vccd1 vccd1 _17230_/A sky130_fd_sc_hd__buf_2
X_12075_ _11582_/A _12074_/X _11713_/X vssd1 vssd1 vccd1 vccd1 _12075_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_173_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15903_ _22938_/Q _15903_/B vssd1 vssd1 vccd1 vccd1 _15903_/X sky130_fd_sc_hd__and2_1
XFILLER_38_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_323_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19671_ _19226_/X _23480_/Q _19671_/S vssd1 vssd1 vccd1 vccd1 _19672_/A sky130_fd_sc_hd__mux2_1
X_16883_ _19233_/A vssd1 vssd1 vccd1 vccd1 _16883_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18622_ _18622_/A vssd1 vssd1 vccd1 vccd1 _23043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_265_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15834_ _15833_/X _14752_/X _14753_/X _22968_/Q vssd1 vssd1 vccd1 vccd1 _15834_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18553_ _19164_/A _19483_/B vssd1 vssd1 vccd1 vccd1 _18610_/A sky130_fd_sc_hd__or2_4
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12977_ _22315_/Q _23451_/Q _12977_/S vssd1 vssd1 vccd1 vccd1 _12977_/X sky130_fd_sc_hd__mux2_1
X_15765_ _22966_/Q vssd1 vssd1 vccd1 vccd1 _18418_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _17504_/A vssd1 vssd1 vccd1 vccd1 _22659_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14716_ _22489_/Q _14232_/X _14247_/A _14715_/X _14071_/A vssd1 vssd1 vccd1 vccd1
+ _14716_/X sky130_fd_sc_hd__o221a_1
X_11928_ _12097_/A _11928_/B vssd1 vssd1 vccd1 vccd1 _11928_/X sky130_fd_sc_hd__or2_1
X_18484_ _22989_/Q _18492_/B vssd1 vssd1 vccd1 vccd1 _18484_/Y sky130_fd_sc_hd__nand2_1
X_15696_ _15003_/X _15684_/X _15695_/X vssd1 vssd1 vccd1 vccd1 _17182_/A sky130_fd_sc_hd__o21ai_4
XFILLER_233_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17435_ _22629_/Q _16255_/X _17443_/S vssd1 vssd1 vccd1 vccd1 _17436_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14647_ _14647_/A _14369_/X vssd1 vssd1 vccd1 vccd1 _14647_/X sky130_fd_sc_hd__or2b_1
XFILLER_268_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11859_ _11267_/A _13745_/A _11858_/X _11828_/B vssd1 vssd1 vccd1 vccd1 _13522_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_348_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14578_ _15057_/S vssd1 vssd1 vccd1 vccd1 _14719_/S sky130_fd_sc_hd__clkbuf_4
X_17366_ _17366_/A vssd1 vssd1 vccd1 vccd1 _22603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_347_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19105_ _23242_/Q _18788_/X _19113_/S vssd1 vssd1 vccd1 vccd1 _19106_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16317_ _16317_/A vssd1 vssd1 vccd1 vccd1 _22326_/D sky130_fd_sc_hd__clkbuf_1
X_13529_ _13621_/A _13621_/B _13621_/C _13625_/A _12162_/Y vssd1 vssd1 vccd1 vccd1
+ _13618_/C sky130_fd_sc_hd__a311o_2
XFILLER_158_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17297_ _22219_/A vssd1 vssd1 vccd1 vccd1 _22193_/A sky130_fd_sc_hd__buf_8
XFILLER_335_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16248_ _16248_/A vssd1 vssd1 vccd1 vccd1 _22305_/D sky130_fd_sc_hd__clkbuf_1
X_19036_ _16838_/X _23212_/Q _19040_/S vssd1 vssd1 vccd1 vccd1 _19037_/A sky130_fd_sc_hd__mux2_1
XFILLER_334_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16179_ _15558_/X _16168_/X _16177_/X _16178_/X _14755_/A vssd1 vssd1 vccd1 vccd1
+ _16179_/X sky130_fd_sc_hd__o32a_4
XFILLER_115_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_350_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_303_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_331_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19938_ _23591_/Q _19938_/B _19938_/C vssd1 vssd1 vccd1 vccd1 _19968_/A sky130_fd_sc_hd__and3_1
XFILLER_303_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19869_ _19869_/A vssd1 vssd1 vccd1 vccd1 _23567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21900_ _21900_/A _21900_/B vssd1 vssd1 vccd1 vccd1 _21900_/X sky130_fd_sc_hd__or2_1
X_22880_ _23584_/CLK _22880_/D vssd1 vssd1 vccd1 vccd1 _22880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21831_ _21831_/A _21831_/B _21922_/A vssd1 vssd1 vccd1 vccd1 _21831_/X sky130_fd_sc_hd__or3b_1
XFILLER_71_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21762_ _21762_/A _21766_/A vssd1 vssd1 vccd1 vccd1 _21763_/B sky130_fd_sc_hd__or2_1
XPHY_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23501_ _23565_/CLK _23501_/D vssd1 vssd1 vccd1 vccd1 _23501_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20713_ _20713_/A _20731_/B vssd1 vssd1 vccd1 vccd1 _20716_/B sky130_fd_sc_hd__and2_2
XFILLER_357_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21693_ _21550_/A _21605_/B _21605_/C _21692_/X _21604_/A vssd1 vssd1 vccd1 vccd1
+ _21693_/X sky130_fd_sc_hd__a41o_1
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23432_ _23526_/CLK _23432_/D vssd1 vssd1 vccd1 vccd1 _23432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_339_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20644_ _21652_/A _20572_/X _20643_/Y vssd1 vssd1 vccd1 vccd1 _20645_/C sky130_fd_sc_hd__a21oi_1
XFILLER_338_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_338_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_354_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23363_ _23459_/CLK _23363_/D vssd1 vssd1 vccd1 vccd1 _23363_/Q sky130_fd_sc_hd__dfxtp_1
X_20575_ _14196_/B _20773_/A _20574_/X vssd1 vssd1 vccd1 vccd1 _20575_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_192_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22314_ _23580_/CLK _22314_/D vssd1 vssd1 vccd1 vccd1 _22314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_353_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_326_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23294_ _23456_/CLK _23294_/D vssd1 vssd1 vccd1 vccd1 _23294_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_46_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23951_/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_194_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_353_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22245_ _17315_/X _21714_/A _22234_/Y _22244_/Y _18135_/X vssd1 vssd1 vccd1 vccd1
+ _23942_/D sky130_fd_sc_hd__o221a_1
XFILLER_105_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22176_ _22176_/A _22163_/B vssd1 vssd1 vccd1 vccd1 _22177_/B sky130_fd_sc_hd__or2b_1
XFILLER_87_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21127_ _23858_/Q _21123_/X _21124_/X _20641_/A vssd1 vssd1 vccd1 vccd1 _21128_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_120_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21058_ _23838_/Q _21068_/B vssd1 vssd1 vccd1 vccd1 _21058_/X sky130_fd_sc_hd__or2_1
XFILLER_86_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12900_ _12900_/A _12900_/B vssd1 vssd1 vccd1 vccd1 _12900_/X sky130_fd_sc_hd__or2_1
XFILLER_246_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20009_ _20009_/A _20009_/B _20014_/D vssd1 vssd1 vccd1 vccd1 _20016_/C sky130_fd_sc_hd__and3_1
X_13880_ _13892_/A _14246_/A vssd1 vssd1 vccd1 vccd1 _13880_/Y sky130_fd_sc_hd__nor2_8
XFILLER_101_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12831_ _23420_/Q _23036_/Q _23388_/Q _23356_/Q _12755_/X _12756_/X vssd1 vssd1 vccd1
+ vccd1 _12831_/X sky130_fd_sc_hd__mux4_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _23668_/Q _15905_/B vssd1 vssd1 vccd1 vccd1 _15550_/X sky130_fd_sc_hd__or2_1
X_12762_ _12886_/A _12761_/X _11232_/A vssd1 vssd1 vccd1 vccd1 _12762_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_261_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14501_ _15726_/B vssd1 vssd1 vccd1 vccd1 _15735_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_203_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11713_ _11713_/A vssd1 vssd1 vccd1 vccd1 _11713_/X sky130_fd_sc_hd__buf_2
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15481_ _23925_/Q vssd1 vssd1 vccd1 vccd1 _21762_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _23416_/Q _23032_/Q _23384_/Q _23352_/Q _12692_/X _12041_/X vssd1 vssd1 vccd1
+ vccd1 _12693_/X sky130_fd_sc_hd__mux4_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _23483_/Q _17220_/B vssd1 vssd1 vccd1 vccd1 _17220_/Y sky130_fd_sc_hd__nand2_1
X_14432_ _22903_/Q _14394_/X _14164_/X _22596_/Q vssd1 vssd1 vccd1 vccd1 _14550_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _12475_/A vssd1 vssd1 vccd1 vccd1 _11919_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_345_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17151_ _21790_/A _17174_/B vssd1 vssd1 vccd1 vccd1 _17151_/Y sky130_fd_sc_hd__nand2_1
XFILLER_357_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14363_ _14357_/X _14360_/Y _15085_/S vssd1 vssd1 vccd1 vccd1 _14363_/Y sky130_fd_sc_hd__a21oi_1
X_11575_ _12119_/S vssd1 vssd1 vccd1 vccd1 _12978_/S sky130_fd_sc_hd__buf_4
XFILLER_11_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 core_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput27 core_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_2
X_16102_ _23682_/Q _16102_/B vssd1 vssd1 vccd1 vccd1 _16102_/X sky130_fd_sc_hd__or2_1
XFILLER_156_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput38 core_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
X_13314_ _13314_/A _14388_/C vssd1 vssd1 vccd1 vccd1 _13427_/B sky130_fd_sc_hd__and2_2
XFILLER_337_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17082_ _17082_/A vssd1 vssd1 vccd1 vccd1 _17324_/A sky130_fd_sc_hd__buf_4
XFILLER_183_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput49 dout0[15] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_2
XFILLER_305_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14294_ _14294_/A vssd1 vssd1 vccd1 vccd1 _14952_/S sky130_fd_sc_hd__buf_4
XFILLER_345_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_316_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16033_ _14835_/A _13561_/A _16032_/X vssd1 vssd1 vccd1 vccd1 _16033_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_183_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13245_ _13542_/A vssd1 vssd1 vccd1 vccd1 _13246_/A sky130_fd_sc_hd__inv_2
XFILLER_313_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13176_ _13180_/A _13176_/B vssd1 vssd1 vccd1 vccd1 _13176_/X sky130_fd_sc_hd__or2_1
XFILLER_272_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12127_ _23409_/Q _23025_/Q _23377_/Q _23345_/Q _11151_/A _11953_/A vssd1 vssd1 vccd1
+ vccd1 _12127_/X sky130_fd_sc_hd__mux4_1
XFILLER_112_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17984_ _22837_/Q _17972_/X _17896_/X _17982_/X _17983_/X vssd1 vssd1 vccd1 vccd1
+ _17984_/X sky130_fd_sc_hd__a221o_1
XFILLER_269_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19723_ _19769_/S vssd1 vssd1 vccd1 vccd1 _19732_/S sky130_fd_sc_hd__buf_4
XFILLER_334_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12058_ _12754_/A _12057_/X _12687_/A vssd1 vssd1 vccd1 vccd1 _12058_/Y sky130_fd_sc_hd__o21ai_1
X_16935_ _16942_/A _16935_/B vssd1 vssd1 vccd1 vccd1 _22246_/A sky130_fd_sc_hd__or2_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19654_ _19201_/X _23472_/Q _19660_/S vssd1 vssd1 vccd1 vccd1 _19655_/A sky130_fd_sc_hd__mux2_1
X_16866_ _16866_/A vssd1 vssd1 vccd1 vccd1 _22536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_350_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18605_ _18605_/A vssd1 vssd1 vccd1 vccd1 _23035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15817_ _14822_/A _15794_/X _15816_/Y _14568_/A vssd1 vssd1 vccd1 vccd1 _15818_/C
+ sky130_fd_sc_hd__a211o_1
X_19585_ _19585_/A vssd1 vssd1 vccd1 vccd1 _23441_/D sky130_fd_sc_hd__clkbuf_1
X_16797_ _22516_/Q _16783_/X _16784_/X input31/X vssd1 vssd1 vccd1 vccd1 _16798_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_34_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_350_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18536_ _18536_/A vssd1 vssd1 vccd1 vccd1 _18549_/B sky130_fd_sc_hd__inv_2
XFILLER_240_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15748_ _18833_/A vssd1 vssd1 vccd1 vccd1 _19226_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18467_ _18480_/A vssd1 vssd1 vccd1 vccd1 _18467_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15679_ _12805_/A _15583_/X _15458_/X _15338_/A _15678_/Y vssd1 vssd1 vccd1 vccd1
+ _15679_/X sky130_fd_sc_hd__o221a_1
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_339_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17418_ _17418_/A vssd1 vssd1 vccd1 vccd1 _22621_/D sky130_fd_sc_hd__clkbuf_1
X_18398_ _15501_/A _18400_/C _18397_/Y vssd1 vssd1 vccd1 vccd1 _22960_/D sky130_fd_sc_hd__o21a_1
XFILLER_193_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_320_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17349_ _17371_/A vssd1 vssd1 vccd1 vccd1 _17358_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_20_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_336_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_307_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20360_ _20445_/A vssd1 vssd1 vccd1 vccd1 _20360_/X sky130_fd_sc_hd__buf_2
XFILLER_134_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_350_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19019_ _19075_/A vssd1 vssd1 vccd1 vccd1 _19088_/S sky130_fd_sc_hd__buf_6
XFILLER_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20291_ _20174_/X _20288_/X _20289_/Y _21790_/B _20147_/X vssd1 vssd1 vccd1 vccd1
+ _21033_/A sky130_fd_sc_hd__o32a_4
XFILLER_134_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22030_ _22030_/A _22030_/B vssd1 vssd1 vccd1 vccd1 _22031_/B sky130_fd_sc_hd__nor2_1
XFILLER_115_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_331_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_303_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_330_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_164_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23866_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22932_ _22961_/CLK _22932_/D vssd1 vssd1 vccd1 vccd1 _22932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_290_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22863_ _23008_/CLK _22863_/D vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_228_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_260_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21814_ _23797_/Q _21814_/B vssd1 vssd1 vccd1 vccd1 _21814_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22794_ _23446_/CLK _22794_/D vssd1 vssd1 vccd1 vccd1 _22794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_358_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21745_ _21737_/A _21479_/X _21729_/Y _21744_/X _21681_/X vssd1 vssd1 vccd1 vccd1
+ _23924_/D sky130_fd_sc_hd__o221a_2
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21676_ _21676_/A _21676_/B vssd1 vssd1 vccd1 vccd1 _21676_/Y sky130_fd_sc_hd__nor2_1
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23415_ _23544_/CLK _23415_/D vssd1 vssd1 vccd1 vccd1 _23415_/Q sky130_fd_sc_hd__dfxtp_1
X_20627_ _23726_/Q _20593_/X _20626_/X _20602_/X vssd1 vssd1 vccd1 vccd1 _23726_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_326_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23346_ _23535_/CLK _23346_/D vssd1 vssd1 vccd1 vccd1 _23346_/Q sky130_fd_sc_hd__dfxtp_1
X_11360_ _12594_/A vssd1 vssd1 vccd1 vccd1 _12156_/A sky130_fd_sc_hd__buf_6
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20558_ _20558_/A _20558_/B _20591_/A vssd1 vssd1 vccd1 vccd1 _20558_/X sky130_fd_sc_hd__or3_1
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_355_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_353_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11291_ _12506_/A vssd1 vssd1 vccd1 vccd1 _12321_/A sky130_fd_sc_hd__buf_2
XFILLER_106_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23277_ _23534_/CLK _23277_/D vssd1 vssd1 vccd1 vccd1 _23277_/Q sky130_fd_sc_hd__dfxtp_1
X_20489_ _23715_/Q _20491_/B vssd1 vssd1 vccd1 vccd1 _20489_/X sky130_fd_sc_hd__or2_1
XFILLER_180_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13030_ _13592_/A _13027_/X _13029_/Y vssd1 vssd1 vccd1 vccd1 _13030_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_341_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22228_ _22207_/A _22207_/B _22206_/A vssd1 vssd1 vccd1 vccd1 _22232_/A sky130_fd_sc_hd__o21a_1
XFILLER_279_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22159_ _22165_/A _22044_/X _22158_/X _22048_/X vssd1 vssd1 vccd1 vccd1 _22161_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_79_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14981_ _22982_/Q _14137_/A _15164_/A input241/X vssd1 vssd1 vccd1 vccd1 _21437_/A
+ sky130_fd_sc_hd__a22o_4
XTAP_6899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16720_ _16723_/A _16720_/B vssd1 vssd1 vccd1 vccd1 _16721_/A sky130_fd_sc_hd__or2_1
XFILLER_219_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13932_ _13918_/X _15123_/A _13931_/Y _13924_/X vssd1 vssd1 vccd1 vccd1 _14093_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_304_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16651_ _22473_/Q _16268_/X _16651_/S vssd1 vssd1 vccd1 vccd1 _16652_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13863_ _13863_/A _13863_/B vssd1 vssd1 vccd1 vccd1 _13863_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_506 _15377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12814_ _12742_/A _12807_/Y _12813_/Y vssd1 vssd1 vccd1 vccd1 _12814_/X sky130_fd_sc_hd__a21o_1
X_15602_ _23701_/Q _15592_/X _15601_/X vssd1 vssd1 vccd1 vccd1 _15602_/X sky130_fd_sc_hd__o21a_4
XINSDIODE2_517 _22512_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19370_ _23346_/Q _18814_/X _19372_/S vssd1 vssd1 vccd1 vccd1 _19371_/A sky130_fd_sc_hd__mux2_1
X_16582_ _15785_/X _22442_/Q _16590_/S vssd1 vssd1 vccd1 vccd1 _16583_/A sky130_fd_sc_hd__mux2_1
XFILLER_290_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13794_ _13790_/X _13842_/A _13792_/Y _13840_/A vssd1 vssd1 vccd1 vccd1 _14043_/C
+ sky130_fd_sc_hd__a211o_4
XINSDIODE2_528 _14024_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_539 _23915_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18321_ _19932_/A vssd1 vssd1 vccd1 vccd1 _18358_/A sky130_fd_sc_hd__buf_2
X_12745_ _12745_/A vssd1 vssd1 vccd1 vccd1 _12745_/X sky130_fd_sc_hd__buf_6
XFILLER_231_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15533_ _15187_/A _15109_/B _15484_/B vssd1 vssd1 vccd1 vccd1 _15533_/Y sky130_fd_sc_hd__o21ai_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ _22864_/Q _18242_/X _18251_/X _18245_/X vssd1 vssd1 vccd1 vccd1 _22912_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15464_ _15436_/X _17122_/A _15463_/X vssd1 vssd1 vccd1 vccd1 _15464_/X sky130_fd_sc_hd__o21a_1
X_12676_ _22473_/Q _22633_/Q _12920_/A vssd1 vssd1 vccd1 vccd1 _12676_/X sky130_fd_sc_hd__mux2_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_336_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17203_ _16989_/X _15767_/X _17170_/B _23481_/Q _17202_/Y vssd1 vssd1 vccd1 vccd1
+ _17203_/X sky130_fd_sc_hd__a221o_1
X_14415_ _23909_/Q _14552_/B _14415_/S vssd1 vssd1 vccd1 vccd1 _14458_/A sky130_fd_sc_hd__mux2_1
XFILLER_318_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11627_ _12661_/A _11627_/B vssd1 vssd1 vccd1 vccd1 _11627_/Y sky130_fd_sc_hd__nand2_1
X_18183_ _18163_/A _18171_/X _18180_/X _18182_/Y _18198_/A vssd1 vssd1 vccd1 vccd1
+ _18183_/X sky130_fd_sc_hd__a221o_1
X_15395_ _22958_/Q _15726_/B vssd1 vssd1 vccd1 vccd1 _15395_/X sky130_fd_sc_hd__or2_1
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_329_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17134_ _17134_/A vssd1 vssd1 vccd1 vccd1 _17134_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14346_ _14635_/A vssd1 vssd1 vccd1 vccd1 _14841_/S sky130_fd_sc_hd__buf_2
XFILLER_317_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11558_ _11558_/A _11558_/B vssd1 vssd1 vccd1 vccd1 _13318_/A sky130_fd_sc_hd__nor2_2
XFILLER_155_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17065_ _13931_/B _17064_/X _17087_/S vssd1 vssd1 vccd1 vccd1 _17065_/X sky130_fd_sc_hd__mux2_1
X_14277_ _14348_/A _12602_/A _14276_/X vssd1 vssd1 vccd1 vccd1 _14277_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_109_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11489_ _13306_/A _11489_/B vssd1 vssd1 vccd1 vccd1 _11489_/Y sky130_fd_sc_hd__nand2_1
XFILLER_171_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_332_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16016_ _16016_/A vssd1 vssd1 vccd1 vccd1 _21077_/A sky130_fd_sc_hd__buf_8
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13228_ _23485_/Q _23581_/Q _22545_/Q _22349_/Q _11517_/A _11527_/A vssd1 vssd1 vccd1
+ vccd1 _13229_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _23486_/Q _23582_/Q _22546_/Q _22350_/Q _11431_/A _13085_/X vssd1 vssd1 vccd1
+ vccd1 _13159_/X sky130_fd_sc_hd__mux4_1
XFILLER_297_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17967_ _22832_/Q _17956_/X _17959_/X input278/X _17966_/X vssd1 vssd1 vccd1 vccd1
+ _17967_/X sky130_fd_sc_hd__a221o_1
XFILLER_285_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19706_ _19172_/X _23495_/Q _19710_/S vssd1 vssd1 vccd1 vccd1 _19707_/A sky130_fd_sc_hd__mux2_1
X_16918_ _22421_/Q _16534_/B _14160_/X _16917_/Y vssd1 vssd1 vccd1 vccd1 _16918_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_214_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17898_ _17983_/A vssd1 vssd1 vccd1 vccd1 _17933_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_266_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_19637_ _19637_/A vssd1 vssd1 vccd1 vccd1 _23464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_254_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16849_ _16847_/X _22531_/Q _16861_/S vssd1 vssd1 vccd1 vccd1 _16850_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19568_ _19625_/S vssd1 vssd1 vccd1 vccd1 _19577_/S sky130_fd_sc_hd__buf_4
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18519_ _18507_/X _18518_/Y _18516_/X vssd1 vssd1 vccd1 vccd1 _23002_/D sky130_fd_sc_hd__a21oi_1
XFILLER_209_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19499_ _19185_/X _23403_/Q _19505_/S vssd1 vssd1 vccd1 vccd1 _19500_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21530_ _23820_/Q vssd1 vssd1 vccd1 vccd1 _21530_/Y sky130_fd_sc_hd__inv_2
XFILLER_221_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_355_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21461_ _21417_/A _21416_/A _21415_/Y vssd1 vssd1 vccd1 vccd1 _21462_/B sky130_fd_sc_hd__o21a_2
XFILLER_309_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_336_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23200_ _23264_/CLK _23200_/D vssd1 vssd1 vccd1 vccd1 _23200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20412_ _20543_/A _20408_/X _20411_/X _20392_/X vssd1 vssd1 vccd1 vccd1 _23685_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21392_ _21342_/A _21342_/B _21345_/A vssd1 vssd1 vccd1 vccd1 _21393_/B sky130_fd_sc_hd__a21oi_1
XFILLER_309_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23131_ _23549_/CLK _23131_/D vssd1 vssd1 vccd1 vccd1 _23131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20343_ _20294_/X _22003_/A _20341_/Y _20342_/X vssd1 vssd1 vccd1 vccd1 _20713_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_311_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23062_ _23574_/CLK _23062_/D vssd1 vssd1 vccd1 vccd1 _23062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_289_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20274_ _17122_/A _20295_/A _20275_/B vssd1 vssd1 vccd1 vccd1 _20274_/Y sky130_fd_sc_hd__o21ai_1
XTAP_6107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22013_ _22013_/A vssd1 vssd1 vccd1 vccd1 _22231_/A sky130_fd_sc_hd__buf_2
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput206 localMemory_wb_adr_i[2] vssd1 vssd1 vccd1 vccd1 input206/X sky130_fd_sc_hd__clkbuf_1
Xinput217 localMemory_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input217/X sky130_fd_sc_hd__buf_6
XTAP_5428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput228 localMemory_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 input228/X sky130_fd_sc_hd__buf_8
XTAP_5439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput239 localMemory_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 input239/X sky130_fd_sc_hd__buf_8
XFILLER_271_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22915_ _23599_/CLK _22915_/D vssd1 vssd1 vccd1 vccd1 _22915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_272_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23895_ _23895_/CLK _23895_/D vssd1 vssd1 vccd1 vccd1 _23895_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_245_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22846_ _23426_/CLK _22846_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22777_ _23555_/CLK _22777_/D vssd1 vssd1 vccd1 vccd1 _22777_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _11127_/A _12523_/Y _12525_/Y _12527_/Y _12529_/Y vssd1 vssd1 vccd1 vccd1
+ _12530_/X sky130_fd_sc_hd__o32a_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21728_ _23794_/Q _21683_/X _21727_/Y _21346_/X vssd1 vssd1 vccd1 vccd1 _21729_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_223_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23541_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12461_ _12534_/A _12456_/Y _12458_/Y _12460_/Y vssd1 vssd1 vccd1 vccd1 _12461_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_200_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21659_ _21658_/A _21658_/B _14713_/C vssd1 vssd1 vccd1 vccd1 _21659_/X sky130_fd_sc_hd__o21a_1
XFILLER_200_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14200_ _20549_/A vssd1 vssd1 vccd1 vccd1 _14200_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_296_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11412_ _12457_/S vssd1 vssd1 vccd1 vccd1 _11413_/A sky130_fd_sc_hd__buf_4
X_15180_ _15180_/A _15483_/B vssd1 vssd1 vccd1 vccd1 _15181_/A sky130_fd_sc_hd__nor2_1
X_12392_ _23914_/Q vssd1 vssd1 vccd1 vccd1 _13901_/A sky130_fd_sc_hd__inv_2
XFILLER_342_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14131_ _14433_/S vssd1 vssd1 vccd1 vccd1 _20191_/A sky130_fd_sc_hd__buf_4
XFILLER_126_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23329_ _23553_/CLK _23329_/D vssd1 vssd1 vccd1 vccd1 _23329_/Q sky130_fd_sc_hd__dfxtp_1
X_11343_ _11343_/A _11343_/B vssd1 vssd1 vccd1 vccd1 _11343_/X sky130_fd_sc_hd__or2_1
XFILLER_315_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_314_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14062_ input233/X _14058_/X _14061_/X vssd1 vssd1 vccd1 vccd1 _14062_/X sky130_fd_sc_hd__a21bo_4
XFILLER_165_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11274_ _11683_/A vssd1 vssd1 vccd1 vccd1 _11275_/A sky130_fd_sc_hd__buf_4
XFILLER_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13013_ _13013_/A vssd1 vssd1 vccd1 vccd1 _13015_/A sky130_fd_sc_hd__inv_2
XFILLER_3_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18870_ _18870_/A vssd1 vssd1 vccd1 vccd1 _23139_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_315_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17821_ _17821_/A vssd1 vssd1 vccd1 vccd1 _22783_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_294_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17752_ _22753_/Q _17572_/X _17754_/S vssd1 vssd1 vccd1 vccd1 _17753_/A sky130_fd_sc_hd__mux2_1
XFILLER_310_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14964_ _15056_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _15380_/A sky130_fd_sc_hd__nand2_1
XTAP_5984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16703_ _22490_/Q _16689_/X _16693_/X input35/X vssd1 vssd1 vccd1 vccd1 _16704_/B
+ sky130_fd_sc_hd__o22a_1
X_13915_ _13910_/X _13913_/Y _13951_/A vssd1 vssd1 vccd1 vccd1 _13991_/B sky130_fd_sc_hd__mux2_8
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17683_ _17683_/A vssd1 vssd1 vccd1 vccd1 _22722_/D sky130_fd_sc_hd__clkbuf_1
X_14895_ _14895_/A vssd1 vssd1 vccd1 vccd1 _22264_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19422_ _23369_/Q _18785_/X _19422_/S vssd1 vssd1 vccd1 vccd1 _19423_/A sky130_fd_sc_hd__mux2_1
XFILLER_263_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_303 _15990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16634_ _22465_/Q _16243_/X _16640_/S vssd1 vssd1 vccd1 vccd1 _16635_/A sky130_fd_sc_hd__mux2_1
X_13846_ _13746_/X _13711_/B _13863_/B vssd1 vssd1 vccd1 vccd1 _13846_/Y sky130_fd_sc_hd__a21oi_1
XINSDIODE2_314 _22139_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_325 _16107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_336 _17084_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_347 _21975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19353_ _23338_/Q _18788_/X _19361_/S vssd1 vssd1 vccd1 vccd1 _19354_/A sky130_fd_sc_hd__mux2_1
XFILLER_250_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16565_ _16565_/A vssd1 vssd1 vccd1 vccd1 _22434_/D sky130_fd_sc_hd__clkbuf_1
X_13777_ _13777_/A _13777_/B vssd1 vssd1 vccd1 vccd1 _13875_/B sky130_fd_sc_hd__nor2_2
XINSDIODE2_358 INSDIODE2_358/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_369 _23476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18304_ _18305_/A _18305_/C _22928_/Q vssd1 vssd1 vccd1 vccd1 _18306_/B sky130_fd_sc_hd__a21oi_1
XFILLER_188_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15516_ _15676_/A _21240_/A _15515_/X _15775_/A vssd1 vssd1 vccd1 vccd1 _15516_/X
+ sky130_fd_sc_hd__o22a_1
X_12728_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12728_/X sky130_fd_sc_hd__buf_4
X_19284_ _19284_/A vssd1 vssd1 vccd1 vccd1 _23307_/D sky130_fd_sc_hd__clkbuf_1
X_16496_ _15625_/X _22405_/Q _16502_/S vssd1 vssd1 vccd1 vccd1 _16497_/A sky130_fd_sc_hd__mux2_1
XFILLER_337_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18235_ hold6/X _18229_/X _18234_/X _18232_/X vssd1 vssd1 vccd1 vccd1 _22905_/D sky130_fd_sc_hd__o211a_1
XFILLER_148_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12659_ _12651_/Y _12653_/Y _12655_/Y _12658_/Y _11559_/A vssd1 vssd1 vccd1 vccd1
+ _12660_/C sky130_fd_sc_hd__o221a_1
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15447_ _23826_/Q _15211_/A _15442_/X _15446_/X _14923_/A vssd1 vssd1 vccd1 vccd1
+ _15447_/X sky130_fd_sc_hd__a221o_2
X_18166_ _18181_/A _18166_/B vssd1 vssd1 vccd1 vccd1 _18179_/A sky130_fd_sc_hd__nor2_1
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15378_ _15329_/A _15376_/C _15377_/X vssd1 vssd1 vccd1 vccd1 _15379_/B sky130_fd_sc_hd__a21oi_1
XFILLER_345_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_345_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17117_ _15377_/X _17116_/X _17137_/S vssd1 vssd1 vccd1 vccd1 _17117_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14329_ _11691_/B _12168_/B _14329_/S vssd1 vssd1 vccd1 vccd1 _14329_/X sky130_fd_sc_hd__mux2_1
X_18097_ _18097_/A vssd1 vssd1 vccd1 vccd1 _18097_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_239_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_289_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17048_ _16951_/X _17046_/X _17078_/A _16996_/X vssd1 vssd1 vccd1 vccd1 _17048_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_332_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18999_ _16889_/X _23196_/Q _19001_/S vssd1 vssd1 vccd1 vccd1 _19000_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_18 _17483_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_29 _21220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20961_ _23803_/Q _20953_/X _20960_/X _20948_/X vssd1 vssd1 vccd1 vccd1 _23803_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22700_ _22801_/CLK _22700_/D vssd1 vssd1 vccd1 vccd1 _22700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23680_ _23684_/CLK _23680_/D vssd1 vssd1 vccd1 vccd1 _23680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20892_ _20969_/A vssd1 vssd1 vccd1 vccd1 _20925_/A sky130_fd_sc_hd__buf_2
XFILLER_241_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22631_ _22632_/CLK _22631_/D vssd1 vssd1 vccd1 vccd1 _22631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22562_ _22600_/CLK _22562_/D vssd1 vssd1 vccd1 vccd1 _22562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_356_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21513_ _21513_/A _21513_/B vssd1 vssd1 vccd1 vccd1 _21514_/B sky130_fd_sc_hd__nor2_1
XFILLER_186_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22493_ _23876_/CLK _22493_/D vssd1 vssd1 vccd1 vccd1 _22493_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_309_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21444_ _21444_/A _21716_/B vssd1 vssd1 vccd1 vccd1 _21444_/Y sky130_fd_sc_hd__nor2_1
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_324_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_309_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_308_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21375_ _21301_/B _21289_/A _20774_/A _21191_/A vssd1 vssd1 vccd1 vccd1 _21634_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_134_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23114_ _23370_/CLK _23114_/D vssd1 vssd1 vccd1 vccd1 _23114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_323_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20326_ _20387_/B vssd1 vssd1 vccd1 vccd1 _20400_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23045_ _23555_/CLK _23045_/D vssd1 vssd1 vccd1 vccd1 _23045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20257_ _20275_/A _20255_/Y _20320_/A vssd1 vssd1 vccd1 vccd1 _20257_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20188_ _15671_/X _21386_/A _20197_/S vssd1 vssd1 vccd1 vccd1 _20190_/B sky130_fd_sc_hd__mux2_1
XTAP_5247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ _11961_/A vssd1 vssd1 vccd1 vccd1 _12056_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _13715_/A _13985_/B _13793_/B vssd1 vssd1 vccd1 vccd1 _13701_/A sky130_fd_sc_hd__and3_4
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14680_ _14682_/A vssd1 vssd1 vccd1 vccd1 _20138_/B sky130_fd_sc_hd__buf_6
XFILLER_244_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11892_ _11723_/A _11891_/X _11706_/X vssd1 vssd1 vccd1 vccd1 _11892_/Y sky130_fd_sc_hd__o21ai_1
X_23878_ _23878_/CLK _23878_/D vssd1 vssd1 vccd1 vccd1 _23878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_352_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13631_ _23931_/Q vssd1 vssd1 vccd1 vccd1 _21950_/A sky130_fd_sc_hd__buf_4
XFILLER_71_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22829_ _22830_/CLK _22829_/D vssd1 vssd1 vccd1 vccd1 _22829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16350_ _16350_/A vssd1 vssd1 vccd1 vccd1 _22341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13562_ _13562_/A _13562_/B vssd1 vssd1 vccd1 vccd1 _13562_/Y sky130_fd_sc_hd__nand2_1
XFILLER_358_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_319_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_358_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15301_ _19977_/B _14901_/X _14902_/X _23631_/Q vssd1 vssd1 vccd1 vccd1 _15301_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_200_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12513_ _23896_/Q _12512_/X _11280_/A vssd1 vssd1 vccd1 vccd1 _12513_/X sky130_fd_sc_hd__o21a_1
X_16281_ _18846_/A vssd1 vssd1 vccd1 vccd1 _16281_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13493_ _13493_/A _13493_/B vssd1 vssd1 vccd1 vccd1 _13493_/Y sky130_fd_sc_hd__nand2_2
XFILLER_346_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18020_ _18053_/A vssd1 vssd1 vccd1 vccd1 _18020_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_200_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15232_ _14215_/X _21225_/A _15231_/X _14882_/X vssd1 vssd1 vccd1 vccd1 _15232_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_12444_ _13364_/A _14294_/A vssd1 vssd1 vccd1 vccd1 _13897_/A sky130_fd_sc_hd__xnor2_4
XFILLER_139_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15163_ _14819_/X _15157_/X _15161_/Y _15162_/X vssd1 vssd1 vccd1 vccd1 _15163_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_342_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12375_ _23464_/Q _23560_/Q _22524_/Q _22328_/Q _11646_/A _11651_/A vssd1 vssd1 vccd1
+ vccd1 _12375_/X sky130_fd_sc_hd__mux4_2
XFILLER_165_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14114_ _22886_/Q _22885_/Q vssd1 vssd1 vccd1 vccd1 _14119_/D sky130_fd_sc_hd__and2_1
XFILLER_126_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11326_ _13278_/A _11326_/B vssd1 vssd1 vccd1 vccd1 _11326_/X sky130_fd_sc_hd__or2_1
XFILLER_153_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19971_ _23605_/Q _19971_/B _19971_/C _19971_/D vssd1 vssd1 vccd1 vccd1 _19980_/C
+ sky130_fd_sc_hd__and4_1
X_15094_ _16057_/A _15092_/X _15093_/X vssd1 vssd1 vccd1 vccd1 _15094_/X sky130_fd_sc_hd__o21ba_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_326_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18922_ _18922_/A vssd1 vssd1 vccd1 vccd1 _23161_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_330_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14045_ _14023_/X _13801_/B _14041_/X input224/X vssd1 vssd1 vccd1 vccd1 _14045_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11257_ _12801_/A vssd1 vssd1 vccd1 vccd1 _11398_/A sky130_fd_sc_hd__clkbuf_8
XTAP_7161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18853_ _18853_/A vssd1 vssd1 vccd1 vccd1 _18866_/S sky130_fd_sc_hd__buf_6
XTAP_6460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11188_ _11424_/A _11188_/B vssd1 vssd1 vccd1 vccd1 _11188_/Y sky130_fd_sc_hd__nor2_1
XFILLER_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_311_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17804_ _19267_/A _17804_/B vssd1 vssd1 vccd1 vccd1 _17861_/A sky130_fd_sc_hd__nor2_8
XFILLER_39_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18784_ _18784_/A vssd1 vssd1 vccd1 vccd1 _23112_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15996_ _15996_/A _15996_/B vssd1 vssd1 vccd1 vccd1 _15996_/Y sky130_fd_sc_hd__nand2_1
XFILLER_342_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_294_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17735_ _22745_/Q _17544_/X _17743_/S vssd1 vssd1 vccd1 vccd1 _17736_/A sky130_fd_sc_hd__mux2_1
XFILLER_342_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14947_ _15456_/A _14855_/B _14767_/X vssd1 vssd1 vccd1 vccd1 _14947_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17666_ _17666_/A vssd1 vssd1 vccd1 vccd1 _22714_/D sky130_fd_sc_hd__clkbuf_1
X_14878_ _22917_/Q _14509_/X _14513_/X _22949_/Q vssd1 vssd1 vccd1 vccd1 _14878_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_223_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_100 _21648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_111 _13875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19405_ _23362_/Q _18865_/X _19405_/S vssd1 vssd1 vccd1 vccd1 _19406_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_122 _13714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16617_ _16617_/A vssd1 vssd1 vccd1 vccd1 _22457_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_133 _13500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13829_ _15576_/A _13829_/B vssd1 vssd1 vccd1 vccd1 _13874_/C sky130_fd_sc_hd__or2_2
XINSDIODE2_144 _21448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17597_ _17597_/A vssd1 vssd1 vccd1 vccd1 _22693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_250_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_155 _14866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_166 _13633_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19336_ _19336_/A vssd1 vssd1 vccd1 vccd1 _23331_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_177 _13701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_188 _13991_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16548_ _16605_/S vssd1 vssd1 vccd1 vccd1 _16557_/S sky130_fd_sc_hd__buf_6
XFILLER_287_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_199 _13951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19267_ _19267_/A _19771_/B vssd1 vssd1 vccd1 vccd1 _19324_/A sky130_fd_sc_hd__or2_4
XFILLER_149_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16479_ _16479_/A vssd1 vssd1 vccd1 vccd1 _22397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_337_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18218_ _22899_/Q _18227_/B vssd1 vssd1 vccd1 vccd1 _18218_/X sky130_fd_sc_hd__or2_1
XFILLER_164_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19198_ _19265_/S vssd1 vssd1 vccd1 vccd1 _19211_/S sky130_fd_sc_hd__buf_4
XFILLER_306_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18149_ _22886_/Q _22879_/Q _18158_/S vssd1 vssd1 vccd1 vccd1 _18150_/B sky130_fd_sc_hd__mux2_1
XFILLER_156_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_333_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21160_ _23868_/Q _21139_/X _21159_/X _21073_/X vssd1 vssd1 vccd1 vccd1 _23868_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20111_ _23644_/Q _20123_/C vssd1 vssd1 vccd1 vccd1 _20114_/B sky130_fd_sc_hd__nor2_1
XFILLER_131_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21091_ _21091_/A _21091_/B vssd1 vssd1 vccd1 vccd1 _23846_/D sky130_fd_sc_hd__nor2_1
XFILLER_160_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_302_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20042_ _23624_/Q _20048_/B _20042_/C _20042_/D vssd1 vssd1 vccd1 vccd1 _20051_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23801_ _23942_/CLK _23801_/D vssd1 vssd1 vccd1 vccd1 _23801_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21993_ _21993_/A _21993_/B vssd1 vssd1 vccd1 vccd1 _21995_/A sky130_fd_sc_hd__nor2_1
XFILLER_227_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23732_ _23918_/CLK _23732_/D vssd1 vssd1 vccd1 vccd1 _23732_/Q sky130_fd_sc_hd__dfxtp_1
X_20944_ _23797_/Q _20939_/X _20943_/X _20934_/X vssd1 vssd1 vccd1 vccd1 _23797_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23663_ _23818_/CLK _23663_/D vssd1 vssd1 vccd1 vccd1 _23663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20875_ _20747_/B _20864_/X _20865_/X _23776_/Q vssd1 vssd1 vccd1 vccd1 _20876_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22614_ _23527_/CLK _22614_/D vssd1 vssd1 vccd1 vccd1 _22614_/Q sky130_fd_sc_hd__dfxtp_1
X_23594_ _23600_/CLK _23594_/D vssd1 vssd1 vccd1 vccd1 _23594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_356_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22545_ _23547_/CLK _22545_/D vssd1 vssd1 vccd1 vccd1 _22545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_324_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22476_ _23577_/CLK _22476_/D vssd1 vssd1 vccd1 vccd1 _22476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21427_ _21344_/A _21344_/B _21425_/X _21391_/B _21426_/X vssd1 vssd1 vccd1 vccd1
+ _21428_/B sky130_fd_sc_hd__a311o_2
XFILLER_324_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12160_ _12160_/A _13497_/A vssd1 vssd1 vccd1 vccd1 _13342_/A sky130_fd_sc_hd__nor2_2
XFILLER_108_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21358_ _23815_/Q _23749_/Q _21456_/A vssd1 vssd1 vccd1 vccd1 _21361_/B sky130_fd_sc_hd__and3_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11111_ _11146_/A vssd1 vssd1 vccd1 vccd1 _11112_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_151_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20309_ _23670_/Q _20338_/B vssd1 vssd1 vccd1 vccd1 _20309_/X sky130_fd_sc_hd__or2_1
XFILLER_311_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12091_ _12091_/A _12091_/B vssd1 vssd1 vccd1 vccd1 _12091_/X sky130_fd_sc_hd__or2_1
X_21289_ _21289_/A _21289_/B vssd1 vssd1 vccd1 vccd1 _21297_/C sky130_fd_sc_hd__and2_1
XFILLER_249_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23028_ _23414_/CLK _23028_/D vssd1 vssd1 vccd1 vccd1 _23028_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15850_ _16034_/A _15850_/B vssd1 vssd1 vccd1 vccd1 _15850_/X sky130_fd_sc_hd__or2_1
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14801_ _14801_/A vssd1 vssd1 vccd1 vccd1 _15345_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15781_ _15781_/A vssd1 vssd1 vccd1 vccd1 _15932_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_218_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _12993_/A _12993_/B vssd1 vssd1 vccd1 vccd1 _12993_/X sky130_fd_sc_hd__or2_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _17520_/A vssd1 vssd1 vccd1 vccd1 _22666_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14732_ _14901_/A vssd1 vssd1 vccd1 vccd1 _14732_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_312_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_291_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11944_ _11944_/A vssd1 vssd1 vccd1 vccd1 _13521_/B sky130_fd_sc_hd__buf_4
XFILLER_206_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17451_ _17451_/A vssd1 vssd1 vccd1 vccd1 _22636_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14663_ _14340_/X _14342_/X _14664_/S vssd1 vssd1 vccd1 vccd1 _14663_/X sky130_fd_sc_hd__mux2_1
X_11875_ _12410_/A _11875_/B vssd1 vssd1 vccd1 vccd1 _11875_/X sky130_fd_sc_hd__or2_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16402_ _16402_/A vssd1 vssd1 vccd1 vccd1 _22363_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13614_ _15492_/S _13619_/A vssd1 vssd1 vccd1 vccd1 _13615_/B sky130_fd_sc_hd__nor2_2
XFILLER_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17382_ _17382_/A vssd1 vssd1 vccd1 vccd1 _20808_/A sky130_fd_sc_hd__inv_2
X_14594_ _19922_/B _14450_/X _14455_/X _23622_/Q vssd1 vssd1 vccd1 vccd1 _14594_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_198_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19121_ _19121_/A vssd1 vssd1 vccd1 vccd1 _23249_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16333_ _15283_/X _22334_/Q _16333_/S vssd1 vssd1 vccd1 vccd1 _16334_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13545_ _13080_/A _13542_/Y _13544_/Y _13082_/B vssd1 vssd1 vccd1 vccd1 _13545_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_185_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19052_ _19052_/A vssd1 vssd1 vccd1 vccd1 _23219_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16264_ _16264_/A vssd1 vssd1 vccd1 vccd1 _22310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13476_ _13476_/A vssd1 vssd1 vccd1 vccd1 _13476_/Y sky130_fd_sc_hd__inv_2
XFILLER_347_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18003_ _22842_/Q _17990_/X _17986_/X _18002_/X _17933_/A vssd1 vssd1 vccd1 vccd1
+ _18003_/X sky130_fd_sc_hd__a221o_1
XFILLER_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15215_ _15215_/A vssd1 vssd1 vccd1 vccd1 _15215_/X sky130_fd_sc_hd__clkbuf_4
X_12427_ _12523_/A _12426_/X _11127_/A vssd1 vssd1 vccd1 vccd1 _12427_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_315_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16195_ _16193_/X _16194_/X _16195_/S vssd1 vssd1 vccd1 vccd1 _18871_/A sky130_fd_sc_hd__mux2_8
XFILLER_327_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput307 _13957_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[12] sky130_fd_sc_hd__buf_2
XFILLER_337_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15146_ _23820_/Q _14464_/X _15142_/X _15145_/X _14612_/X vssd1 vssd1 vccd1 vccd1
+ _15146_/X sky130_fd_sc_hd__a221o_2
Xoutput318 _13978_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[23] sky130_fd_sc_hd__buf_2
X_12358_ _23304_/Q _23272_/Q _23240_/Q _23528_/Q _11413_/A _11702_/A vssd1 vssd1 vccd1
+ vccd1 _12359_/B sky130_fd_sc_hd__mux4_2
Xoutput329 _13941_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[8] sky130_fd_sc_hd__buf_2
XFILLER_330_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_288_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_287_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_342_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_315_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11309_ _11532_/A vssd1 vssd1 vccd1 vccd1 _11517_/A sky130_fd_sc_hd__buf_4
XFILLER_4_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19954_ _19981_/A _19959_/C vssd1 vssd1 vccd1 vccd1 _19954_/Y sky130_fd_sc_hd__nor2_1
X_15077_ _15003_/X _15064_/X _15076_/X vssd1 vssd1 vccd1 vccd1 _17052_/A sky130_fd_sc_hd__o21ai_4
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12289_ _13928_/A _13920_/A vssd1 vssd1 vccd1 vccd1 _12289_/Y sky130_fd_sc_hd__nor2_1
XFILLER_206_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18905_ _23154_/Q _18814_/X _18907_/S vssd1 vssd1 vccd1 vccd1 _18906_/A sky130_fd_sc_hd__mux2_1
X_14028_ _13754_/B _14049_/A vssd1 vssd1 vccd1 vccd1 _14028_/X sky130_fd_sc_hd__and2b_1
XFILLER_302_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19885_ _16265_/X _23575_/Q _19887_/S vssd1 vssd1 vccd1 vccd1 _19886_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_295_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18836_ _18836_/A vssd1 vssd1 vccd1 vccd1 _18836_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_255_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18767_ _16914_/X _23108_/Q _18767_/S vssd1 vssd1 vccd1 vccd1 _18768_/A sky130_fd_sc_hd__mux2_1
X_15979_ _15575_/X _15287_/Y _15942_/X vssd1 vssd1 vccd1 vccd1 _21272_/A sky130_fd_sc_hd__a21oi_4
XFILLER_49_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17718_ _22738_/Q _17626_/X _17726_/S vssd1 vssd1 vccd1 vccd1 _17719_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18698_ _18754_/A vssd1 vssd1 vccd1 vccd1 _18767_/S sky130_fd_sc_hd__buf_6
XFILLER_270_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17649_ _17655_/B vssd1 vssd1 vccd1 vccd1 _17653_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_212_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20660_ _20660_/A vssd1 vssd1 vccd1 vccd1 _20661_/A sky130_fd_sc_hd__clkinv_2
XFILLER_338_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_189_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23493_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19319_ _19319_/A vssd1 vssd1 vccd1 vccd1 _23323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_338_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20591_ _20591_/A _20591_/B _20591_/C vssd1 vssd1 vccd1 vccd1 _20591_/X sky130_fd_sc_hd__or3_1
XFILLER_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_118_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23592_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22330_ _23530_/CLK _22330_/D vssd1 vssd1 vccd1 vccd1 _22330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22261_ _23903_/CLK _22261_/D vssd1 vssd1 vccd1 vccd1 _22261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_352_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21212_ _21215_/A _21212_/B vssd1 vssd1 vccd1 vccd1 _21213_/A sky130_fd_sc_hd__and2_1
XFILLER_340_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22192_ _22193_/A _22197_/A vssd1 vssd1 vccd1 vccd1 _22195_/A sky130_fd_sc_hd__nor2_1
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21143_ _20675_/A _21140_/X _21142_/X _20520_/B _21135_/X vssd1 vssd1 vccd1 vccd1
+ _21143_/X sky130_fd_sc_hd__a221o_1
XFILLER_133_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21074_ _20765_/A _21008_/A _21072_/X _21073_/X vssd1 vssd1 vccd1 vccd1 _23844_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_330_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20025_ _20041_/A _20025_/B _20025_/C vssd1 vssd1 vccd1 vccd1 _23619_/D sky130_fd_sc_hd__nor3_1
XFILLER_259_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_274_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21976_ _23932_/Q _21979_/A vssd1 vssd1 vccd1 vccd1 _21977_/B sky130_fd_sc_hd__or2_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23715_ _23871_/CLK _23715_/D vssd1 vssd1 vccd1 vccd1 _23715_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20927_ _13951_/B _20922_/X _20635_/B _20926_/X vssd1 vssd1 vccd1 vccd1 _20927_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_270_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _12334_/A vssd1 vssd1 vccd1 vccd1 _12406_/A sky130_fd_sc_hd__clkbuf_4
X_23646_ _23646_/CLK _23646_/D vssd1 vssd1 vccd1 vccd1 _23646_/Q sky130_fd_sc_hd__dfxtp_1
X_20858_ _20861_/A _20858_/B vssd1 vssd1 vccd1 vccd1 _20859_/A sky130_fd_sc_hd__and2_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_357_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11591_ _12073_/A vssd1 vssd1 vccd1 vccd1 _12041_/A sky130_fd_sc_hd__buf_4
XFILLER_211_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23577_ _23577_/CLK _23577_/D vssd1 vssd1 vccd1 vccd1 _23577_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_288_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20789_ _20888_/C _20785_/X _20786_/X _20788_/X vssd1 vssd1 vccd1 vccd1 _23752_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_357_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13330_ _13532_/D _13330_/B vssd1 vssd1 vccd1 vccd1 _13387_/A sky130_fd_sc_hd__xnor2_4
XFILLER_195_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22528_ _23500_/CLK _22528_/D vssd1 vssd1 vccd1 vccd1 _22528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_298_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_316_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13261_ _13268_/A _13260_/X _11236_/X vssd1 vssd1 vccd1 vccd1 _13261_/Y sky130_fd_sc_hd__o21ai_1
X_22459_ _23368_/CLK _22459_/D vssd1 vssd1 vccd1 vccd1 _22459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15000_ _15000_/A vssd1 vssd1 vccd1 vccd1 _15000_/X sky130_fd_sc_hd__clkbuf_2
X_12212_ _12387_/A _12211_/X _11819_/A vssd1 vssd1 vccd1 vccd1 _12212_/X sky130_fd_sc_hd__o21a_1
XFILLER_142_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13192_ _11195_/A _13191_/X _13091_/A vssd1 vssd1 vccd1 vccd1 _13192_/X sky130_fd_sc_hd__a21o_1
XFILLER_182_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12143_ _23409_/Q _23025_/Q _23377_/Q _23345_/Q _11637_/A _11742_/A vssd1 vssd1 vccd1
+ vccd1 _12144_/B sky130_fd_sc_hd__mux4_1
XFILLER_151_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16951_ _16951_/A vssd1 vssd1 vccd1 vccd1 _16951_/X sky130_fd_sc_hd__clkbuf_2
X_12074_ _22790_/Q _22758_/Q _22659_/Q _22726_/Q _11894_/S _11566_/A vssd1 vssd1 vccd1
+ vccd1 _12074_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15902_ _15633_/X _15189_/Y _15942_/A vssd1 vssd1 vccd1 vccd1 _21267_/A sky130_fd_sc_hd__a21oi_4
X_19670_ _19670_/A vssd1 vssd1 vccd1 vccd1 _23479_/D sky130_fd_sc_hd__clkbuf_1
X_16882_ _16882_/A vssd1 vssd1 vccd1 vccd1 _22541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_265_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_293_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18621_ _16911_/X _23043_/Q _18623_/S vssd1 vssd1 vccd1 vccd1 _18622_/A sky130_fd_sc_hd__mux2_1
X_15833_ _22936_/Q vssd1 vssd1 vccd1 vccd1 _15833_/X sky130_fd_sc_hd__buf_2
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18552_ _19090_/B _18770_/B _17471_/B vssd1 vssd1 vccd1 vccd1 _19483_/B sky130_fd_sc_hd__or3b_4
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _22966_/Q _15763_/X _16144_/S vssd1 vssd1 vccd1 vccd1 _15764_/X sky130_fd_sc_hd__mux2_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _22799_/Q _22767_/Q _22668_/Q _22735_/Q _12921_/S _12749_/X vssd1 vssd1 vccd1
+ vccd1 _12976_/X sky130_fd_sc_hd__mux4_2
XFILLER_205_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_346_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17503_ _22659_/Q _16249_/X _17505_/S vssd1 vssd1 vccd1 vccd1 _17504_/A sky130_fd_sc_hd__mux2_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ input134/X input129/X _15033_/S vssd1 vssd1 vccd1 vccd1 _14715_/X sky130_fd_sc_hd__mux2_8
XFILLER_233_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18483_ _18480_/X _18482_/Y _18476_/X vssd1 vssd1 vccd1 vccd1 _22988_/D sky130_fd_sc_hd__a21oi_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _23469_/Q _23565_/Q _22529_/Q _22333_/Q _11821_/X _11317_/A vssd1 vssd1 vccd1
+ vccd1 _11928_/B sky130_fd_sc_hd__mux4_1
X_15695_ _22932_/Q _15259_/B _15685_/X _15694_/Y _14727_/X vssd1 vssd1 vccd1 vccd1
+ _15695_/X sky130_fd_sc_hd__a221o_1
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17434_ _17456_/A vssd1 vssd1 vccd1 vccd1 _17443_/S sky130_fd_sc_hd__buf_4
XFILLER_178_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14646_ _14283_/X _14286_/X _14646_/S vssd1 vssd1 vccd1 vccd1 _14646_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11858_ _14179_/A _11910_/A vssd1 vssd1 vccd1 vccd1 _11858_/X sky130_fd_sc_hd__or2_1
XFILLER_199_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17365_ _22603_/Q input197/X _17369_/S vssd1 vssd1 vccd1 vccd1 _17366_/A sky130_fd_sc_hd__mux2_1
X_14577_ _14725_/A _15243_/A vssd1 vssd1 vccd1 vccd1 _14577_/X sky130_fd_sc_hd__or2_1
XFILLER_186_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11789_ _11905_/A _11789_/B vssd1 vssd1 vccd1 vccd1 _11789_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19104_ _19161_/S vssd1 vssd1 vccd1 vccd1 _19113_/S sky130_fd_sc_hd__buf_4
XFILLER_348_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16316_ _14706_/X _22326_/Q _16322_/S vssd1 vssd1 vccd1 vccd1 _16317_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13528_ _13528_/A _13528_/B _13528_/C vssd1 vssd1 vccd1 vccd1 _13621_/C sky130_fd_sc_hd__or3_2
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_335_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17296_ input100/X input64/X _17314_/S vssd1 vssd1 vccd1 vccd1 _17296_/X sky130_fd_sc_hd__mux2_8
XFILLER_334_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_348_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19035_ _19035_/A vssd1 vssd1 vccd1 vccd1 _23211_/D sky130_fd_sc_hd__clkbuf_1
X_16247_ _22305_/Q _16246_/X _16253_/S vssd1 vssd1 vccd1 vccd1 _16248_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_2_wb_clk_i clkbuf_1_0_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_334_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13459_ _13459_/A vssd1 vssd1 vccd1 vccd1 _14820_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_284_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_322_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16178_ _16168_/A _14752_/A _14753_/A _22977_/Q vssd1 vssd1 vccd1 vccd1 _16178_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_303_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_343_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15129_ _14851_/X _14853_/X _15129_/S vssd1 vssd1 vccd1 vccd1 _15538_/B sky130_fd_sc_hd__mux2_2
XFILLER_342_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_331_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19937_ _23596_/Q _23595_/Q _23592_/Q vssd1 vssd1 vccd1 vccd1 _19938_/C sky130_fd_sc_hd__and3_1
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_287_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19868_ _16239_/X _23567_/Q _19876_/S vssd1 vssd1 vccd1 vccd1 _19869_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18819_ _18819_/A vssd1 vssd1 vccd1 vccd1 _23123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19799_ _19799_/A vssd1 vssd1 vccd1 vccd1 _23536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_271_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21830_ _21594_/B _21828_/Y _21829_/Y _21677_/X vssd1 vssd1 vccd1 vccd1 _21831_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_83_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21761_ _21762_/A _21766_/A vssd1 vssd1 vccd1 vccd1 _21763_/A sky130_fd_sc_hd__nand2_1
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23500_ _23500_/CLK _23500_/D vssd1 vssd1 vccd1 vccd1 _23500_/Q sky130_fd_sc_hd__dfxtp_1
X_20712_ _23738_/Q _20697_/X _20711_/X _20706_/X vssd1 vssd1 vccd1 vccd1 _23738_/D
+ sky130_fd_sc_hd__o211a_1
X_21692_ _16118_/A _21550_/B _21599_/Y _21601_/Y vssd1 vssd1 vccd1 vccd1 _21692_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_357_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_339_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23431_ _23527_/CLK _23431_/D vssd1 vssd1 vccd1 vccd1 _23431_/Q sky130_fd_sc_hd__dfxtp_1
X_20643_ _14535_/X _20642_/X _20574_/X vssd1 vssd1 vccd1 vccd1 _20643_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_339_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23362_ _23489_/CLK _23362_/D vssd1 vssd1 vccd1 vccd1 _23362_/Q sky130_fd_sc_hd__dfxtp_1
X_20574_ _20733_/A vssd1 vssd1 vccd1 vccd1 _20574_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_258_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22313_ _22666_/CLK _22313_/D vssd1 vssd1 vccd1 vccd1 _22313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_325_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23293_ _23549_/CLK _23293_/D vssd1 vssd1 vccd1 vccd1 _23293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_354_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22244_ _22237_/Y _22238_/X _22243_/X vssd1 vssd1 vccd1 vccd1 _22244_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_306_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22175_ _22166_/A _21366_/X _22174_/X _22122_/X vssd1 vssd1 vccd1 vccd1 _23939_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_86_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _22801_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21126_ _21134_/A _21126_/B vssd1 vssd1 vccd1 vccd1 _23857_/D sky130_fd_sc_hd__nor2_1
XFILLER_105_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23503_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_293_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21057_ _20723_/A _21047_/X _21056_/X _21049_/X vssd1 vssd1 vccd1 vccd1 _23837_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20008_ _20008_/A _20008_/B _20021_/C vssd1 vssd1 vccd1 vccd1 _23614_/D sky130_fd_sc_hd__nor3_1
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12830_ _12836_/A _12830_/B vssd1 vssd1 vccd1 vccd1 _12830_/Y sky130_fd_sc_hd__nor2_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _22375_/Q _22407_/Q _22696_/Q _23063_/Q _12922_/S _12746_/X vssd1 vssd1 vccd1
+ vccd1 _12761_/X sky130_fd_sc_hd__mux4_2
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21959_ _20334_/A _22045_/A _15793_/B _22046_/A vssd1 vssd1 vccd1 vccd1 _21959_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_70_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14500_ _14500_/A _14510_/B _15068_/C vssd1 vssd1 vccd1 vccd1 _15726_/B sky130_fd_sc_hd__or3_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11712_ _22788_/Q _22756_/Q _22657_/Q _22724_/Q _11700_/X _11590_/A vssd1 vssd1 vccd1
+ vccd1 _11712_/X sky130_fd_sc_hd__mux4_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12755_/A vssd1 vssd1 vccd1 vccd1 _12692_/X sky130_fd_sc_hd__buf_4
XFILLER_230_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15480_ _15480_/A vssd1 vssd1 vccd1 vccd1 _15480_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_230_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11643_ _23318_/Q _23286_/Q _23254_/Q _23542_/Q _11637_/X _12777_/A vssd1 vssd1 vccd1
+ vccd1 _11643_/X sky130_fd_sc_hd__mux4_2
X_14431_ _14431_/A vssd1 vssd1 vccd1 vccd1 _14431_/X sky130_fd_sc_hd__buf_2
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23629_ _23632_/CLK _23629_/D vssd1 vssd1 vccd1 vccd1 _23629_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17150_ _17148_/X _17149_/Y _17163_/B vssd1 vssd1 vccd1 vccd1 _17150_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_174_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11574_ _11574_/A vssd1 vssd1 vccd1 vccd1 _12119_/S sky130_fd_sc_hd__buf_2
XFILLER_196_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14362_ _14949_/S vssd1 vssd1 vccd1 vccd1 _15085_/S sky130_fd_sc_hd__buf_2
XFILLER_317_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 core_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16101_ _23618_/Q _15589_/X _15590_/X _23650_/Q vssd1 vssd1 vccd1 vccd1 _16101_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput28 core_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput39 core_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_1
X_13313_ _13403_/A _13310_/X _13312_/X vssd1 vssd1 vccd1 vccd1 _14388_/C sky130_fd_sc_hd__o21ai_2
X_17081_ _22561_/Q _17038_/X _17028_/X _17080_/X vssd1 vssd1 vccd1 vccd1 _22561_/D
+ sky130_fd_sc_hd__a211o_1
X_14293_ _14285_/X _14291_/X _14635_/A vssd1 vssd1 vccd1 vccd1 _14293_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13244_ _13187_/A _13240_/Y _13243_/X vssd1 vssd1 vccd1 vccd1 _13244_/X sky130_fd_sc_hd__a21o_1
X_16032_ _13082_/B _16054_/B _14761_/A _13080_/A _14836_/A vssd1 vssd1 vccd1 vccd1
+ _16032_/X sky130_fd_sc_hd__a221o_1
XFILLER_115_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_344_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_297_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13175_ _23230_/Q _23198_/Q _23166_/Q _23134_/Q _11532_/X _13127_/X vssd1 vssd1 vccd1
+ vccd1 _13176_/B sky130_fd_sc_hd__mux4_1
XFILLER_272_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_324_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_313_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_340_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12126_ _12130_/A _12126_/B vssd1 vssd1 vccd1 vccd1 _12126_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17983_ _17983_/A vssd1 vssd1 vccd1 vccd1 _17983_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_334_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19722_ _19722_/A vssd1 vssd1 vccd1 vccd1 _23502_/D sky130_fd_sc_hd__clkbuf_1
X_12057_ _23475_/Q _23571_/Q _22535_/Q _22339_/Q _12825_/A _12756_/A vssd1 vssd1 vccd1
+ vccd1 _12057_/X sky130_fd_sc_hd__mux4_1
X_16934_ _22249_/C vssd1 vssd1 vccd1 vccd1 _16958_/B sky130_fd_sc_hd__inv_2
XFILLER_266_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19653_ _19653_/A vssd1 vssd1 vccd1 vccd1 _23471_/D sky130_fd_sc_hd__clkbuf_1
X_16865_ _16863_/X _22536_/Q _16877_/S vssd1 vssd1 vccd1 vccd1 _16866_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18604_ _16886_/X _23035_/Q _18608_/S vssd1 vssd1 vccd1 vccd1 _18605_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15816_ _15802_/X _15815_/Y _11099_/A vssd1 vssd1 vccd1 vccd1 _15816_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_350_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19584_ _23441_/Q _19204_/A _19588_/S vssd1 vssd1 vccd1 vccd1 _19585_/A sky130_fd_sc_hd__mux2_1
X_16796_ _16796_/A vssd1 vssd1 vccd1 vccd1 _22515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18535_ _18480_/A _18534_/Y _18264_/A vssd1 vssd1 vccd1 vccd1 _23009_/D sky130_fd_sc_hd__a21oi_1
XFILLER_281_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_350_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15747_ _15744_/Y _21920_/A _16047_/S vssd1 vssd1 vccd1 vccd1 _18833_/A sky130_fd_sc_hd__mux2_8
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _12993_/A _12956_/X _12958_/X _12721_/X vssd1 vssd1 vccd1 vccd1 _12959_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18466_ _18451_/X _18465_/Y _18463_/X vssd1 vssd1 vccd1 vccd1 _22982_/D sky130_fd_sc_hd__a21oi_1
XFILLER_34_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15678_ _15678_/A _15996_/B vssd1 vssd1 vccd1 vccd1 _15678_/Y sky130_fd_sc_hd__nand2_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17417_ _22621_/Q _16230_/X _17421_/S vssd1 vssd1 vccd1 vccd1 _17418_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14629_ _14629_/A vssd1 vssd1 vccd1 vccd1 _14629_/Y sky130_fd_sc_hd__inv_2
XFILLER_221_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18397_ _15501_/A _18400_/C _18380_/X vssd1 vssd1 vccd1 vccd1 _18397_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_159_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17348_ _17348_/A vssd1 vssd1 vccd1 vccd1 _22595_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_295_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_307_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17279_ _17279_/A vssd1 vssd1 vccd1 vccd1 _17279_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19018_ _19267_/A _19018_/B vssd1 vssd1 vccd1 vccd1 _19075_/A sky130_fd_sc_hd__or2_4
XFILLER_106_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_350_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20290_ _21791_/B vssd1 vssd1 vccd1 vccd1 _21790_/B sky130_fd_sc_hd__clkinv_4
XFILLER_228_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_322_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_288_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_331_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22931_ _22961_/CLK _22931_/D vssd1 vssd1 vccd1 vccd1 _22931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22862_ _23008_/CLK _22862_/D vssd1 vssd1 vccd1 vccd1 _22862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_260_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21813_ _21813_/A _21853_/B _21813_/C vssd1 vssd1 vccd1 vccd1 _21813_/X sky130_fd_sc_hd__or3_1
X_22793_ _23446_/CLK _22793_/D vssd1 vssd1 vccd1 vccd1 _22793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_133_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _22974_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_184_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21744_ _21491_/X _21735_/X _21743_/Y vssd1 vssd1 vccd1 vccd1 _21744_/X sky130_fd_sc_hd__a21o_1
XFILLER_358_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_358_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21675_ _21675_/A _21675_/B vssd1 vssd1 vccd1 vccd1 _21675_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_237_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23414_ _23414_/CLK _23414_/D vssd1 vssd1 vccd1 vccd1 _23414_/Q sky130_fd_sc_hd__dfxtp_1
X_20626_ _20626_/A _20626_/B _20626_/C vssd1 vssd1 vccd1 vccd1 _20626_/X sky130_fd_sc_hd__or3_1
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_327_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23345_ _23537_/CLK _23345_/D vssd1 vssd1 vccd1 vccd1 _23345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_338_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20557_ _20768_/A vssd1 vssd1 vccd1 vccd1 _20591_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_137_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_353_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_342_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_354_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23276_ _23950_/A _23276_/D vssd1 vssd1 vccd1 vccd1 _23276_/Q sky130_fd_sc_hd__dfxtp_1
X_11290_ _12511_/A vssd1 vssd1 vccd1 vccd1 _12506_/A sky130_fd_sc_hd__buf_2
XFILLER_342_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20488_ _20754_/A _20428_/A _20487_/X _20483_/X vssd1 vssd1 vccd1 vccd1 _23714_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_279_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22227_ _22217_/A _21366_/X _22226_/Y _22122_/X vssd1 vssd1 vccd1 vccd1 _23941_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_322_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22158_ _22046_/X _16079_/B _21900_/B _20381_/A vssd1 vssd1 vccd1 vccd1 _22158_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_6834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput490 _23918_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[7] sky130_fd_sc_hd__buf_2
XFILLER_294_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21109_ _21122_/A vssd1 vssd1 vccd1 vccd1 _21121_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_6867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14980_ _14980_/A vssd1 vssd1 vccd1 vccd1 _15164_/A sky130_fd_sc_hd__clkbuf_2
X_22089_ _22086_/X _22087_/Y _22065_/A _22085_/Y vssd1 vssd1 vccd1 vccd1 _22090_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_121_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13931_ _13931_/A _13931_/B vssd1 vssd1 vccd1 vccd1 _13931_/Y sky130_fd_sc_hd__nor2_1
XFILLER_275_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16650_ _16650_/A vssd1 vssd1 vccd1 vccd1 _22472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13862_ _13893_/A vssd1 vssd1 vccd1 vccd1 _13892_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_47_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15601_ _23829_/Q _15593_/X _15594_/X _15600_/X _14738_/X vssd1 vssd1 vccd1 vccd1
+ _15601_/X sky130_fd_sc_hd__a221o_1
XINSDIODE2_507 _15606_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12813_ _12809_/Y _12812_/Y _13599_/A vssd1 vssd1 vccd1 vccd1 _12813_/Y sky130_fd_sc_hd__a21oi_1
X_16581_ _16592_/A vssd1 vssd1 vccd1 vccd1 _16590_/S sky130_fd_sc_hd__clkbuf_4
XINSDIODE2_518 _22491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13793_ _13821_/A _13793_/B vssd1 vssd1 vccd1 vccd1 _13840_/A sky130_fd_sc_hd__nor2_1
XFILLER_216_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_529 _14026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18320_ _15724_/X _18323_/C _18319_/Y vssd1 vssd1 vccd1 vccd1 _22933_/D sky130_fd_sc_hd__o21a_1
X_15532_ _15532_/A _15485_/B vssd1 vssd1 vccd1 vccd1 _15865_/B sky130_fd_sc_hd__or2b_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _13532_/C vssd1 vssd1 vccd1 vccd1 _13599_/A sky130_fd_sc_hd__buf_4
XFILLER_215_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18251_ _22912_/Q _18253_/B vssd1 vssd1 vccd1 vccd1 _18251_/X sky130_fd_sc_hd__or2_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _15454_/X _15462_/X _14690_/A vssd1 vssd1 vccd1 vccd1 _15463_/X sky130_fd_sc_hd__a21o_1
X_12675_ _12675_/A vssd1 vssd1 vccd1 vccd1 _12920_/A sky130_fd_sc_hd__buf_4
XFILLER_230_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17202_ _17248_/A vssd1 vssd1 vccd1 vccd1 _17202_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14414_ _22906_/Q _14153_/X _14151_/X _22599_/Q vssd1 vssd1 vccd1 vccd1 _14552_/B
+ sky130_fd_sc_hd__a22o_1
X_18182_ _18162_/A _18167_/X _18165_/X _18195_/A vssd1 vssd1 vccd1 vccd1 _18182_/Y
+ sky130_fd_sc_hd__o211ai_1
X_11626_ _11559_/X _11601_/Y _11625_/X _13718_/A vssd1 vssd1 vccd1 vccd1 _11627_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_329_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15394_ _22926_/Q _14931_/A _14933_/A _22958_/Q vssd1 vssd1 vccd1 vccd1 _15394_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_345_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17133_ _21762_/A vssd1 vssd1 vccd1 vccd1 _17133_/X sky130_fd_sc_hd__buf_8
X_14345_ _14342_/X _14343_/X _14660_/S vssd1 vssd1 vccd1 vccd1 _14345_/X sky130_fd_sc_hd__mux2_1
X_11557_ _11557_/A _11557_/B vssd1 vssd1 vccd1 vccd1 _11558_/B sky130_fd_sc_hd__and2_1
XFILLER_318_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_344_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17064_ _14548_/X _17063_/X _17144_/A vssd1 vssd1 vccd1 vccd1 _17064_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_305_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14276_ _14288_/A _14276_/B vssd1 vssd1 vccd1 vccd1 _14276_/X sky130_fd_sc_hd__or2_1
X_11488_ _13306_/B vssd1 vssd1 vccd1 vccd1 _11489_/B sky130_fd_sc_hd__clkinv_2
XFILLER_109_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_345_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16015_ _16015_/A vssd1 vssd1 vccd1 vccd1 _22287_/D sky130_fd_sc_hd__clkbuf_1
X_13227_ _13218_/A _13226_/X _11537_/A vssd1 vssd1 vccd1 vccd1 _13227_/X sky130_fd_sc_hd__o21a_1
XFILLER_171_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_350_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13158_ _13158_/A _13158_/B vssd1 vssd1 vccd1 vccd1 _13158_/Y sky130_fd_sc_hd__nor2_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12109_ _12156_/A _12109_/B _12109_/C vssd1 vssd1 vccd1 vccd1 _21716_/A sky130_fd_sc_hd__nand3_4
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17966_ _17983_/A vssd1 vssd1 vccd1 vccd1 _17966_/X sky130_fd_sc_hd__clkbuf_2
X_13089_ _13089_/A vssd1 vssd1 vccd1 vccd1 _13090_/S sky130_fd_sc_hd__buf_4
XFILLER_214_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16917_ _16917_/A vssd1 vssd1 vccd1 vccd1 _16917_/Y sky130_fd_sc_hd__inv_2
X_19705_ _19705_/A vssd1 vssd1 vccd1 vccd1 _23494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17897_ _17908_/A _18021_/B vssd1 vssd1 vccd1 vccd1 _17983_/A sky130_fd_sc_hd__or2_1
XFILLER_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16848_ _16915_/S vssd1 vssd1 vccd1 vccd1 _16861_/S sky130_fd_sc_hd__buf_4
X_19636_ _19175_/X _23464_/Q _19638_/S vssd1 vssd1 vccd1 vccd1 _19637_/A sky130_fd_sc_hd__mux2_1
XFILLER_254_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19567_ _19567_/A vssd1 vssd1 vccd1 vccd1 _23433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16779_ _16779_/A vssd1 vssd1 vccd1 vccd1 _16795_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18518_ _23002_/Q _18518_/B vssd1 vssd1 vccd1 vccd1 _18518_/Y sky130_fd_sc_hd__nand2_1
XFILLER_222_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19498_ _19498_/A vssd1 vssd1 vccd1 vccd1 _23402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18449_ _16945_/A _18449_/B vssd1 vssd1 vccd1 vccd1 _18520_/A sky130_fd_sc_hd__nand2b_4
XFILLER_179_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_309_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21460_ _21460_/A _21459_/Y vssd1 vssd1 vccd1 vccd1 _21462_/A sky130_fd_sc_hd__or2b_1
XFILLER_239_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_348_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20411_ _23685_/Q _20482_/B vssd1 vssd1 vccd1 vccd1 _20411_/X sky130_fd_sc_hd__or2_1
XFILLER_336_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21391_ _21391_/A _21391_/B vssd1 vssd1 vccd1 vccd1 _21393_/A sky130_fd_sc_hd__nor2_1
XFILLER_308_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23130_ _23420_/CLK _23130_/D vssd1 vssd1 vccd1 vccd1 _23130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20342_ _20227_/X _20340_/X _20320_/A vssd1 vssd1 vccd1 vccd1 _20342_/X sky130_fd_sc_hd__o21a_1
XFILLER_135_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23061_ _23414_/CLK _23061_/D vssd1 vssd1 vccd1 vccd1 _23061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20273_ _21716_/A _20387_/B vssd1 vssd1 vccd1 vccd1 _20275_/B sky130_fd_sc_hd__or2_1
XFILLER_134_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_289_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22012_ _22012_/A _22012_/B vssd1 vssd1 vccd1 vccd1 _22013_/A sky130_fd_sc_hd__or2_1
XFILLER_310_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput207 localMemory_wb_adr_i[3] vssd1 vssd1 vccd1 vccd1 input207/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput218 localMemory_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input218/X sky130_fd_sc_hd__buf_6
XTAP_5429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput229 localMemory_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 input229/X sky130_fd_sc_hd__buf_6
XFILLER_25_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22914_ _23599_/CLK _22914_/D vssd1 vssd1 vccd1 vccd1 _22914_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_272_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23894_ _23895_/CLK _23894_/D vssd1 vssd1 vccd1 vccd1 _23894_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_327_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22845_ _23005_/CLK _22845_/D vssd1 vssd1 vccd1 vccd1 _22845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_260_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22776_ _23588_/CLK _22776_/D vssd1 vssd1 vccd1 vccd1 _22776_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21727_ _21801_/B _21727_/B vssd1 vssd1 vccd1 vccd1 _21727_/Y sky130_fd_sc_hd__xnor2_2
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_318_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21658_ _21658_/A _21658_/B vssd1 vssd1 vccd1 vccd1 _21658_/Y sky130_fd_sc_hd__nand2_1
X_12460_ _12465_/A _12459_/X _11843_/A vssd1 vssd1 vccd1 vccd1 _12460_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_339_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11411_ _11411_/A vssd1 vssd1 vccd1 vccd1 _12457_/S sky130_fd_sc_hd__buf_2
XFILLER_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20609_ _23723_/Q _20593_/X _20608_/X _20602_/X vssd1 vssd1 vccd1 vccd1 _23723_/D
+ sky130_fd_sc_hd__o211a_1
X_12391_ _12594_/A _12391_/B _12391_/C vssd1 vssd1 vccd1 vccd1 _21386_/A sky130_fd_sc_hd__and3_4
X_21589_ _21630_/A _21587_/Y _21973_/S vssd1 vssd1 vccd1 vccd1 _21589_/X sky130_fd_sc_hd__mux2_4
XFILLER_342_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11342_ _22485_/Q _22645_/Q _22324_/Q _23460_/Q _11364_/A _11365_/A vssd1 vssd1 vccd1
+ vccd1 _11343_/B sky130_fd_sc_hd__mux4_1
X_14130_ _14415_/S vssd1 vssd1 vccd1 vccd1 _14433_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_299_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23328_ _23424_/CLK _23328_/D vssd1 vssd1 vccd1 vccd1 _23328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_299_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_30_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23577_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_341_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14061_ _14064_/A _14066_/B _14061_/C vssd1 vssd1 vccd1 vccd1 _14061_/X sky130_fd_sc_hd__or3_1
X_11273_ _11273_/A vssd1 vssd1 vccd1 vccd1 _11683_/A sky130_fd_sc_hd__buf_4
X_23259_ _23549_/CLK _23259_/D vssd1 vssd1 vccd1 vccd1 _23259_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_7321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13012_ _13026_/A _14307_/B vssd1 vssd1 vccd1 vccd1 _13013_/A sky130_fd_sc_hd__nand2_1
XTAP_7354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17820_ _22783_/Q _17566_/X _17826_/S vssd1 vssd1 vccd1 vccd1 _17821_/A sky130_fd_sc_hd__mux2_1
XTAP_6653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17751_ _17751_/A vssd1 vssd1 vccd1 vccd1 _22752_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_14963_ _22515_/Q _14231_/A _14246_/B _14962_/X vssd1 vssd1 vccd1 vccd1 _14964_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16702_ _16702_/A vssd1 vssd1 vccd1 vccd1 _22489_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13914_ _21293_/A vssd1 vssd1 vccd1 vccd1 _13951_/A sky130_fd_sc_hd__clkbuf_2
X_17682_ _22722_/Q _17575_/X _17682_/S vssd1 vssd1 vccd1 vccd1 _17683_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14894_ _14893_/X _22264_/Q _14985_/S vssd1 vssd1 vccd1 vccd1 _14895_/A sky130_fd_sc_hd__mux2_1
XFILLER_331_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19421_ _19421_/A vssd1 vssd1 vccd1 vccd1 _23368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16633_ _16633_/A vssd1 vssd1 vccd1 vccd1 _22464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13845_ _13861_/A _14059_/C vssd1 vssd1 vccd1 vccd1 _13845_/Y sky130_fd_sc_hd__nor2_1
XINSDIODE2_304 _15990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_315 _16068_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_326 _16107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_337 _17100_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19352_ _19409_/S vssd1 vssd1 vccd1 vccd1 _19361_/S sky130_fd_sc_hd__buf_4
X_16564_ _15422_/X _22434_/Q _16568_/S vssd1 vssd1 vccd1 vccd1 _16565_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_348 _21975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13776_ _13776_/A _14207_/A vssd1 vssd1 vccd1 vccd1 _13777_/A sky130_fd_sc_hd__or2_4
XFILLER_62_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_359 _23791_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18303_ _18305_/A _18305_/C _18302_/Y vssd1 vssd1 vccd1 vccd1 _22927_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_349_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15515_ _14690_/A _15498_/X _17134_/A _15436_/X vssd1 vssd1 vccd1 vccd1 _15515_/X
+ sky130_fd_sc_hd__o22a_1
X_12727_ _12733_/A vssd1 vssd1 vccd1 vccd1 _12727_/X sky130_fd_sc_hd__buf_4
X_19283_ _19185_/X _23307_/Q _19289_/S vssd1 vssd1 vccd1 vccd1 _19284_/A sky130_fd_sc_hd__mux2_1
X_16495_ _16495_/A vssd1 vssd1 vccd1 vccd1 _22404_/D sky130_fd_sc_hd__clkbuf_1
X_18234_ _22905_/Q _18240_/B vssd1 vssd1 vccd1 vccd1 _18234_/X sky130_fd_sc_hd__or2_1
XFILLER_337_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15446_ _23762_/Q _15215_/A _15216_/A _15444_/X _15445_/X vssd1 vssd1 vccd1 vccd1
+ _15446_/X sky130_fd_sc_hd__a221o_1
X_12658_ _12683_/A _12658_/B vssd1 vssd1 vccd1 vccd1 _12658_/Y sky130_fd_sc_hd__nor2_1
XFILLER_175_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18165_ _18144_/B _18162_/X _18164_/Y vssd1 vssd1 vccd1 vccd1 _18165_/X sky130_fd_sc_hd__o21a_1
X_11609_ _11609_/A vssd1 vssd1 vccd1 vccd1 _12292_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15377_ _21708_/A vssd1 vssd1 vccd1 vccd1 _15377_/X sky130_fd_sc_hd__buf_12
XFILLER_306_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12589_ _22781_/Q _22749_/Q _22650_/Q _22717_/Q _12324_/X _12329_/X vssd1 vssd1 vccd1
+ vccd1 _12590_/B sky130_fd_sc_hd__mux4_1
XFILLER_239_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17116_ _15081_/A _17115_/X _17116_/S vssd1 vssd1 vccd1 vccd1 _17116_/X sky130_fd_sc_hd__mux2_1
X_14328_ _14326_/X _14327_/X _14331_/S vssd1 vssd1 vccd1 vccd1 _14328_/X sky130_fd_sc_hd__mux2_1
X_18096_ _18096_/A vssd1 vssd1 vccd1 vccd1 _18096_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_209_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17047_ _17047_/A vssd1 vssd1 vccd1 vccd1 _17078_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_292_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14259_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14259_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_292_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_289_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_332_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_314_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18998_ _18998_/A vssd1 vssd1 vccd1 vccd1 _23195_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_286_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_19 _17559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17949_ _22827_/Q _17932_/X _17945_/X _17948_/X vssd1 vssd1 vccd1 vccd1 _22827_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_273_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_300_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20960_ _21999_/A _20950_/X _20716_/B _20954_/X vssd1 vssd1 vccd1 vccd1 _20960_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19619_ _23457_/Q _19255_/A _19621_/S vssd1 vssd1 vccd1 vccd1 _19620_/A sky130_fd_sc_hd__mux2_1
XFILLER_226_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20891_ _20891_/A _20895_/B vssd1 vssd1 vccd1 vccd1 _20969_/A sky130_fd_sc_hd__or2_4
XFILLER_246_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22630_ _23575_/CLK _22630_/D vssd1 vssd1 vccd1 vccd1 _22630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22561_ _22977_/CLK _22561_/D vssd1 vssd1 vccd1 vccd1 _22561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21512_ _21472_/A _21468_/Y _21472_/C _21501_/B _21470_/B vssd1 vssd1 vccd1 vccd1
+ _21513_/B sky130_fd_sc_hd__o311a_1
XFILLER_22_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22492_ _23876_/CLK _22492_/D vssd1 vssd1 vccd1 vccd1 _22492_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_356_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_355_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21443_ _21443_/A vssd1 vssd1 vccd1 vccd1 _21716_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_175_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_308_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21374_ _21418_/A _21374_/B vssd1 vssd1 vccd1 vccd1 _21374_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_324_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_323_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_308_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23113_ _23561_/CLK _23113_/D vssd1 vssd1 vccd1 vccd1 _23113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20325_ _23672_/Q _20177_/A _20323_/Y _20324_/X vssd1 vssd1 vccd1 vccd1 _23672_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23044_ _23556_/CLK _23044_/D vssd1 vssd1 vccd1 vccd1 _23044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20256_ _17103_/A _20295_/A _20255_/Y vssd1 vssd1 vccd1 vccd1 _20256_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_304_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_304_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20187_ _20220_/A vssd1 vssd1 vccd1 vccd1 _20187_/X sky130_fd_sc_hd__buf_2
XTAP_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ _12047_/A _11960_/B vssd1 vssd1 vccd1 vccd1 _11960_/Y sky130_fd_sc_hd__nor2_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23946_ _23946_/CLK _23946_/D vssd1 vssd1 vccd1 vccd1 _23946_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_229_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23877_ _23877_/CLK _23877_/D vssd1 vssd1 vccd1 vccd1 _23877_/Q sky130_fd_sc_hd__dfxtp_1
X_11891_ _22365_/Q _22397_/Q _22686_/Q _23053_/Q _11777_/S _11590_/A vssd1 vssd1 vccd1
+ vccd1 _11891_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13630_ _23929_/Q _13588_/A _13629_/Y _13594_/A vssd1 vssd1 vccd1 vccd1 _13967_/A
+ sky130_fd_sc_hd__a22o_4
X_22828_ _22830_/CLK _22828_/D vssd1 vssd1 vccd1 vccd1 _22828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13561_ _13561_/A _13561_/B vssd1 vssd1 vccd1 vccd1 _13562_/B sky130_fd_sc_hd__xor2_4
X_22759_ _23578_/CLK _22759_/D vssd1 vssd1 vccd1 vccd1 _22759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15300_ _23599_/Q vssd1 vssd1 vccd1 vccd1 _19977_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_346_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12512_ _23205_/Q _23173_/Q _23141_/Q _23109_/Q _12501_/X _12502_/X vssd1 vssd1 vccd1
+ vccd1 _12512_/X sky130_fd_sc_hd__mux4_1
XFILLER_319_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16280_ _16280_/A vssd1 vssd1 vccd1 vccd1 _22315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13492_ _13492_/A _13492_/B _13632_/A _13492_/D vssd1 vssd1 vccd1 vccd1 _13492_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_8_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15231_ _15345_/A _15204_/X _15230_/X _15815_/A vssd1 vssd1 vccd1 vccd1 _15231_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_12443_ _12443_/A vssd1 vssd1 vccd1 vccd1 _14294_/A sky130_fd_sc_hd__buf_2
XFILLER_139_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_327_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15162_ _15162_/A vssd1 vssd1 vccd1 vccd1 _15162_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_354_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12374_ _12378_/A _12374_/B vssd1 vssd1 vccd1 vccd1 _12374_/X sky130_fd_sc_hd__or2_1
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14113_ _22887_/Q vssd1 vssd1 vccd1 vccd1 _14119_/C sky130_fd_sc_hd__clkbuf_2
X_11325_ _22388_/Q _22420_/Q _22709_/Q _23076_/Q _11468_/A _11469_/A vssd1 vssd1 vccd1
+ vccd1 _11326_/B sky130_fd_sc_hd__mux4_1
XFILLER_114_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19970_ _20008_/A _19970_/B _19985_/C vssd1 vssd1 vccd1 vccd1 _23604_/D sky130_fd_sc_hd__nor3_1
XFILLER_299_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15093_ _12287_/A _16054_/B _14674_/A _13920_/A _14836_/A vssd1 vssd1 vccd1 vccd1
+ _15093_/X sky130_fd_sc_hd__a221o_1
XFILLER_126_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_342_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18921_ _23161_/Q _18836_/X _18929_/S vssd1 vssd1 vccd1 vccd1 _18922_/A sky130_fd_sc_hd__mux2_1
X_14044_ input223/X _14038_/X _14043_/X vssd1 vssd1 vccd1 vccd1 _14044_/X sky130_fd_sc_hd__a21bo_4
X_11256_ _11763_/B vssd1 vssd1 vccd1 vccd1 _12801_/A sky130_fd_sc_hd__buf_6
XTAP_7140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_326_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18852_ _18852_/A vssd1 vssd1 vccd1 vccd1 _18852_/X sky130_fd_sc_hd__clkbuf_2
X_11187_ _22388_/Q _22420_/Q _22709_/Q _23076_/Q _13434_/A _11170_/X vssd1 vssd1 vccd1
+ vccd1 _11188_/B sky130_fd_sc_hd__mux4_1
XFILLER_95_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17803_ _17803_/A vssd1 vssd1 vccd1 vccd1 _22776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18783_ _23112_/Q _18782_/X _18786_/S vssd1 vssd1 vccd1 vccd1 _18784_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15995_ _15995_/A _15995_/B vssd1 vssd1 vccd1 vccd1 _15995_/Y sky130_fd_sc_hd__nand2_1
XTAP_5771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17734_ _17802_/S vssd1 vssd1 vccd1 vccd1 _17743_/S sky130_fd_sc_hd__buf_6
XTAP_5793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14946_ _15339_/S vssd1 vssd1 vccd1 vccd1 _15456_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_208_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17665_ _22714_/Q _17550_/X _17671_/S vssd1 vssd1 vccd1 vccd1 _17666_/A sky130_fd_sc_hd__mux2_1
X_14877_ _22949_/Q _14876_/X _15360_/A vssd1 vssd1 vccd1 vccd1 _14877_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_101 _21648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_112 _21773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19404_ _19404_/A vssd1 vssd1 vccd1 vccd1 _23361_/D sky130_fd_sc_hd__clkbuf_1
X_16616_ _22457_/Q _16217_/X _16618_/S vssd1 vssd1 vccd1 vccd1 _16617_/A sky130_fd_sc_hd__mux2_1
X_13828_ _13828_/A vssd1 vssd1 vccd1 vccd1 _13828_/X sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_123 _21386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17596_ _22693_/Q _17594_/X _17608_/S vssd1 vssd1 vccd1 vccd1 _17597_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_134 _20347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_145 _20362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_156 _21079_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19335_ _19261_/X _23331_/Q _19337_/S vssd1 vssd1 vccd1 vccd1 _19336_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16547_ _16547_/A vssd1 vssd1 vccd1 vccd1 _22426_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_167 _13972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13759_ _13810_/B _13739_/X _13758_/X _13730_/X vssd1 vssd1 vccd1 vccd1 _14032_/C
+ sky130_fd_sc_hd__a22oi_4
XINSDIODE2_178 _13701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_338_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_189 _13991_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19266_ _19266_/A vssd1 vssd1 vccd1 vccd1 _23300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16478_ _15240_/X _22397_/Q _16480_/S vssd1 vssd1 vccd1 vccd1 _16479_/A sky130_fd_sc_hd__mux2_1
XFILLER_349_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18217_ _18243_/A vssd1 vssd1 vccd1 vccd1 _18227_/B sky130_fd_sc_hd__clkbuf_1
X_15429_ _21738_/A vssd1 vssd1 vccd1 vccd1 _21737_/A sky130_fd_sc_hd__buf_12
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19197_ _19197_/A vssd1 vssd1 vccd1 vccd1 _19197_/X sky130_fd_sc_hd__buf_2
X_18148_ _18148_/A vssd1 vssd1 vccd1 vccd1 _22885_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_306_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_356_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_333_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_345_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_333_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18079_ _22864_/Q _18067_/X _18068_/X _22997_/Q _18069_/X vssd1 vssd1 vccd1 vccd1
+ _18079_/X sky130_fd_sc_hd__a221o_1
XFILLER_172_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20110_ _23643_/Q _23640_/Q _20110_/C _20112_/D vssd1 vssd1 vccd1 vccd1 _20123_/C
+ sky130_fd_sc_hd__and4_1
X_21090_ _21075_/Y _21085_/Y _21301_/D _20058_/X vssd1 vssd1 vccd1 vccd1 _21091_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20041_ _20041_/A _20041_/B _20056_/C vssd1 vssd1 vccd1 vccd1 _23624_/D sky130_fd_sc_hd__nor3_1
XFILLER_320_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_302_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_298_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23800_ _23942_/CLK _23800_/D vssd1 vssd1 vccd1 vccd1 _23800_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_65_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21992_ _23835_/Q _23769_/Q vssd1 vssd1 vccd1 vccd1 _21993_/B sky130_fd_sc_hd__nor2_1
XFILLER_273_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23731_ _23861_/CLK _23731_/D vssd1 vssd1 vccd1 vccd1 _23731_/Q sky130_fd_sc_hd__dfxtp_1
X_20943_ _17163_/A _20936_/X _20678_/B _20940_/X vssd1 vssd1 vccd1 vccd1 _20943_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23662_ _23818_/CLK _23662_/D vssd1 vssd1 vccd1 vccd1 _23662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ _20874_/A vssd1 vssd1 vccd1 vccd1 _23775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22613_ _22968_/CLK _22613_/D vssd1 vssd1 vccd1 vccd1 _22613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23593_ _23600_/CLK _23593_/D vssd1 vssd1 vccd1 vccd1 _23593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22544_ _23576_/CLK _22544_/D vssd1 vssd1 vccd1 vccd1 _22544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_329_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22475_ _23578_/CLK _22475_/D vssd1 vssd1 vccd1 vccd1 _22475_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_194_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_355_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21426_ _21425_/A _21425_/B _21342_/A _21342_/B vssd1 vssd1 vccd1 vccd1 _21426_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21357_ _23814_/Q _23813_/Q _21357_/C vssd1 vssd1 vccd1 vccd1 _21456_/A sky130_fd_sc_hd__and3b_4
XFILLER_135_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11110_ _23899_/Q vssd1 vssd1 vccd1 vccd1 _11146_/A sky130_fd_sc_hd__buf_4
XFILLER_107_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20308_ _20302_/X _20304_/Y _20306_/X _21861_/A _20307_/X vssd1 vssd1 vccd1 vccd1
+ _20680_/A sky130_fd_sc_hd__a32o_4
X_12090_ _22274_/Q _23090_/Q _23506_/Q _22435_/Q _11637_/A _11755_/A vssd1 vssd1 vccd1
+ vccd1 _12091_/B sky130_fd_sc_hd__mux4_1
X_21288_ _20544_/A _21191_/B _13603_/X vssd1 vssd1 vccd1 vccd1 _21297_/B sky130_fd_sc_hd__a21oi_1
XFILLER_311_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23027_ _23507_/CLK _23027_/D vssd1 vssd1 vccd1 vccd1 _23027_/Q sky130_fd_sc_hd__dfxtp_1
X_20239_ _23661_/Q _20277_/B vssd1 vssd1 vccd1 vccd1 _20239_/X sky130_fd_sc_hd__or2_1
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_295_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14800_ _14800_/A vssd1 vssd1 vccd1 vccd1 _14801_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_292_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_291_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _15780_/A vssd1 vssd1 vccd1 vccd1 _15931_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12992_ _22283_/Q _23099_/Q _23515_/Q _22444_/Q _12727_/X _12728_/X vssd1 vssd1 vccd1
+ vccd1 _12993_/B sky130_fd_sc_hd__mux4_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14731_ _14731_/A vssd1 vssd1 vccd1 vccd1 _14901_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_291_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23929_ _23936_/CLK _23929_/D vssd1 vssd1 vccd1 vccd1 _23929_/Q sky130_fd_sc_hd__dfxtp_4
X_11943_ _13392_/A _11943_/B vssd1 vssd1 vccd1 vccd1 _11943_/Y sky130_fd_sc_hd__nor2_1
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17450_ _22636_/Q _16278_/X _17454_/S vssd1 vssd1 vccd1 vccd1 _17451_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _14660_/X _14661_/X _14665_/S vssd1 vssd1 vccd1 vccd1 _14662_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11874_ _23214_/Q _23182_/Q _23150_/Q _23118_/Q _11305_/A _11869_/X vssd1 vssd1 vccd1
+ vccd1 _11875_/B sky130_fd_sc_hd__mux4_2
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16401_ _15104_/X _22363_/Q _16407_/S vssd1 vssd1 vccd1 vccd1 _16402_/A sky130_fd_sc_hd__mux2_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ _23927_/Q _13588_/A _13612_/X _13451_/A vssd1 vssd1 vccd1 vccd1 _13965_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_17381_ _17381_/A vssd1 vssd1 vccd1 vccd1 _22610_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14593_ _23590_/Q vssd1 vssd1 vccd1 vccd1 _19922_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_214_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19120_ _23249_/Q _18811_/X _19124_/S vssd1 vssd1 vccd1 vccd1 _19121_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16332_ _16332_/A vssd1 vssd1 vccd1 vccd1 _22333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13544_ _13188_/A _13543_/Y _15996_/A vssd1 vssd1 vccd1 vccd1 _13544_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_201_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_319_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19051_ _16860_/X _23219_/Q _19051_/S vssd1 vssd1 vccd1 vccd1 _19052_/A sky130_fd_sc_hd__mux2_1
X_16263_ _22310_/Q _16262_/X _16269_/S vssd1 vssd1 vccd1 vccd1 _16264_/A sky130_fd_sc_hd__mux2_1
XFILLER_335_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13475_ _13470_/X _13603_/A _13879_/A vssd1 vssd1 vccd1 vccd1 _13890_/A sky130_fd_sc_hd__a21oi_2
XFILLER_9_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18002_ input7/X input282/X _18005_/S vssd1 vssd1 vccd1 vccd1 _18002_/X sky130_fd_sc_hd__mux2_1
X_15214_ _23661_/Q _16021_/B vssd1 vssd1 vccd1 vccd1 _15214_/X sky130_fd_sc_hd__or2_1
XFILLER_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12426_ _22779_/Q _22747_/Q _22648_/Q _22715_/Q _12535_/S _11609_/A vssd1 vssd1 vccd1
+ vccd1 _12426_/X sky130_fd_sc_hd__mux4_1
X_16194_ _23009_/Q _16944_/A _16085_/X input239/X vssd1 vssd1 vccd1 vccd1 _16194_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_154_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15145_ _23756_/Q _14482_/X _14478_/X _15143_/X _15144_/X vssd1 vssd1 vccd1 vccd1
+ _15145_/X sky130_fd_sc_hd__a221o_1
Xoutput308 _13962_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[13] sky130_fd_sc_hd__buf_2
Xoutput319 _13980_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[24] sky130_fd_sc_hd__buf_2
X_12357_ _12241_/A _12354_/X _12356_/X vssd1 vssd1 vccd1 vccd1 _12357_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_337_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ _11308_/A vssd1 vssd1 vccd1 vccd1 _11532_/A sky130_fd_sc_hd__clkbuf_4
X_19953_ _23600_/Q _19977_/B _19953_/C vssd1 vssd1 vccd1 vccd1 _19959_/C sky130_fd_sc_hd__and3_1
XFILLER_287_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15076_ _22920_/Q _14868_/B _15075_/X _14727_/X vssd1 vssd1 vccd1 vccd1 _15076_/X
+ sky130_fd_sc_hd__a211o_1
X_12288_ _13510_/B vssd1 vssd1 vccd1 vccd1 _13920_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_142_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18904_ _18904_/A vssd1 vssd1 vccd1 vccd1 _23153_/D sky130_fd_sc_hd__clkbuf_1
X_14027_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14027_/X sky130_fd_sc_hd__buf_2
XFILLER_141_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11239_ _11424_/A _11239_/B vssd1 vssd1 vccd1 vccd1 _11239_/Y sky130_fd_sc_hd__nor2_1
X_19884_ _19884_/A vssd1 vssd1 vccd1 vccd1 _23574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18835_ _18835_/A vssd1 vssd1 vccd1 vccd1 _23128_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15978_ _15978_/A vssd1 vssd1 vccd1 vccd1 _22286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18766_ _18766_/A vssd1 vssd1 vccd1 vccd1 _23107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14929_ _22950_/Q _14926_/X _15885_/A vssd1 vssd1 vccd1 vccd1 _14929_/X sky130_fd_sc_hd__mux2_1
X_17717_ _17717_/A vssd1 vssd1 vccd1 vccd1 _17726_/S sky130_fd_sc_hd__buf_6
XFILLER_222_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18697_ _19699_/A _19843_/B vssd1 vssd1 vccd1 vccd1 _18754_/A sky130_fd_sc_hd__or2_4
XFILLER_282_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17648_ _17648_/A _17648_/B _17648_/C vssd1 vssd1 vccd1 vccd1 _17655_/B sky130_fd_sc_hd__and3_1
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17579_ _17646_/S vssd1 vssd1 vccd1 vccd1 _17592_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_338_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19318_ _19236_/X _23323_/Q _19322_/S vssd1 vssd1 vccd1 vccd1 _19319_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20590_ _17033_/A _20572_/X _20589_/Y vssd1 vssd1 vccd1 vccd1 _20591_/C sky130_fd_sc_hd__a21oi_2
XFILLER_176_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_338_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19249_ _19249_/A vssd1 vssd1 vccd1 vccd1 _19249_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22260_ _22260_/A _22260_/B vssd1 vssd1 vccd1 vccd1 _23946_/D sky130_fd_sc_hd__nor2_1
XFILLER_118_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21211_ _13440_/C _14970_/X _21214_/S vssd1 vssd1 vccd1 vccd1 _21212_/B sky130_fd_sc_hd__mux2_8
XFILLER_352_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_158_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23704_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22191_ _21838_/A _22189_/X _22190_/Y _21361_/A vssd1 vssd1 vccd1 vccd1 _22191_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_105_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21142_ _21142_/A vssd1 vssd1 vccd1 vccd1 _21142_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_321_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21073_ _21163_/A vssd1 vssd1 vccd1 vccd1 _21073_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_321_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20024_ _20034_/B _20034_/C vssd1 vssd1 vccd1 vccd1 _20025_/C sky130_fd_sc_hd__and2_1
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21975_ _21975_/A _21979_/A vssd1 vssd1 vccd1 vccd1 _21977_/A sky130_fd_sc_hd__nand2_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23714_ _23714_/CLK _23714_/D vssd1 vssd1 vccd1 vccd1 _23714_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20926_ _20926_/A vssd1 vssd1 vccd1 vccd1 _20926_/X sky130_fd_sc_hd__clkbuf_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23645_ _23646_/CLK _23645_/D vssd1 vssd1 vccd1 vccd1 _23645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20857_ _20716_/B _20846_/X _20847_/X _23771_/Q vssd1 vssd1 vccd1 vccd1 _20858_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_357_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23576_ _23576_/CLK _23576_/D vssd1 vssd1 vccd1 vccd1 _23576_/Q sky130_fd_sc_hd__dfxtp_1
X_11590_ _11590_/A vssd1 vssd1 vccd1 vccd1 _12073_/A sky130_fd_sc_hd__buf_4
XFILLER_356_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20788_ _20948_/A vssd1 vssd1 vccd1 vccd1 _20788_/X sky130_fd_sc_hd__buf_2
XFILLER_357_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_317_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22527_ _23467_/CLK _22527_/D vssd1 vssd1 vccd1 vccd1 _22527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_344_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13260_ _22385_/Q _22417_/Q _22706_/Q _23073_/Q _11206_/X _11208_/X vssd1 vssd1 vccd1
+ vccd1 _13260_/X sky130_fd_sc_hd__mux4_2
XFILLER_108_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_309_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22458_ _22618_/CLK _22458_/D vssd1 vssd1 vccd1 vccd1 _22458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_339_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_325_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_308_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12211_ _23468_/Q _23564_/Q _22528_/Q _22332_/Q _12209_/X _12210_/X vssd1 vssd1 vccd1
+ vccd1 _12211_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21409_ _21398_/X _21404_/Y _21406_/Y _21408_/X vssd1 vssd1 vccd1 vccd1 _21409_/X
+ sky130_fd_sc_hd__a211o_1
X_13191_ _22478_/Q _22638_/Q _13191_/S vssd1 vssd1 vccd1 vccd1 _13191_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22389_ _23902_/CLK _22389_/D vssd1 vssd1 vccd1 vccd1 _22389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_340_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_312_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12142_ _23313_/Q _23281_/Q _23249_/Q _23537_/Q _11457_/C _12020_/A vssd1 vssd1 vccd1
+ vccd1 _12142_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16950_ _17244_/C _16950_/B vssd1 vssd1 vccd1 vccd1 _16951_/A sky130_fd_sc_hd__and2_1
X_12073_ _12073_/A _12073_/B vssd1 vssd1 vccd1 vccd1 _12073_/Y sky130_fd_sc_hd__nand2_1
XFILLER_150_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15901_ _15901_/A _15901_/B vssd1 vssd1 vccd1 vccd1 _15942_/A sky130_fd_sc_hd__nor2_4
X_16881_ _16879_/X _22541_/Q _16893_/S vssd1 vssd1 vccd1 vccd1 _16882_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18620_ _18620_/A vssd1 vssd1 vccd1 vccd1 _23042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15832_ _15832_/A vssd1 vssd1 vccd1 vccd1 _15964_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_264_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18551_ _18551_/A vssd1 vssd1 vccd1 vccd1 _23012_/D sky130_fd_sc_hd__clkbuf_1
X_15763_ _15440_/X _15756_/X _15762_/X _14497_/A vssd1 vssd1 vccd1 vccd1 _15763_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _12968_/Y _12970_/Y _12972_/Y _12974_/Y _11246_/A vssd1 vssd1 vccd1 vccd1
+ _12988_/A sky130_fd_sc_hd__o221a_2
XFILLER_280_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_2_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_346_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ _17502_/A vssd1 vssd1 vccd1 vccd1 _22658_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14714_ _21339_/B _21339_/C vssd1 vssd1 vccd1 vccd1 _14714_/X sky130_fd_sc_hd__and2_1
X_18482_ _22988_/Q _18492_/B vssd1 vssd1 vccd1 vccd1 _18482_/Y sky130_fd_sc_hd__nand2_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ _11926_/A _11926_/B vssd1 vssd1 vccd1 vccd1 _11926_/X sky130_fd_sc_hd__or2_1
X_15694_ _16028_/A _15694_/B vssd1 vssd1 vccd1 vccd1 _15694_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _17433_/A vssd1 vssd1 vccd1 vccd1 _22628_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _14643_/X _14644_/X _14853_/S vssd1 vssd1 vccd1 vccd1 _14645_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _12260_/A _11857_/B _11857_/C vssd1 vssd1 vccd1 vccd1 _13745_/A sky130_fd_sc_hd__nor3_4
XFILLER_348_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_348_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17364_ _17364_/A vssd1 vssd1 vccd1 vccd1 _22602_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14576_ _14724_/A _14576_/B vssd1 vssd1 vccd1 vccd1 _15243_/A sky130_fd_sc_hd__nand2_1
XFILLER_158_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11788_ _22271_/Q _23087_/Q _23503_/Q _22432_/Q _11893_/S _11621_/X vssd1 vssd1 vccd1
+ vccd1 _11789_/B sky130_fd_sc_hd__mux4_1
XFILLER_198_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_348_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19103_ _19103_/A vssd1 vssd1 vccd1 vccd1 _23241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16315_ _16315_/A vssd1 vssd1 vccd1 vccd1 _22325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13527_ _13524_/Y _13526_/X _11940_/A vssd1 vssd1 vccd1 vccd1 _13528_/C sky130_fd_sc_hd__a21oi_1
X_17295_ _22581_/Q _17255_/X _17240_/X _17294_/X vssd1 vssd1 vccd1 vccd1 _22581_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_203_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_348_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_319_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19034_ _16835_/X _23211_/Q _19040_/S vssd1 vssd1 vccd1 vccd1 _19035_/A sky130_fd_sc_hd__mux2_1
X_16246_ _18811_/A vssd1 vssd1 vccd1 vccd1 _16246_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_348_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13458_ _23945_/Q vssd1 vssd1 vccd1 vccd1 _13570_/A sky130_fd_sc_hd__buf_2
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12409_ _22779_/Q _22747_/Q _22648_/Q _22715_/Q _11305_/A _11869_/X vssd1 vssd1 vccd1
+ vccd1 _12410_/B sky130_fd_sc_hd__mux4_1
X_16177_ _22977_/Q _16176_/X _16177_/S vssd1 vssd1 vccd1 vccd1 _16177_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13389_ _13329_/A _13322_/C _13388_/Y vssd1 vssd1 vccd1 vccd1 _13389_/X sky130_fd_sc_hd__a21o_1
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15128_ _15089_/S _15127_/Y _14860_/X vssd1 vssd1 vccd1 vccd1 _15915_/B sky130_fd_sc_hd__a21o_1
XFILLER_217_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_330_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19936_ _23594_/Q _23593_/Q _23590_/Q _23589_/Q vssd1 vssd1 vccd1 vccd1 _19938_/B
+ sky130_fd_sc_hd__and4_1
X_15059_ input156/X _13650_/A _14967_/S input121/X _14235_/A vssd1 vssd1 vccd1 vccd1
+ _15059_/X sky130_fd_sc_hd__a221o_4
XFILLER_330_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_330_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19867_ _19913_/S vssd1 vssd1 vccd1 vccd1 _19876_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_255_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18818_ _23123_/Q _18817_/X _18818_/S vssd1 vssd1 vccd1 vccd1 _18819_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19798_ _23536_/Q _19201_/A _19804_/S vssd1 vssd1 vccd1 vccd1 _19799_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18749_ _18749_/A vssd1 vssd1 vccd1 vccd1 _23099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21760_ _22215_/A _21760_/B vssd1 vssd1 vccd1 vccd1 _21760_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20711_ _20727_/A _20711_/B _20711_/C vssd1 vssd1 vccd1 vccd1 _20711_/X sky130_fd_sc_hd__or3_1
XFILLER_196_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21691_ _21548_/A _21548_/B _21690_/X vssd1 vssd1 vccd1 vccd1 _21696_/A sky130_fd_sc_hd__o21a_1
XFILLER_52_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23430_ _23558_/CLK _23430_/D vssd1 vssd1 vccd1 vccd1 _23430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_339_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20642_ _20642_/A vssd1 vssd1 vccd1 vccd1 _20642_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_338_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_354_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23361_ _23451_/CLK _23361_/D vssd1 vssd1 vccd1 vccd1 _23361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20573_ _20642_/A vssd1 vssd1 vccd1 vccd1 _20773_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_338_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_339_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22312_ _23580_/CLK _22312_/D vssd1 vssd1 vccd1 vccd1 _22312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23292_ _23545_/CLK _23292_/D vssd1 vssd1 vccd1 vccd1 _23292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_258_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22243_ _21361_/A _22241_/Y _22242_/X _21410_/A vssd1 vssd1 vccd1 vccd1 _22243_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_127_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_306_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22174_ _21491_/X _22154_/X _22173_/X vssd1 vssd1 vccd1 vccd1 _22174_/X sky130_fd_sc_hd__a21bo_1
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21125_ _23857_/Q _21123_/X _21124_/X _20631_/A vssd1 vssd1 vccd1 vccd1 _21126_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_322_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_321_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_294_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21056_ _23837_/Q _21068_/B vssd1 vssd1 vccd1 vccd1 _21056_/X sky130_fd_sc_hd__or2_1
XFILLER_293_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20007_ _20009_/A _23611_/Q _20007_/C _20014_/D vssd1 vssd1 vccd1 vccd1 _20021_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_247_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_55_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _22695_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_235_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12760_ _12825_/A vssd1 vssd1 vccd1 vccd1 _12922_/S sky130_fd_sc_hd__buf_6
XFILLER_43_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21958_ _21949_/A _21714_/A _21942_/Y _21957_/X _18135_/X vssd1 vssd1 vccd1 vccd1
+ _23931_/D sky130_fd_sc_hd__o221a_1
XFILLER_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11711_ _12071_/A _11708_/X _11710_/X vssd1 vssd1 vccd1 vccd1 _11711_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_199_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20909_ _21431_/A _20908_/X _20591_/B _20897_/X vssd1 vssd1 vccd1 vccd1 _20909_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12836_/A _12691_/B vssd1 vssd1 vccd1 vccd1 _12691_/Y sky130_fd_sc_hd__nor2_1
XFILLER_215_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21889_ _21889_/A _21889_/B vssd1 vssd1 vccd1 vccd1 _21892_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14897_/A vssd1 vssd1 vccd1 vccd1 _14431_/A sky130_fd_sc_hd__buf_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23628_ _23632_/CLK _23628_/D vssd1 vssd1 vccd1 vccd1 _23628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_329_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11642_ _12028_/A vssd1 vssd1 vccd1 vccd1 _12842_/A sky130_fd_sc_hd__buf_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14361_ _14952_/S vssd1 vssd1 vccd1 vccd1 _14949_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23559_ _23559_/CLK _23559_/D vssd1 vssd1 vccd1 vccd1 _23559_/Q sky130_fd_sc_hd__dfxtp_1
X_11573_ _11719_/A vssd1 vssd1 vccd1 vccd1 _11574_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_356_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16100_ _22975_/Q _16144_/S vssd1 vssd1 vccd1 vccd1 _16100_/X sky130_fd_sc_hd__or2_1
Xinput18 core_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_317_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13312_ _13314_/A _13311_/X _11489_/Y _13427_/A vssd1 vssd1 vccd1 vccd1 _13312_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_329_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17080_ _17070_/X _17071_/X _17079_/X _17057_/X vssd1 vssd1 vccd1 vccd1 _17080_/X
+ sky130_fd_sc_hd__o211a_4
Xinput29 core_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14292_ _14292_/A vssd1 vssd1 vccd1 vccd1 _14635_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16031_ _13406_/Y _13562_/B _16031_/S vssd1 vssd1 vccd1 vccd1 _16031_/X sky130_fd_sc_hd__mux2_1
X_13243_ _13188_/A _13543_/A _13242_/X vssd1 vssd1 vccd1 vccd1 _13243_/X sky130_fd_sc_hd__o21a_1
XFILLER_182_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13174_ _11288_/A _13167_/X _13169_/X _13173_/X _11379_/A vssd1 vssd1 vccd1 vccd1
+ _13184_/B sky130_fd_sc_hd__a311o_1
XFILLER_312_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12125_ _23313_/Q _23281_/Q _23249_/Q _23537_/Q _11561_/A _11613_/X vssd1 vssd1 vccd1
+ vccd1 _12126_/B sky130_fd_sc_hd__mux4_1
XFILLER_233_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17982_ input2/X input268/X _17987_/S vssd1 vssd1 vccd1 vccd1 _17982_/X sky130_fd_sc_hd__mux2_1
XFILLER_269_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_312_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19721_ _19194_/X _23502_/Q _19721_/S vssd1 vssd1 vccd1 vccd1 _19722_/A sky130_fd_sc_hd__mux2_1
XFILLER_334_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_313_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12056_ _12056_/A _12056_/B vssd1 vssd1 vccd1 vccd1 _12056_/Y sky130_fd_sc_hd__nor2_1
X_16933_ _22908_/Q _14160_/X _16929_/A _22601_/Q _14553_/C vssd1 vssd1 vccd1 vccd1
+ _22249_/C sky130_fd_sc_hd__a221oi_4
XFILLER_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19652_ _19197_/X _23471_/Q _19660_/S vssd1 vssd1 vccd1 vccd1 _19653_/A sky130_fd_sc_hd__mux2_1
X_16864_ _16896_/A vssd1 vssd1 vccd1 vccd1 _16877_/S sky130_fd_sc_hd__buf_4
XFILLER_93_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18603_ _18603_/A vssd1 vssd1 vccd1 vccd1 _23034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_280_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15815_ _15815_/A _15815_/B vssd1 vssd1 vccd1 vccd1 _15815_/Y sky130_fd_sc_hd__nand2_1
X_19583_ _19583_/A vssd1 vssd1 vccd1 vccd1 _23440_/D sky130_fd_sc_hd__clkbuf_1
X_16795_ _16795_/A _16795_/B vssd1 vssd1 vccd1 vccd1 _16796_/A sky130_fd_sc_hd__or2_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_350_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18534_ _23009_/Q _18534_/B vssd1 vssd1 vccd1 vccd1 _18534_/Y sky130_fd_sc_hd__nand2_1
X_15746_ _15746_/A vssd1 vssd1 vccd1 vccd1 _16047_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_92_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12958_ _12958_/A _12958_/B vssd1 vssd1 vccd1 vccd1 _12958_/X sky130_fd_sc_hd__or2_1
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11909_ _12134_/A _11909_/B _11909_/C vssd1 vssd1 vccd1 vccd1 _13778_/A sky130_fd_sc_hd__nor3_4
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18465_ _22982_/Q _18465_/B vssd1 vssd1 vccd1 vccd1 _18465_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15677_ _15674_/X _15675_/Y _15676_/X vssd1 vssd1 vccd1 vccd1 _15677_/Y sky130_fd_sc_hd__a21oi_1
X_12889_ _12882_/Y _12884_/Y _12886_/Y _12888_/Y _11559_/X vssd1 vssd1 vccd1 vccd1
+ _12889_/X sky130_fd_sc_hd__o221a_2
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14628_ _15339_/S _14627_/X _14767_/A vssd1 vssd1 vccd1 vccd1 _14629_/A sky130_fd_sc_hd__o21a_1
X_17416_ _17416_/A vssd1 vssd1 vccd1 vccd1 _22620_/D sky130_fd_sc_hd__clkbuf_1
X_18396_ _22959_/Q _18394_/B _18395_/Y vssd1 vssd1 vccd1 vccd1 _22959_/D sky130_fd_sc_hd__o21a_1
XFILLER_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17347_ _22595_/Q input212/X _17347_/S vssd1 vssd1 vccd1 vccd1 _17348_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14559_ _19699_/A _19627_/A vssd1 vssd1 vccd1 vccd1 _15976_/A sky130_fd_sc_hd__or2_4
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_336_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_308_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_308_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17278_ _23938_/Q vssd1 vssd1 vccd1 vccd1 _22139_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_307_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_323_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_307_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19017_ _19017_/A vssd1 vssd1 vccd1 vccd1 _23204_/D sky130_fd_sc_hd__clkbuf_1
X_16229_ _16229_/A vssd1 vssd1 vccd1 vccd1 _22299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_350_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_288_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19919_ _19915_/X _19916_/X _19922_/B vssd1 vssd1 vccd1 vccd1 _19919_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_229_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22930_ _22961_/CLK _22930_/D vssd1 vssd1 vccd1 vccd1 _22930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_290_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22861_ _23008_/CLK _22861_/D vssd1 vssd1 vccd1 vccd1 _22861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21812_ _21934_/A _21812_/B vssd1 vssd1 vccd1 vccd1 _21813_/C sky130_fd_sc_hd__and2b_1
XFILLER_25_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22792_ _23450_/CLK _22792_/D vssd1 vssd1 vccd1 vccd1 _22792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21743_ _21981_/A _21743_/B vssd1 vssd1 vccd1 vccd1 _21743_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21674_ _21674_/A _21674_/B vssd1 vssd1 vccd1 vccd1 _21675_/B sky130_fd_sc_hd__nor2_1
XFILLER_106_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23413_ _23541_/CLK _23413_/D vssd1 vssd1 vccd1 vccd1 _23413_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_173_wb_clk_i _23917_/CLK vssd1 vssd1 vccd1 vccd1 _23804_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_184_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20625_ _21601_/A _20572_/X _20624_/Y vssd1 vssd1 vccd1 vccd1 _20626_/C sky130_fd_sc_hd__a21oi_2
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_339_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_338_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_326_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_102_wb_clk_i _22899_/CLK vssd1 vssd1 vccd1 vccd1 _23264_/CLK sky130_fd_sc_hd__clkbuf_16
X_23344_ _23951_/A _23344_/D vssd1 vssd1 vccd1 vccd1 _23344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20556_ _20730_/A vssd1 vssd1 vccd1 vccd1 _20768_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_354_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_342_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_295_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_314_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23275_ _23467_/CLK _23275_/D vssd1 vssd1 vccd1 vccd1 _23275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_354_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_353_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20487_ _23714_/Q _20487_/B vssd1 vssd1 vccd1 vccd1 _20487_/X sky130_fd_sc_hd__or2_1
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_307_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_298_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_353_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_341_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_313_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22226_ _21379_/X _22208_/X _22215_/Y _22225_/X _21410_/X vssd1 vssd1 vccd1 vccd1
+ _22226_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_118_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_341_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22157_ _22053_/A _22155_/X _22156_/X vssd1 vssd1 vccd1 vccd1 _22176_/A sky130_fd_sc_hd__a21oi_4
XFILLER_310_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput480 _23938_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[27] sky130_fd_sc_hd__buf_2
XFILLER_133_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput491 _23919_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[8] sky130_fd_sc_hd__buf_2
XTAP_6857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21108_ _21108_/A _21108_/B vssd1 vssd1 vccd1 vccd1 _23851_/D sky130_fd_sc_hd__nor2_1
XTAP_6868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22088_ _22065_/A _22085_/Y _22086_/X _22087_/Y vssd1 vssd1 vccd1 vccd1 _22090_/A
+ sky130_fd_sc_hd__a211o_1
XTAP_6879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13930_ _21522_/A vssd1 vssd1 vccd1 vccd1 _13931_/B sky130_fd_sc_hd__buf_6
X_21039_ _23830_/Q _21048_/B vssd1 vssd1 vccd1 vccd1 _21039_/X sky130_fd_sc_hd__or2_1
X_13861_ _13861_/A _14064_/C vssd1 vssd1 vccd1 vccd1 _13861_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15600_ _23765_/Q _15595_/X _15596_/X _15598_/X _15599_/X vssd1 vssd1 vccd1 vccd1
+ _15600_/X sky130_fd_sc_hd__a221o_2
XFILLER_290_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12812_ _13629_/A _12812_/B vssd1 vssd1 vccd1 vccd1 _12812_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16580_ _16580_/A vssd1 vssd1 vccd1 vccd1 _22441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_508 _15656_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13792_ _11627_/B _13798_/B _13709_/A vssd1 vssd1 vccd1 vccd1 _13792_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_222_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_519 _22493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15531_ _15611_/B _15531_/B vssd1 vssd1 vccd1 vccd1 _15531_/X sky130_fd_sc_hd__or2_4
XFILLER_215_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _12741_/Y _12743_/B vssd1 vssd1 vccd1 vccd1 _13532_/C sky130_fd_sc_hd__and2b_1
XFILLER_349_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ hold5/X _18242_/X _18249_/X _18245_/X vssd1 vssd1 vccd1 vccd1 _22911_/D sky130_fd_sc_hd__o211a_1
XFILLER_188_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ _16034_/A _15458_/X _15459_/X _14621_/A _15461_/X vssd1 vssd1 vccd1 vccd1
+ _15462_/X sky130_fd_sc_hd__o221a_2
X_12674_ _22312_/Q _23448_/Q _12819_/S vssd1 vssd1 vccd1 vccd1 _12674_/X sky130_fd_sc_hd__mux2_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _21950_/A vssd1 vssd1 vccd1 vccd1 _21949_/A sky130_fd_sc_hd__clkbuf_16
X_14413_ _14178_/A _14552_/C _14415_/S vssd1 vssd1 vccd1 vccd1 _14458_/B sky130_fd_sc_hd__mux2_1
XFILLER_203_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18181_ _18181_/A vssd1 vssd1 vccd1 vccd1 _18195_/A sky130_fd_sc_hd__clkbuf_2
X_11625_ _12700_/A _11615_/X _11619_/X _11624_/X _11217_/A vssd1 vssd1 vccd1 vccd1
+ _11625_/X sky130_fd_sc_hd__a311o_2
X_15393_ _14621_/A _15384_/X _15390_/X _15392_/X vssd1 vssd1 vccd1 vccd1 _15393_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_318_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_329_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_317_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17132_ input83/X input48/X _17132_/S vssd1 vssd1 vccd1 vccd1 _17132_/X sky130_fd_sc_hd__mux2_8
XFILLER_345_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14344_ _14369_/A vssd1 vssd1 vccd1 vccd1 _14660_/S sky130_fd_sc_hd__clkbuf_4
X_11556_ _11557_/A _11557_/B vssd1 vssd1 vccd1 vccd1 _11558_/A sky130_fd_sc_hd__nor2_1
XFILLER_344_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17063_ _23468_/Q _17061_/X _17062_/X _17042_/X _15155_/X vssd1 vssd1 vccd1 vccd1
+ _17063_/X sky130_fd_sc_hd__a32o_1
X_14275_ _14343_/S _13514_/B _14274_/Y vssd1 vssd1 vccd1 vccd1 _14275_/X sky130_fd_sc_hd__a21o_1
XFILLER_333_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11487_ _16005_/A _20394_/A _11486_/X vssd1 vssd1 vccd1 vccd1 _13306_/B sky130_fd_sc_hd__o21ai_4
XFILLER_137_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_344_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16014_ _16013_/X _22287_/Q _16125_/S vssd1 vssd1 vccd1 vccd1 _16015_/A sky130_fd_sc_hd__mux2_1
X_13226_ _23421_/Q _23037_/Q _23389_/Q _23357_/Q _11526_/A _11519_/A vssd1 vssd1 vccd1
+ vccd1 _13226_/X sky130_fd_sc_hd__mux4_2
XFILLER_298_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_350_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13157_ _22286_/Q _23102_/Q _23518_/Q _22447_/Q _13034_/S _13096_/X vssd1 vssd1 vccd1
+ vccd1 _13158_/B sky130_fd_sc_hd__mux4_1
XFILLER_301_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12108_ _12101_/X _12103_/X _12105_/X _12107_/X _11275_/A vssd1 vssd1 vccd1 vccd1
+ _12109_/C sky130_fd_sc_hd__a221o_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17965_ _17981_/A vssd1 vssd1 vccd1 vccd1 _17965_/X sky130_fd_sc_hd__clkbuf_2
X_13088_ _22319_/Q _23455_/Q _13088_/S vssd1 vssd1 vccd1 vccd1 _13088_/X sky130_fd_sc_hd__mux2_1
XFILLER_312_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_300_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19704_ _19169_/X _23494_/Q _19710_/S vssd1 vssd1 vccd1 vccd1 _19705_/A sky130_fd_sc_hd__mux2_1
X_12039_ _22791_/Q _22759_/Q _22660_/Q _22727_/Q _12675_/A _12746_/A vssd1 vssd1 vccd1
+ vccd1 _12040_/B sky130_fd_sc_hd__mux4_1
X_16916_ _16916_/A vssd1 vssd1 vccd1 vccd1 _22552_/D sky130_fd_sc_hd__clkbuf_1
X_17896_ _17986_/A vssd1 vssd1 vccd1 vccd1 _17896_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19635_ _19635_/A vssd1 vssd1 vccd1 vccd1 _23463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16847_ _19197_/A vssd1 vssd1 vccd1 vccd1 _16847_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19566_ _23433_/Q _19178_/A _19566_/S vssd1 vssd1 vccd1 vccd1 _19567_/A sky130_fd_sc_hd__mux2_1
X_16778_ _16778_/A vssd1 vssd1 vccd1 vccd1 _22510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18517_ _18507_/X _18515_/Y _18516_/X vssd1 vssd1 vccd1 vccd1 _23001_/D sky130_fd_sc_hd__a21oi_1
XFILLER_280_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15729_ _23736_/Q _23866_/Q _15729_/S vssd1 vssd1 vccd1 vccd1 _15729_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_0_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23530_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19497_ _19181_/X _23402_/Q _19505_/S vssd1 vssd1 vccd1 vccd1 _19498_/A sky130_fd_sc_hd__mux2_1
XFILLER_233_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18448_ _22977_/Q _18445_/B _18447_/Y vssd1 vssd1 vccd1 vccd1 _22977_/D sky130_fd_sc_hd__o21a_1
XFILLER_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18379_ _22953_/Q _18377_/B _18378_/Y vssd1 vssd1 vccd1 vccd1 _22953_/D sky130_fd_sc_hd__o21a_1
XFILLER_187_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20410_ _20470_/A vssd1 vssd1 vccd1 vccd1 _20482_/B sky130_fd_sc_hd__buf_4
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21390_ _21425_/A _21425_/B vssd1 vssd1 vccd1 vccd1 _21391_/B sky130_fd_sc_hd__and2_1
XFILLER_239_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20341_ _15846_/Y _20295_/X _20340_/X vssd1 vssd1 vccd1 vccd1 _20341_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_323_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_323_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23060_ _23572_/CLK _23060_/D vssd1 vssd1 vccd1 vccd1 _23060_/Q sky130_fd_sc_hd__dfxtp_1
X_20272_ _20333_/A vssd1 vssd1 vccd1 vccd1 _20272_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_332_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_288_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22011_ _21989_/A _21989_/B _22010_/Y vssd1 vssd1 vccd1 vccd1 _22017_/A sky130_fd_sc_hd__o21ai_1
XTAP_6109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_289_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_289_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput208 localMemory_wb_adr_i[4] vssd1 vssd1 vccd1 vccd1 input208/X sky130_fd_sc_hd__clkbuf_1
Xinput219 localMemory_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input219/X sky130_fd_sc_hd__buf_6
XFILLER_76_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22913_ _22956_/CLK _22913_/D vssd1 vssd1 vccd1 vccd1 _22913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23893_ _23893_/CLK _23893_/D vssd1 vssd1 vccd1 vccd1 _23893_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_272_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22844_ _22893_/CLK _22844_/D vssd1 vssd1 vccd1 vccd1 _22844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22775_ _23893_/CLK _22775_/D vssd1 vssd1 vccd1 vccd1 _22775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_347_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21726_ _21801_/A _21697_/B _21725_/X vssd1 vssd1 vccd1 vccd1 _21727_/B sky130_fd_sc_hd__a21o_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_303_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21657_ _21624_/A _21624_/B _21624_/C _21694_/A vssd1 vssd1 vccd1 vccd1 _21658_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_33_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_339_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11410_ _23899_/Q vssd1 vssd1 vccd1 vccd1 _11411_/A sky130_fd_sc_hd__buf_4
X_20608_ _20626_/A _20608_/B _20608_/C vssd1 vssd1 vccd1 vccd1 _20608_/X sky130_fd_sc_hd__or3_1
X_12390_ _12383_/X _12385_/X _12387_/X _12389_/X _11273_/A vssd1 vssd1 vccd1 vccd1
+ _12391_/C sky130_fd_sc_hd__a221o_1
X_21588_ _21816_/A vssd1 vssd1 vccd1 vccd1 _21973_/S sky130_fd_sc_hd__buf_6
XFILLER_32_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23327_ _23327_/CLK _23327_/D vssd1 vssd1 vccd1 vccd1 _23327_/Q sky130_fd_sc_hd__dfxtp_1
X_11341_ _22808_/Q _22776_/Q _22677_/Q _22744_/Q _11468_/A _11469_/A vssd1 vssd1 vccd1
+ vccd1 _11341_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20539_ _20759_/B vssd1 vssd1 vccd1 vccd1 _21301_/C sky130_fd_sc_hd__buf_4
XFILLER_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_314_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14060_ input232/X _14058_/X _14059_/X vssd1 vssd1 vccd1 vccd1 _14060_/X sky130_fd_sc_hd__a21bo_4
XTAP_7300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23258_ _23420_/CLK _23258_/D vssd1 vssd1 vccd1 vccd1 _23258_/Q sky130_fd_sc_hd__dfxtp_1
X_11272_ _11272_/A vssd1 vssd1 vccd1 vccd1 _11273_/A sky130_fd_sc_hd__clkbuf_8
XTAP_7311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13011_ _17224_/A _20340_/A _13500_/A vssd1 vssd1 vccd1 vccd1 _14307_/B sky130_fd_sc_hd__mux2_4
XTAP_7333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22209_ _23843_/Q _23777_/Q vssd1 vssd1 vccd1 vccd1 _22211_/A sky130_fd_sc_hd__and2_1
XTAP_7344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23189_ _23349_/CLK _23189_/D vssd1 vssd1 vccd1 vccd1 _23189_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_70_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23546_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14962_ input163/X input127/X _15114_/S vssd1 vssd1 vccd1 vccd1 _14962_/X sky130_fd_sc_hd__mux2_8
XTAP_5953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17750_ _22752_/Q _17569_/X _17754_/S vssd1 vssd1 vccd1 vccd1 _17751_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_94_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16701_ _16704_/A _16701_/B vssd1 vssd1 vccd1 vccd1 _16702_/A sky130_fd_sc_hd__or2_1
XFILLER_59_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13913_ _13913_/A _13913_/B vssd1 vssd1 vccd1 vccd1 _13913_/Y sky130_fd_sc_hd__xnor2_4
X_14893_ _19175_/A vssd1 vssd1 vccd1 vccd1 _14893_/X sky130_fd_sc_hd__clkbuf_2
X_17681_ _17681_/A vssd1 vssd1 vccd1 vccd1 _22721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19420_ _23368_/Q _18782_/X _19422_/S vssd1 vssd1 vccd1 vccd1 _19421_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13844_ _13840_/Y _13842_/Y _13843_/X vssd1 vssd1 vccd1 vccd1 _14059_/C sky130_fd_sc_hd__o21ai_4
X_16632_ _22464_/Q _16239_/X _16640_/S vssd1 vssd1 vccd1 vccd1 _16633_/A sky130_fd_sc_hd__mux2_1
XFILLER_262_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_305 _15990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_316 _17289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_327 _16107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19351_ _19351_/A vssd1 vssd1 vccd1 vccd1 _23337_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_338 _17110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16563_ _16563_/A vssd1 vssd1 vccd1 vccd1 _22433_/D sky130_fd_sc_hd__clkbuf_1
X_13775_ _13775_/A _13775_/B _20148_/A _13775_/D vssd1 vssd1 vccd1 vccd1 _13776_/A
+ sky130_fd_sc_hd__or4_2
XINSDIODE2_349 _21975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18302_ _18305_/A _18305_/C _18292_/X vssd1 vssd1 vccd1 vccd1 _18302_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_215_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12726_ _12949_/A vssd1 vssd1 vccd1 vccd1 _12993_/A sky130_fd_sc_hd__buf_2
X_15514_ _14755_/A _15500_/X _15513_/X vssd1 vssd1 vccd1 vccd1 _17134_/A sky130_fd_sc_hd__o21ai_4
XFILLER_204_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16494_ _15570_/X _22404_/Q _16502_/S vssd1 vssd1 vccd1 vccd1 _16495_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19282_ _19282_/A vssd1 vssd1 vccd1 vccd1 _23306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18233_ hold4/X _18229_/X _18231_/X _18232_/X vssd1 vssd1 vccd1 vccd1 _22904_/D sky130_fd_sc_hd__o211a_1
XFILLER_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15445_ _23794_/Q _15219_/A _14919_/A vssd1 vssd1 vccd1 vccd1 _15445_/X sky130_fd_sc_hd__a21o_1
X_12657_ _22277_/Q _23093_/Q _23509_/Q _22438_/Q _12751_/S _12685_/A vssd1 vssd1 vccd1
+ vccd1 _12658_/B sky130_fd_sc_hd__mux4_2
XFILLER_129_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11608_ _11893_/S vssd1 vssd1 vccd1 vccd1 _12043_/S sky130_fd_sc_hd__buf_4
XFILLER_175_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18164_ _18164_/A _18164_/B vssd1 vssd1 vccd1 vccd1 _18164_/Y sky130_fd_sc_hd__nor2_1
XFILLER_191_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15376_ _21708_/A _21673_/A _15376_/C vssd1 vssd1 vccd1 vccd1 _15430_/B sky130_fd_sc_hd__and3_2
XFILLER_318_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12588_ _12590_/A _12587_/X _11282_/A vssd1 vssd1 vccd1 vccd1 _12588_/X sky130_fd_sc_hd__o21a_1
XFILLER_345_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17115_ _23473_/Q _17113_/X _17114_/X _17094_/X _15408_/Y vssd1 vssd1 vccd1 vccd1
+ _17115_/X sky130_fd_sc_hd__a32o_1
X_14327_ _12166_/X _12809_/B _14330_/S vssd1 vssd1 vccd1 vccd1 _14327_/X sky130_fd_sc_hd__mux2_1
X_18095_ _22870_/Q _18081_/X _18094_/X _18090_/X vssd1 vssd1 vccd1 vccd1 _22870_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_305_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11539_ _11288_/A _11521_/X _11529_/X _11538_/X _11483_/A vssd1 vssd1 vccd1 vccd1
+ _11552_/B sky130_fd_sc_hd__a311o_1
XFILLER_172_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_356_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_317_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17046_ _13910_/X _17044_/X _17087_/S vssd1 vssd1 vccd1 vccd1 _17046_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14258_ _14760_/A vssd1 vssd1 vccd1 vccd1 _14259_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_356_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13209_ _13202_/Y _13204_/Y _13206_/Y _13208_/Y _11246_/A vssd1 vssd1 vccd1 vccd1
+ _13210_/B sky130_fd_sc_hd__o221a_1
XFILLER_174_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14189_ _21335_/B _14815_/B _14815_/C vssd1 vssd1 vccd1 vccd1 _21443_/A sky130_fd_sc_hd__nand3_4
XFILLER_286_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _16886_/X _23195_/Q _19001_/S vssd1 vssd1 vccd1 vccd1 _18998_/A sky130_fd_sc_hd__mux2_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _18029_/A vssd1 vssd1 vccd1 vccd1 _17948_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_305_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17879_ _17879_/A vssd1 vssd1 vccd1 vccd1 _22810_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_281_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19618_ _19618_/A vssd1 vssd1 vccd1 vccd1 _23456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20890_ _20890_/A _20890_/B vssd1 vssd1 vccd1 vccd1 _20895_/B sky130_fd_sc_hd__nor2_2
XFILLER_326_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19549_ _19258_/X _23426_/Q _19549_/S vssd1 vssd1 vccd1 vccd1 _19550_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22560_ _22977_/CLK _22560_/D vssd1 vssd1 vccd1 vccd1 _22560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21511_ _21509_/Y _21511_/B vssd1 vssd1 vccd1 vccd1 _21514_/A sky130_fd_sc_hd__and2b_1
XFILLER_194_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22491_ _23841_/CLK _22491_/D vssd1 vssd1 vccd1 vccd1 _22491_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_349_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_15_0_wb_clk_i clkbuf_3_7_1_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_15_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_309_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21442_ _21520_/A _21442_/B vssd1 vssd1 vccd1 vccd1 _21442_/Y sky130_fd_sc_hd__nor2_1
XFILLER_348_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21373_ _21373_/A _21373_/B vssd1 vssd1 vccd1 vccd1 _21374_/B sky130_fd_sc_hd__xnor2_1
XFILLER_108_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_324_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_292_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23112_ _23368_/CLK _23112_/D vssd1 vssd1 vccd1 vccd1 _23112_/Q sky130_fd_sc_hd__dfxtp_1
X_20324_ _20324_/A vssd1 vssd1 vccd1 vccd1 _20324_/X sky130_fd_sc_hd__buf_2
XFILLER_351_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_323_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23043_ _23555_/CLK _23043_/D vssd1 vssd1 vccd1 vccd1 _23043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_333_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20255_ _21648_/A _20279_/B vssd1 vssd1 vccd1 vccd1 _20255_/Y sky130_fd_sc_hd__nand2_1
XFILLER_320_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_289_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_288_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20186_ _20186_/A _20186_/B vssd1 vssd1 vccd1 vccd1 _20220_/A sky130_fd_sc_hd__nor2_1
XTAP_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23945_ _23945_/CLK _23945_/D vssd1 vssd1 vccd1 vccd1 _23945_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_291_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _11890_/A _11890_/B vssd1 vssd1 vccd1 vccd1 _11890_/Y sky130_fd_sc_hd__nor2_1
X_23876_ _23876_/CLK _23876_/D vssd1 vssd1 vccd1 vccd1 _23876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_301_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22827_ _22830_/CLK _22827_/D vssd1 vssd1 vccd1 vccd1 _22827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_260_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13560_ _13569_/A _13569_/B _15996_/A vssd1 vssd1 vccd1 vccd1 _13561_/B sky130_fd_sc_hd__a21oi_2
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22758_ _23570_/CLK _22758_/D vssd1 vssd1 vccd1 vccd1 _22758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12511_ _12511_/A _12511_/B vssd1 vssd1 vccd1 vccd1 _12511_/X sky130_fd_sc_hd__or2_1
X_21709_ _21709_/A _21709_/B vssd1 vssd1 vccd1 vccd1 _21711_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13491_ _13491_/A _15996_/A vssd1 vssd1 vccd1 vccd1 _13569_/A sky130_fd_sc_hd__nor2_4
XFILLER_347_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22689_ _23058_/CLK _22689_/D vssd1 vssd1 vccd1 vccd1 _22689_/Q sky130_fd_sc_hd__dfxtp_1
X_15230_ _14898_/X _15206_/X _15228_/X _15229_/X _14937_/X vssd1 vssd1 vccd1 vccd1
+ _15230_/X sky130_fd_sc_hd__o32a_4
XFILLER_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12442_ _11957_/A _12371_/B _12441_/X _12283_/B vssd1 vssd1 vccd1 vccd1 _12443_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15161_ _15161_/A _15161_/B vssd1 vssd1 vccd1 vccd1 _15161_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_354_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12373_ _22264_/Q _23080_/Q _23496_/Q _22425_/Q _12209_/X _12210_/X vssd1 vssd1 vccd1
+ vccd1 _12374_/B sky130_fd_sc_hd__mux4_1
XFILLER_327_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_354_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14112_ _22888_/Q vssd1 vssd1 vccd1 vccd1 _14119_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_315_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11324_ _11365_/A vssd1 vssd1 vccd1 vccd1 _11469_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15092_ _15292_/S _15091_/Y _14860_/X vssd1 vssd1 vccd1 vccd1 _15092_/X sky130_fd_sc_hd__a21o_1
XFILLER_342_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18920_ _18931_/A vssd1 vssd1 vccd1 vccd1 _18929_/S sky130_fd_sc_hd__buf_2
X_14043_ _14046_/A _14052_/B _14043_/C vssd1 vssd1 vccd1 vccd1 _14043_/X sky130_fd_sc_hd__or3_1
XTAP_7130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11255_ _11884_/B vssd1 vssd1 vccd1 vccd1 _11763_/B sky130_fd_sc_hd__buf_2
XTAP_7141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18851_ _18851_/A vssd1 vssd1 vccd1 vccd1 _23133_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11186_ _11492_/S vssd1 vssd1 vccd1 vccd1 _13434_/A sky130_fd_sc_hd__buf_4
XFILLER_122_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17802_ _22776_/Q _17645_/X _17802_/S vssd1 vssd1 vccd1 vccd1 _17803_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18782_ _18782_/A vssd1 vssd1 vccd1 vccd1 _18782_/X sky130_fd_sc_hd__clkbuf_2
XTAP_6495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15994_ _14755_/X _15981_/X _15993_/X vssd1 vssd1 vccd1 vccd1 _17269_/A sky130_fd_sc_hd__o21ai_4
XTAP_5761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17733_ _17789_/A vssd1 vssd1 vccd1 vccd1 _17802_/S sky130_fd_sc_hd__buf_6
XFILLER_10_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_294_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14945_ _15387_/S vssd1 vssd1 vccd1 vccd1 _15089_/S sky130_fd_sc_hd__clkbuf_2
XTAP_5794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_205_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23950_/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_91_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17664_ _17664_/A vssd1 vssd1 vccd1 vccd1 _22713_/D sky130_fd_sc_hd__clkbuf_1
X_14876_ _14936_/A _14869_/X _14875_/X _14498_/X vssd1 vssd1 vccd1 vccd1 _14876_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19403_ _23361_/Q _18862_/X _19405_/S vssd1 vssd1 vccd1 vccd1 _19404_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_102 _21616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_290_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16615_ _16615_/A vssd1 vssd1 vccd1 vccd1 _22456_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_113 _20264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13827_ _13855_/A _13827_/B vssd1 vssd1 vccd1 vccd1 _13828_/A sky130_fd_sc_hd__and2_1
XINSDIODE2_124 _21386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17595_ _17627_/A vssd1 vssd1 vccd1 vccd1 _17608_/S sky130_fd_sc_hd__clkbuf_8
XINSDIODE2_135 _20347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_146 _20362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19334_ _19334_/A vssd1 vssd1 vccd1 vccd1 _23330_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_157 _16016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_168 _17385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13758_ _13858_/A _13771_/B vssd1 vssd1 vccd1 vccd1 _13758_/X sky130_fd_sc_hd__and2_1
X_16546_ _14984_/X _22426_/Q _16546_/S vssd1 vssd1 vccd1 vccd1 _16547_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_179 _13713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ _12709_/A vssd1 vssd1 vccd1 vccd1 _12709_/X sky130_fd_sc_hd__buf_4
XFILLER_189_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_337_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19265_ _19264_/X _23300_/Q _19265_/S vssd1 vssd1 vccd1 vccd1 _19266_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13689_ _14231_/A vssd1 vssd1 vccd1 vccd1 _14219_/A sky130_fd_sc_hd__buf_2
X_16477_ _16477_/A vssd1 vssd1 vccd1 vccd1 _22396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18216_ _18242_/A vssd1 vssd1 vccd1 vccd1 _18216_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15428_ _21738_/A _15430_/B vssd1 vssd1 vccd1 vccd1 _15529_/C sky130_fd_sc_hd__and2_2
XFILLER_318_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19196_ _19196_/A vssd1 vssd1 vccd1 vccd1 _23278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_318_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_346_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18147_ _18159_/A _18147_/B vssd1 vssd1 vccd1 vccd1 _18148_/A sky130_fd_sc_hd__and2_1
X_15359_ _15346_/A _15352_/X _15358_/Y _15150_/X vssd1 vssd1 vccd1 vccd1 _15360_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_346_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18078_ _22864_/Q _18066_/X _18077_/X _18075_/X vssd1 vssd1 vccd1 vccd1 _22864_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_305_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17029_ input72/X input87/X _17029_/S vssd1 vssd1 vccd1 vccd1 _17029_/X sky130_fd_sc_hd__mux2_8
XFILLER_299_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20040_ _23624_/Q _23623_/Q _20040_/C _20042_/D vssd1 vssd1 vccd1 vccd1 _20056_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_299_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21991_ _23835_/Q _23769_/Q vssd1 vssd1 vccd1 vccd1 _21993_/A sky130_fd_sc_hd__and2_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23730_ _23861_/CLK _23730_/D vssd1 vssd1 vccd1 vccd1 _23730_/Q sky130_fd_sc_hd__dfxtp_1
X_20942_ _23796_/Q _20939_/X _20941_/X _20934_/X vssd1 vssd1 vccd1 vccd1 _23796_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_226_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23661_ _23700_/CLK _23661_/D vssd1 vssd1 vccd1 vccd1 _23661_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20873_ _20879_/A _20873_/B vssd1 vssd1 vccd1 vccd1 _20874_/A sky130_fd_sc_hd__and2_1
X_22612_ _23851_/CLK _22612_/D vssd1 vssd1 vccd1 vccd1 _22612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23592_ _23592_/CLK _23592_/D vssd1 vssd1 vccd1 vccd1 _23592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22543_ _23515_/CLK _22543_/D vssd1 vssd1 vccd1 vccd1 _22543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22474_ _22666_/CLK _22474_/D vssd1 vssd1 vccd1 vccd1 _22474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_337_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21425_ _21425_/A _21425_/B vssd1 vssd1 vccd1 vccd1 _21425_/X sky130_fd_sc_hd__or2_1
XFILLER_336_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21356_ _21301_/B _21289_/A _20774_/A _21191_/A vssd1 vssd1 vccd1 vccd1 _21361_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_190_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20307_ _20307_/A vssd1 vssd1 vccd1 vccd1 _20307_/X sky130_fd_sc_hd__buf_2
X_21287_ _21287_/A _21287_/B vssd1 vssd1 vccd1 vccd1 _22257_/B sky130_fd_sc_hd__and2_1
XFILLER_116_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23026_ _23535_/CLK _23026_/D vssd1 vssd1 vccd1 vccd1 _23026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_311_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20238_ _20344_/A vssd1 vssd1 vccd1 vccd1 _20277_/B sky130_fd_sc_hd__buf_2
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20169_ _20169_/A vssd1 vssd1 vccd1 vccd1 _20169_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12991_ _23933_/Q vssd1 vssd1 vccd1 vccd1 _17224_/A sky130_fd_sc_hd__inv_6
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14730_ _14730_/A vssd1 vssd1 vccd1 vccd1 _14730_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11942_ _13382_/B _11937_/X _13380_/A vssd1 vssd1 vccd1 vccd1 _11943_/B sky130_fd_sc_hd__a21oi_1
XFILLER_217_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23928_ _23942_/CLK _23928_/D vssd1 vssd1 vccd1 vccd1 _23928_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _14350_/X _14339_/X _14664_/S vssd1 vssd1 vccd1 vccd1 _14661_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _12387_/A vssd1 vssd1 vccd1 vccd1 _12410_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23859_ _23862_/CLK _23859_/D vssd1 vssd1 vccd1 vccd1 _23859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _13612_/A _13611_/X vssd1 vssd1 vccd1 vccd1 _13612_/X sky130_fd_sc_hd__or2b_4
X_16400_ _16400_/A vssd1 vssd1 vccd1 vccd1 _22362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ _22610_/Q _13662_/B _17380_/S vssd1 vssd1 vccd1 vccd1 _17381_/A sky130_fd_sc_hd__mux2_1
X_14592_ _14592_/A vssd1 vssd1 vccd1 vccd1 _14592_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16331_ _15240_/X _22333_/Q _16333_/S vssd1 vssd1 vccd1 vccd1 _16332_/A sky130_fd_sc_hd__mux2_1
X_13543_ _13543_/A _13573_/A vssd1 vssd1 vccd1 vccd1 _13543_/Y sky130_fd_sc_hd__nor2_1
XFILLER_319_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16262_ _18827_/A vssd1 vssd1 vccd1 vccd1 _16262_/X sky130_fd_sc_hd__buf_2
XFILLER_201_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19050_ _19050_/A vssd1 vssd1 vccd1 vccd1 _23218_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13474_ _13474_/A _13884_/B vssd1 vssd1 vccd1 vccd1 _13879_/A sky130_fd_sc_hd__nor2_2
X_18001_ _22842_/Q _17981_/X _17999_/X _18000_/X vssd1 vssd1 vccd1 vccd1 _22842_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_328_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15213_ _15905_/B vssd1 vssd1 vccd1 vccd1 _16021_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_346_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12425_ _12425_/A _12425_/B vssd1 vssd1 vccd1 vccd1 _12425_/Y sky130_fd_sc_hd__nand2_1
XFILLER_200_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16193_ _21079_/A _15478_/X _16192_/X vssd1 vssd1 vccd1 vccd1 _16193_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_337_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_315_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15144_ _23788_/Q _14605_/X _14486_/X vssd1 vssd1 vccd1 vccd1 _15144_/X sky130_fd_sc_hd__a21o_1
XFILLER_343_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12356_ _12365_/A _12355_/X _11229_/A vssd1 vssd1 vccd1 vccd1 _12356_/X sky130_fd_sc_hd__o21a_1
XFILLER_153_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput309 _13963_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[14] sky130_fd_sc_hd__buf_2
XFILLER_342_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11307_ _12843_/A vssd1 vssd1 vccd1 vccd1 _11308_/A sky130_fd_sc_hd__buf_4
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19952_ _19987_/A vssd1 vssd1 vccd1 vccd1 _19981_/A sky130_fd_sc_hd__clkbuf_2
X_15075_ _22952_/Q _15074_/X _15835_/B vssd1 vssd1 vccd1 vccd1 _15075_/X sky130_fd_sc_hd__mux2_1
XFILLER_236_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12287_ _12287_/A _12287_/B vssd1 vssd1 vccd1 vccd1 _13510_/B sky130_fd_sc_hd__nor2_2
XFILLER_342_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18903_ _23153_/Q _18811_/X _18907_/S vssd1 vssd1 vccd1 vccd1 _18904_/A sky130_fd_sc_hd__mux2_1
X_14026_ input246/X _14004_/X _14025_/X vssd1 vssd1 vccd1 vccd1 _14026_/X sky130_fd_sc_hd__a21o_4
XFILLER_113_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11238_ _22292_/Q _23108_/Q _23524_/Q _22453_/Q _13434_/A _14393_/A vssd1 vssd1 vccd1
+ vccd1 _11239_/B sky130_fd_sc_hd__mux4_1
XFILLER_353_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19883_ _16262_/X _23574_/Q _19887_/S vssd1 vssd1 vccd1 vccd1 _19884_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_296_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18834_ _23128_/Q _18833_/X _18834_/S vssd1 vssd1 vccd1 vccd1 _18835_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11169_ _11169_/A vssd1 vssd1 vccd1 vccd1 _11200_/A sky130_fd_sc_hd__buf_2
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18765_ _16911_/X _23107_/Q _18767_/S vssd1 vssd1 vccd1 vccd1 _18766_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15977_ _15975_/X _22286_/Q _16125_/S vssd1 vssd1 vccd1 vccd1 _15978_/A sky130_fd_sc_hd__mux2_1
XTAP_5580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17716_ _17716_/A vssd1 vssd1 vccd1 vccd1 _22737_/D sky130_fd_sc_hd__clkbuf_1
X_14928_ _16177_/S vssd1 vssd1 vccd1 vccd1 _15885_/A sky130_fd_sc_hd__buf_2
XFILLER_208_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18696_ _18696_/A vssd1 vssd1 vccd1 vccd1 _23076_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17647_ _17647_/A vssd1 vssd1 vccd1 vccd1 _22709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14859_ _15339_/S _14858_/X _14767_/A vssd1 vssd1 vccd1 vccd1 _14859_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_298_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17578_ _18804_/A vssd1 vssd1 vccd1 vccd1 _17578_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_211_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19317_ _19317_/A vssd1 vssd1 vccd1 vccd1 _23322_/D sky130_fd_sc_hd__clkbuf_1
X_16529_ _16529_/A vssd1 vssd1 vccd1 vccd1 _22420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_338_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_337_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19248_ _19248_/A vssd1 vssd1 vccd1 vccd1 _23294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_326_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19179_ _19178_/X _23273_/Q _19179_/S vssd1 vssd1 vccd1 vccd1 _19180_/A sky130_fd_sc_hd__mux2_1
XFILLER_319_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21210_ _21210_/A vssd1 vssd1 vccd1 vccd1 _23882_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_345_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22190_ _23842_/Q _22190_/B vssd1 vssd1 vccd1 vccd1 _22190_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21141_ _23845_/Q _21148_/A vssd1 vssd1 vccd1 vccd1 _21142_/A sky130_fd_sc_hd__and2_2
Xclkbuf_leaf_198_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _22618_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21072_ _23844_/Q _21072_/B vssd1 vssd1 vccd1 vccd1 _21072_/X sky130_fd_sc_hd__or2_1
XFILLER_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20023_ _20034_/B _20034_/C vssd1 vssd1 vccd1 vccd1 _20025_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_127_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _22947_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21974_ _21951_/B _21953_/B _21951_/A vssd1 vssd1 vccd1 vccd1 _21978_/A sky130_fd_sc_hd__a21bo_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23713_ _23714_/CLK _23713_/D vssd1 vssd1 vccd1 vccd1 _23713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20925_ _20925_/A vssd1 vssd1 vccd1 vccd1 _20925_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23644_ _23652_/CLK _23644_/D vssd1 vssd1 vccd1 vccd1 _23644_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20856_ _20856_/A vssd1 vssd1 vccd1 vccd1 _23770_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23575_ _23575_/CLK _23575_/D vssd1 vssd1 vccd1 vccd1 _23575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_298_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20787_ _20963_/A vssd1 vssd1 vccd1 vccd1 _20948_/A sky130_fd_sc_hd__buf_4
XFILLER_357_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22526_ _23466_/CLK _22526_/D vssd1 vssd1 vccd1 vccd1 _22526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_344_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_343_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22457_ _22618_/CLK _22457_/D vssd1 vssd1 vccd1 vccd1 _22457_/Q sky130_fd_sc_hd__dfxtp_1
X_12210_ _12476_/A vssd1 vssd1 vccd1 vccd1 _12210_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21408_ _21767_/A vssd1 vssd1 vccd1 vccd1 _21408_/X sky130_fd_sc_hd__buf_2
XFILLER_325_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13190_ _22317_/Q _23453_/Q _13190_/S vssd1 vssd1 vccd1 vccd1 _13190_/X sky130_fd_sc_hd__mux2_1
X_22388_ _23577_/CLK _22388_/D vssd1 vssd1 vccd1 vccd1 _22388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_352_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12141_ _12141_/A _12141_/B vssd1 vssd1 vccd1 vccd1 _12141_/X sky130_fd_sc_hd__or2_1
XFILLER_2_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21339_ _21555_/A _21339_/B _21339_/C vssd1 vssd1 vccd1 vccd1 _21339_/X sky130_fd_sc_hd__and3_1
XFILLER_297_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_340_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12072_ _22306_/Q _23442_/Q _12120_/S vssd1 vssd1 vccd1 vccd1 _12073_/B sky130_fd_sc_hd__mux2_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23009_ _23009_/CLK _23009_/D vssd1 vssd1 vccd1 vccd1 _23009_/Q sky130_fd_sc_hd__dfxtp_4
X_15900_ _15900_/A vssd1 vssd1 vccd1 vccd1 _22284_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16880_ _16896_/A vssd1 vssd1 vccd1 vccd1 _16893_/S sky130_fd_sc_hd__buf_4
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_323_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15831_ _15674_/X _15830_/Y _14570_/X vssd1 vssd1 vccd1 vccd1 _15831_/Y sky130_fd_sc_hd__a21oi_2
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_293_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ _23010_/Q _20790_/A _18550_/C _18550_/D vssd1 vssd1 vccd1 vccd1 _18551_/A
+ sky130_fd_sc_hd__and4_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_346_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12974_ _12926_/A _12973_/X _11133_/A vssd1 vssd1 vccd1 vccd1 _12974_/Y sky130_fd_sc_hd__o21ai_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15762_ _23705_/Q _14905_/A _15761_/X vssd1 vssd1 vccd1 vccd1 _15762_/X sky130_fd_sc_hd__o21a_4
XFILLER_206_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _22658_/Q _16246_/X _17505_/S vssd1 vssd1 vccd1 vccd1 _17502_/A sky130_fd_sc_hd__mux2_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14713_ _14713_/A _16980_/A _14713_/C vssd1 vssd1 vccd1 vccd1 _21339_/C sky130_fd_sc_hd__or3_1
X_18481_ _18534_/B vssd1 vssd1 vccd1 vccd1 _18492_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_205_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11925_ _22269_/Q _23085_/Q _23501_/Q _22430_/Q _11799_/X _11800_/X vssd1 vssd1 vccd1
+ vccd1 _11926_/B sky130_fd_sc_hd__mux4_1
X_15693_ _14730_/X _15686_/X _15692_/Y _15150_/X vssd1 vssd1 vccd1 vccd1 _15694_/B
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _22628_/Q _16252_/X _17432_/S vssd1 vssd1 vccd1 vccd1 _17433_/A sky130_fd_sc_hd__mux2_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14644_ _14277_/Y _14282_/X _14646_/S vssd1 vssd1 vccd1 vccd1 _14644_/X sky130_fd_sc_hd__mux2_1
X_11856_ _11849_/Y _11851_/Y _11853_/Y _11855_/Y _11243_/A vssd1 vssd1 vccd1 vccd1
+ _11857_/C sky130_fd_sc_hd__o221a_1
XFILLER_221_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17363_ _22602_/Q input196/X _17369_/S vssd1 vssd1 vccd1 vccd1 _17364_/A sky130_fd_sc_hd__mux2_1
X_14575_ _22512_/Q _14232_/A _14223_/X _14574_/X vssd1 vssd1 vccd1 vccd1 _14576_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_159_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11787_ _11774_/A _11786_/X _12371_/A vssd1 vssd1 vccd1 vccd1 _11787_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_14_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_319_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_348_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19102_ _23241_/Q _18785_/X _19102_/S vssd1 vssd1 vccd1 vccd1 _19103_/A sky130_fd_sc_hd__mux2_1
X_16314_ _14534_/X _22325_/Q _16322_/S vssd1 vssd1 vccd1 vccd1 _16315_/A sky130_fd_sc_hd__mux2_1
X_13526_ _13526_/A _13942_/A vssd1 vssd1 vccd1 vccd1 _13526_/X sky130_fd_sc_hd__or2_1
X_17294_ _17242_/X _17287_/X _17293_/X _16997_/X vssd1 vssd1 vccd1 vccd1 _17294_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_185_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_348_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19033_ _19033_/A vssd1 vssd1 vccd1 vccd1 _23210_/D sky130_fd_sc_hd__clkbuf_1
X_16245_ _16245_/A vssd1 vssd1 vccd1 vccd1 _22304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13457_ _13457_/A vssd1 vssd1 vccd1 vccd1 _16680_/A sky130_fd_sc_hd__clkinv_2
XFILLER_127_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12408_ _12397_/A _12407_/X _11282_/A vssd1 vssd1 vccd1 vccd1 _12408_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_316_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16176_ _15440_/X _16169_/X _16175_/X _14497_/A vssd1 vssd1 vccd1 vccd1 _16176_/X
+ sky130_fd_sc_hd__o22a_1
X_13388_ _13492_/B _13388_/B vssd1 vssd1 vccd1 vccd1 _13388_/Y sky130_fd_sc_hd__nand2_1
XFILLER_353_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_331_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15127_ _15456_/A _14296_/X _14767_/X vssd1 vssd1 vccd1 vccd1 _15127_/Y sky130_fd_sc_hd__o21ai_1
X_12339_ _12110_/S _21444_/A _12338_/Y vssd1 vssd1 vccd1 vccd1 _12340_/B sky130_fd_sc_hd__a21o_2
XFILLER_342_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_303_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_288_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_330_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19935_ _20008_/A _19935_/B _19935_/C vssd1 vssd1 vccd1 vccd1 _23595_/D sky130_fd_sc_hd__nor3_1
X_15058_ _22501_/Q _14232_/A _14238_/A _15057_/X _15179_/A vssd1 vssd1 vccd1 vccd1
+ _15483_/A sky130_fd_sc_hd__o221a_2
XFILLER_130_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_287_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_331_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14009_ _14041_/A vssd1 vssd1 vccd1 vccd1 _14009_/X sky130_fd_sc_hd__buf_2
XFILLER_123_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_296_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19866_ _19866_/A vssd1 vssd1 vccd1 vccd1 _23566_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_295_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18817_ _18817_/A vssd1 vssd1 vccd1 vccd1 _18817_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_295_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19797_ _19797_/A vssd1 vssd1 vccd1 vccd1 _23535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18748_ _16886_/X _23099_/Q _18752_/S vssd1 vssd1 vccd1 vccd1 _18749_/A sky130_fd_sc_hd__mux2_1
XFILLER_255_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18679_ _18679_/A vssd1 vssd1 vccd1 vccd1 _23068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20710_ _12893_/Y _20701_/X _20709_/Y vssd1 vssd1 vccd1 vccd1 _20711_/C sky130_fd_sc_hd__a21oi_2
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21690_ _21559_/B _21690_/B _21690_/C vssd1 vssd1 vccd1 vccd1 _21690_/X sky130_fd_sc_hd__and3b_1
XFILLER_251_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20641_ _20641_/A _20669_/B vssd1 vssd1 vccd1 vccd1 _20645_/B sky130_fd_sc_hd__nor2_2
XFILLER_189_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_338_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23360_ _23554_/CLK _23360_/D vssd1 vssd1 vccd1 vccd1 _23360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20572_ _20732_/A vssd1 vssd1 vccd1 vccd1 _20572_/X sky130_fd_sc_hd__buf_2
XFILLER_220_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_338_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22311_ _22632_/CLK _22311_/D vssd1 vssd1 vccd1 vccd1 _22311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_258_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23291_ _23419_/CLK _23291_/D vssd1 vssd1 vccd1 vccd1 _23291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_325_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22242_ _23844_/Q _22242_/B _22242_/C vssd1 vssd1 vccd1 vccd1 _22242_/X sky130_fd_sc_hd__and3_1
XFILLER_118_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22173_ _21379_/A _22164_/X _22172_/X _21465_/A vssd1 vssd1 vccd1 vccd1 _22173_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_279_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21124_ _21124_/A vssd1 vssd1 vccd1 vccd1 _21124_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21055_ _23836_/Q _20996_/B _21054_/Y _21049_/X vssd1 vssd1 vccd1 vccd1 _23836_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_259_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_290_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20006_ _23614_/Q _23613_/Q vssd1 vssd1 vccd1 vccd1 _20014_/D sky130_fd_sc_hd__and2_1
XFILLER_59_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_290_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_290_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21957_ _21491_/X _21948_/X _21956_/Y vssd1 vssd1 vccd1 vccd1 _21957_/X sky130_fd_sc_hd__a21o_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_95_wb_clk_i _22899_/CLK vssd1 vssd1 vccd1 vccd1 _23489_/CLK sky130_fd_sc_hd__clkbuf_16
X_11710_ _11621_/X _11709_/X _12256_/A vssd1 vssd1 vccd1 vccd1 _11710_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _20936_/A vssd1 vssd1 vccd1 vccd1 _20908_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _23320_/Q _23288_/Q _23256_/Q _23544_/Q _12977_/S _12685_/X vssd1 vssd1 vccd1
+ vccd1 _12691_/B sky130_fd_sc_hd__mux4_2
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21888_ _21888_/A _21888_/B vssd1 vssd1 vccd1 vccd1 _21889_/B sky130_fd_sc_hd__or2_1
XFILLER_299_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23555_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23627_ _23632_/CLK _23627_/D vssd1 vssd1 vccd1 vccd1 _23627_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_306_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11641_ _11986_/A _11641_/B vssd1 vssd1 vccd1 vccd1 _11641_/X sky130_fd_sc_hd__or2_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20839_ _20683_/B _20828_/X _20829_/X _23766_/Q vssd1 vssd1 vccd1 vccd1 _20840_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_357_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14360_ _14351_/S _14359_/X _14840_/S vssd1 vssd1 vccd1 vccd1 _14360_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_345_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_320_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23558_ _23558_/CLK _23558_/D vssd1 vssd1 vccd1 vccd1 _23558_/Q sky130_fd_sc_hd__dfxtp_1
X_11572_ _12556_/A vssd1 vssd1 vccd1 vccd1 _11719_/A sky130_fd_sc_hd__buf_4
XFILLER_211_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_317_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13311_ _13311_/A _13316_/B vssd1 vssd1 vccd1 vccd1 _13311_/X sky130_fd_sc_hd__or2_1
XFILLER_357_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22509_ _23693_/CLK _22509_/D vssd1 vssd1 vccd1 vccd1 _22509_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput19 core_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_317_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14291_ _14286_/X _14373_/A _14369_/A vssd1 vssd1 vccd1 vccd1 _14291_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23489_ _23489_/CLK _23489_/D vssd1 vssd1 vccd1 vccd1 _23489_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16030_ _15003_/X _16018_/X _16029_/X vssd1 vssd1 vccd1 vccd1 _17279_/A sky130_fd_sc_hd__o21ai_4
X_13242_ _13242_/A _13242_/B vssd1 vssd1 vccd1 vccd1 _13242_/X sky130_fd_sc_hd__and2_1
XFILLER_136_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_331_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13173_ _13216_/A _13170_/X _13172_/X _11352_/A vssd1 vssd1 vccd1 vccd1 _13173_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_340_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12124_ _11131_/A _12115_/Y _12117_/Y _12123_/Y _11216_/A vssd1 vssd1 vccd1 vccd1
+ _12134_/B sky130_fd_sc_hd__o311a_1
XFILLER_151_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17981_ _17981_/A vssd1 vssd1 vccd1 vccd1 _17981_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19720_ _19720_/A vssd1 vssd1 vccd1 vccd1 _23501_/D sky130_fd_sc_hd__clkbuf_1
X_12055_ _22275_/Q _23091_/Q _23507_/Q _22436_/Q _11972_/X _11973_/X vssd1 vssd1 vccd1
+ vccd1 _12056_/B sky130_fd_sc_hd__mux4_1
X_16932_ _16932_/A vssd1 vssd1 vccd1 vccd1 _17648_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_238_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19651_ _19697_/S vssd1 vssd1 vccd1 vccd1 _19660_/S sky130_fd_sc_hd__clkbuf_4
X_16863_ _19213_/A vssd1 vssd1 vccd1 vccd1 _16863_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_293_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18602_ _16883_/X _23034_/Q _18608_/S vssd1 vssd1 vccd1 vccd1 _18603_/A sky130_fd_sc_hd__mux2_1
XFILLER_265_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15814_ _14431_/A _15803_/X _15812_/X _15813_/X _14518_/A vssd1 vssd1 vccd1 vccd1
+ _15815_/B sky130_fd_sc_hd__o32a_4
XFILLER_293_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19582_ _23440_/Q _19201_/A _19588_/S vssd1 vssd1 vccd1 vccd1 _19583_/A sky130_fd_sc_hd__mux2_1
X_16794_ _22515_/Q _16783_/X _16784_/X input30/X vssd1 vssd1 vccd1 vccd1 _16795_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18533_ _18480_/A _18532_/Y _18264_/A vssd1 vssd1 vccd1 vccd1 _23008_/D sky130_fd_sc_hd__a21oi_1
XFILLER_80_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_350_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15745_ _22997_/Q _15780_/A _15781_/A input225/X vssd1 vssd1 vccd1 vccd1 _21920_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_19_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _23417_/Q _23033_/Q _23385_/Q _23353_/Q _12029_/X _12009_/X vssd1 vssd1 vccd1
+ vccd1 _12958_/B sky130_fd_sc_hd__mux4_2
XFILLER_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18464_ _18451_/X _18462_/Y _18463_/X vssd1 vssd1 vccd1 vccd1 _22981_/D sky130_fd_sc_hd__a21oi_1
XFILLER_261_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11908_ _11901_/Y _11903_/Y _11905_/Y _11907_/Y _11244_/A vssd1 vssd1 vccd1 vccd1
+ _11909_/C sky130_fd_sc_hd__o221a_1
XFILLER_221_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ _15676_/A vssd1 vssd1 vccd1 vccd1 _15676_/X sky130_fd_sc_hd__buf_2
X_12888_ _12871_/A _12887_/X _11232_/A vssd1 vssd1 vccd1 vccd1 _12888_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_261_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17415_ _22620_/Q _16227_/X _17421_/S vssd1 vssd1 vccd1 vccd1 _17416_/A sky130_fd_sc_hd__mux2_1
X_14627_ _14854_/S _14626_/X _14376_/X vssd1 vssd1 vccd1 vccd1 _14627_/X sky130_fd_sc_hd__o21a_1
X_18395_ _18403_/A _18400_/C vssd1 vssd1 vccd1 vccd1 _18395_/Y sky130_fd_sc_hd__nor2_1
X_11839_ _11839_/A _11839_/B vssd1 vssd1 vccd1 vccd1 _11839_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_348_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17346_ _17346_/A vssd1 vssd1 vccd1 vccd1 _22594_/D sky130_fd_sc_hd__clkbuf_1
X_14558_ _16203_/B _16457_/B _16457_/C vssd1 vssd1 vccd1 vccd1 _19627_/A sky130_fd_sc_hd__or3b_2
XFILLER_146_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13509_ _13503_/Y _14794_/A _13902_/B _13508_/Y vssd1 vssd1 vccd1 vccd1 _13906_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_347_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17277_ input97/X input62/X _17314_/S vssd1 vssd1 vccd1 vccd1 _17277_/X sky130_fd_sc_hd__mux2_8
X_14489_ _21097_/A _20989_/B vssd1 vssd1 vccd1 vccd1 _20409_/A sky130_fd_sc_hd__or2_4
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19016_ _16914_/X _23204_/Q _19016_/S vssd1 vssd1 vccd1 vccd1 _19017_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16228_ _22299_/Q _16227_/X _16237_/S vssd1 vssd1 vccd1 vccd1 _16229_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16159_ _16156_/X _16157_/X _22224_/A _15708_/S vssd1 vssd1 vccd1 vccd1 _18868_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_304_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19918_ _19915_/X _19916_/X _19917_/Y vssd1 vssd1 vccd1 vccd1 _23589_/D sky130_fd_sc_hd__o21a_1
XFILLER_275_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19849_ _19849_/A vssd1 vssd1 vccd1 vccd1 _23558_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_284_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22860_ _22923_/CLK _22860_/D vssd1 vssd1 vccd1 vccd1 _22860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21811_ _21812_/B _21934_/A vssd1 vssd1 vccd1 vccd1 _21853_/B sky130_fd_sc_hd__and2b_1
XFILLER_272_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22791_ _23578_/CLK _22791_/D vssd1 vssd1 vccd1 vccd1 _22791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21742_ _21569_/X _21740_/X _21741_/Y _21577_/X vssd1 vssd1 vccd1 vccd1 _21743_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_52_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21673_ _21673_/A _21676_/A vssd1 vssd1 vccd1 vccd1 _21674_/B sky130_fd_sc_hd__nor2_1
XFILLER_225_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23412_ _23414_/CLK _23412_/D vssd1 vssd1 vccd1 vccd1 _23412_/Q sky130_fd_sc_hd__dfxtp_1
X_20624_ _14541_/X _20773_/A _20574_/X vssd1 vssd1 vccd1 vccd1 _20624_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_178_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23343_ _23407_/CLK _23343_/D vssd1 vssd1 vccd1 vccd1 _23343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20555_ _14468_/B _20143_/A _21308_/B vssd1 vssd1 vccd1 vccd1 _20730_/A sky130_fd_sc_hd__o21a_2
XFILLER_137_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23274_ _23466_/CLK _23274_/D vssd1 vssd1 vccd1 vccd1 _23274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20486_ _20749_/A _20467_/X _20485_/X _20483_/X vssd1 vssd1 vccd1 vccd1 _23713_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_142_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _23851_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_146_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22225_ _21398_/X _22223_/X _22224_/Y _21408_/X vssd1 vssd1 vccd1 vccd1 _22225_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_180_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_350_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22156_ _22161_/A _22127_/B _22102_/Y _22101_/A vssd1 vssd1 vccd1 vccd1 _22156_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_6814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput470 _23929_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[18] sky130_fd_sc_hd__buf_2
XFILLER_350_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21107_ _23851_/Q _21096_/X _21098_/X _20588_/A vssd1 vssd1 vccd1 vccd1 _21108_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xoutput481 _23939_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[28] sky130_fd_sc_hd__buf_2
Xoutput492 _23920_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[9] sky130_fd_sc_hd__buf_2
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22087_ _22087_/A _22087_/B vssd1 vssd1 vccd1 vccd1 _22087_/Y sky130_fd_sc_hd__nor2_1
XTAP_6869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_304_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21038_ _20675_/A _21027_/X _21035_/X _21037_/X vssd1 vssd1 vccd1 vccd1 _23829_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_75_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13860_ _13857_/X _13858_/X _13859_/X vssd1 vssd1 vccd1 vccd1 _14064_/C sky130_fd_sc_hd__o21ai_4
X_12811_ _13608_/A _12664_/A _12636_/X _11691_/B _13536_/A vssd1 vssd1 vccd1 vccd1
+ _12812_/B sky130_fd_sc_hd__a32o_1
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22989_ _23009_/CLK _22989_/D vssd1 vssd1 vccd1 vccd1 _22989_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_250_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_509 _17232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13791_ _13808_/A vssd1 vssd1 vccd1 vccd1 _13798_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15530_ _21762_/A _15529_/C _21791_/A vssd1 vssd1 vccd1 vccd1 _15531_/B sky130_fd_sc_hd__a21oi_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12742_/A _12807_/A vssd1 vssd1 vccd1 vccd1 _12743_/B sky130_fd_sc_hd__nand2_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12673_ _12820_/S vssd1 vssd1 vccd1 vccd1 _12819_/S sky130_fd_sc_hd__buf_4
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15461_ _12113_/B _15583_/A _14793_/A _12162_/Y _15460_/Y vssd1 vssd1 vccd1 vccd1
+ _15461_/X sky130_fd_sc_hd__o221a_1
XFILLER_179_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17200_ input90/X input55/X _17200_/S vssd1 vssd1 vccd1 vccd1 _17200_/X sky130_fd_sc_hd__mux2_8
X_11624_ _11141_/A _11620_/X _11623_/X _11131_/A vssd1 vssd1 vccd1 vccd1 _11624_/X
+ sky130_fd_sc_hd__o211a_1
X_14412_ _22907_/Q _14153_/X _14151_/X _22600_/Q vssd1 vssd1 vccd1 vccd1 _14552_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18180_ _18144_/B _18167_/X _18178_/X _18179_/Y vssd1 vssd1 vccd1 vccd1 _18180_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_187_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15392_ _13379_/C _16180_/B _15391_/Y _20532_/A vssd1 vssd1 vccd1 vccd1 _15392_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_357_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17131_ _17324_/A vssd1 vssd1 vccd1 vccd1 _17131_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14343_ _12233_/B _13241_/A _14343_/S vssd1 vssd1 vccd1 vccd1 _14343_/X sky130_fd_sc_hd__mux2_1
X_11555_ _11555_/A vssd1 vssd1 vccd1 vccd1 _11557_/B sky130_fd_sc_hd__inv_2
XFILLER_317_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_305_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17062_ _17231_/A vssd1 vssd1 vccd1 vccd1 _17062_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14274_ _14326_/S _14274_/B vssd1 vssd1 vccd1 vccd1 _14274_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11486_ _23941_/Q _11486_/B vssd1 vssd1 vccd1 vccd1 _11486_/X sky130_fd_sc_hd__or2_1
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16013_ _19249_/A vssd1 vssd1 vccd1 vccd1 _16013_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_326_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13225_ _13225_/A _13225_/B vssd1 vssd1 vccd1 vccd1 _13225_/X sky130_fd_sc_hd__or2_1
XFILLER_344_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_345_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_313_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13156_ _13199_/A _13155_/X _11134_/A vssd1 vssd1 vccd1 vccd1 _13156_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_312_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12107_ _12028_/A _12106_/X _11681_/A vssd1 vssd1 vccd1 vccd1 _12107_/X sky130_fd_sc_hd__o21a_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17964_ _22832_/Q _17950_/X _17962_/X _17963_/X vssd1 vssd1 vccd1 vccd1 _22832_/D
+ sky130_fd_sc_hd__o211a_1
X_13087_ _13149_/A _13087_/B vssd1 vssd1 vccd1 vccd1 _13087_/Y sky130_fd_sc_hd__nor2_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_300_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19703_ _19703_/A vssd1 vssd1 vccd1 vccd1 _23493_/D sky130_fd_sc_hd__clkbuf_1
X_16915_ _16914_/X _22552_/Q _16915_/S vssd1 vssd1 vccd1 vccd1 _16916_/A sky130_fd_sc_hd__mux2_1
X_12038_ _23925_/Q _20279_/A _12739_/A vssd1 vssd1 vccd1 vccd1 _12168_/B sky130_fd_sc_hd__mux2_8
XFILLER_239_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17895_ _17908_/A _17971_/A vssd1 vssd1 vccd1 vccd1 _17986_/A sky130_fd_sc_hd__nor2_1
XFILLER_266_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19634_ _19172_/X _23463_/Q _19638_/S vssd1 vssd1 vccd1 vccd1 _19635_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16846_ _16846_/A vssd1 vssd1 vccd1 vccd1 _22530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_265_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19565_ _19565_/A vssd1 vssd1 vccd1 vccd1 _23432_/D sky130_fd_sc_hd__clkbuf_1
X_16777_ _16777_/A _16777_/B vssd1 vssd1 vccd1 vccd1 _16778_/A sky130_fd_sc_hd__or2_1
XFILLER_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13989_ _13990_/A _14085_/A vssd1 vssd1 vccd1 vccd1 _13989_/Y sky130_fd_sc_hd__nor2_8
XFILLER_92_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18516_ _18516_/A vssd1 vssd1 vccd1 vccd1 _18516_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_207_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15728_ _23672_/Q _16170_/B vssd1 vssd1 vccd1 vccd1 _15728_/X sky130_fd_sc_hd__or2_1
XFILLER_80_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19496_ _19553_/S vssd1 vssd1 vccd1 vccd1 _19505_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_280_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18447_ _22977_/Q _18445_/B _18423_/X vssd1 vssd1 vccd1 vccd1 _18447_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_34_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15659_ _23928_/Q vssd1 vssd1 vccd1 vccd1 _21856_/A sky130_fd_sc_hd__buf_4
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18378_ _18403_/A _18384_/C vssd1 vssd1 vccd1 vccd1 _18378_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17329_ _22587_/Q input190/X _17335_/S vssd1 vssd1 vccd1 vccd1 _17330_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_335_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20340_ _20340_/A _20340_/B vssd1 vssd1 vccd1 vccd1 _20340_/X sky130_fd_sc_hd__or2_1
XFILLER_146_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20271_ _23665_/Q _20165_/X _20270_/Y _20246_/X vssd1 vssd1 vccd1 vccd1 _23665_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_351_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_304_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22010_ _22205_/A _22041_/C vssd1 vssd1 vccd1 vccd1 _22010_/Y sky130_fd_sc_hd__nand2_1
XFILLER_255_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_288_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_331_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_288_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput209 localMemory_wb_adr_i[5] vssd1 vssd1 vccd1 vccd1 input209/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22912_ _22956_/CLK _22912_/D vssd1 vssd1 vccd1 vccd1 _22912_/Q sky130_fd_sc_hd__dfxtp_1
X_23892_ _23893_/CLK _23892_/D vssd1 vssd1 vccd1 vccd1 _23892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22843_ _22893_/CLK _22843_/D vssd1 vssd1 vccd1 vccd1 _22843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22774_ _23585_/CLK _22774_/D vssd1 vssd1 vccd1 vccd1 _22774_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21725_ _21688_/B _21725_/B vssd1 vssd1 vccd1 vccd1 _21725_/X sky130_fd_sc_hd__and2b_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_358_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_358_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21656_ _21618_/Y _21619_/X _14180_/B _21605_/B vssd1 vssd1 vccd1 vccd1 _21694_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_303_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_296_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20607_ _13923_/B _20563_/X _20606_/X vssd1 vssd1 vccd1 vccd1 _20608_/C sky130_fd_sc_hd__o21a_1
XFILLER_339_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21587_ _21587_/A _21587_/B vssd1 vssd1 vccd1 vccd1 _21587_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_137_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_327_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23326_ _23391_/CLK _23326_/D vssd1 vssd1 vccd1 vccd1 _23326_/Q sky130_fd_sc_hd__dfxtp_1
X_11340_ _13291_/A _11340_/B vssd1 vssd1 vccd1 vccd1 _11340_/X sky130_fd_sc_hd__or2_1
X_20538_ _21308_/B vssd1 vssd1 vccd1 vccd1 _20759_/B sky130_fd_sc_hd__buf_2
XFILLER_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_354_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_308_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23257_ _23545_/CLK _23257_/D vssd1 vssd1 vccd1 vccd1 _23257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_314_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_298_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11271_ _23898_/Q vssd1 vssd1 vccd1 vccd1 _11272_/A sky130_fd_sc_hd__clkinv_4
XFILLER_341_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20469_ _20708_/A _20467_/X _20468_/X _20459_/X vssd1 vssd1 vccd1 vccd1 _23706_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13010_ _13184_/A _13010_/B _13010_/C vssd1 vssd1 vccd1 vccd1 _20340_/A sky130_fd_sc_hd__nand3_4
XTAP_7323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22208_ _23811_/Q _21381_/X _22207_/Y _21395_/X vssd1 vssd1 vccd1 vccd1 _22208_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_7334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23188_ _23543_/CLK _23188_/D vssd1 vssd1 vccd1 vccd1 _23188_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22139_ _22139_/A _22139_/B vssd1 vssd1 vccd1 vccd1 _22168_/A sky130_fd_sc_hd__nor2_1
XTAP_7389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14961_ _22491_/Q _14232_/X _14247_/X _14960_/X _14072_/A vssd1 vssd1 vccd1 vccd1
+ _14961_/X sky130_fd_sc_hd__o221a_1
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16700_ _22489_/Q _16689_/X _16693_/X input32/X vssd1 vssd1 vccd1 vccd1 _16701_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13912_ _13355_/A _13911_/X _12600_/A vssd1 vssd1 vccd1 vccd1 _13913_/B sky130_fd_sc_hd__a21oi_2
XTAP_5987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17680_ _22721_/Q _17572_/X _17682_/S vssd1 vssd1 vccd1 vccd1 _17681_/A sky130_fd_sc_hd__mux2_1
XTAP_5998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14892_ _18782_/A vssd1 vssd1 vccd1 vccd1 _19175_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16631_ _16677_/S vssd1 vssd1 vccd1 vccd1 _16640_/S sky130_fd_sc_hd__buf_4
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13843_ _13163_/B _13808_/X _13781_/X vssd1 vssd1 vccd1 vccd1 _13843_/X sky130_fd_sc_hd__a21o_1
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_306 _15990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_290_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19350_ _23337_/Q _18785_/X _19350_/S vssd1 vssd1 vccd1 vccd1 _19351_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_317 _17289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_328 _17298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16562_ _15372_/X _22433_/Q _16568_/S vssd1 vssd1 vccd1 vccd1 _16563_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13774_ _14675_/A vssd1 vssd1 vccd1 vccd1 _13775_/A sky130_fd_sc_hd__buf_4
XINSDIODE2_339 _17112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18301_ _22926_/Q _18297_/C _18300_/Y vssd1 vssd1 vccd1 vccd1 _22926_/D sky130_fd_sc_hd__o21a_1
X_15513_ _22928_/Q _16168_/B _15501_/X _15512_/Y _14897_/A vssd1 vssd1 vccd1 vccd1
+ _15513_/X sky130_fd_sc_hd__a221o_1
X_12725_ _12995_/A _12725_/B vssd1 vssd1 vccd1 vccd1 _12725_/X sky130_fd_sc_hd__or2_1
XFILLER_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19281_ _19181_/X _23306_/Q _19289_/S vssd1 vssd1 vccd1 vccd1 _19282_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16493_ _16515_/A vssd1 vssd1 vccd1 vccd1 _16502_/S sky130_fd_sc_hd__buf_6
X_18232_ _18245_/A vssd1 vssd1 vccd1 vccd1 _18232_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15444_ _23730_/Q _23860_/Q _16138_/S vssd1 vssd1 vccd1 vccd1 _15444_/X sky130_fd_sc_hd__mux2_1
X_12656_ _12656_/A vssd1 vssd1 vccd1 vccd1 _12683_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18163_ _18163_/A _18163_/B _22893_/Q vssd1 vssd1 vccd1 vccd1 _18164_/B sky130_fd_sc_hd__nor3b_1
X_11607_ _11723_/A vssd1 vssd1 vccd1 vccd1 _12656_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12587_ _23209_/Q _23177_/Q _23145_/Q _23113_/Q _12324_/X _12325_/X vssd1 vssd1 vccd1
+ vccd1 _12587_/X sky130_fd_sc_hd__mux4_1
X_15375_ _15478_/A vssd1 vssd1 vccd1 vccd1 _15375_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_357_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_317_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17114_ _17231_/A vssd1 vssd1 vccd1 vccd1 _17114_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_345_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14326_ _12163_/Y _12807_/Y _14326_/S vssd1 vssd1 vccd1 vccd1 _14326_/X sky130_fd_sc_hd__mux2_1
X_18094_ _22869_/Q _18082_/X _18083_/X _23002_/Q _18084_/X vssd1 vssd1 vccd1 vccd1
+ _18094_/X sky130_fd_sc_hd__a221o_1
X_11538_ _13064_/A _11530_/X _11536_/X _11537_/X vssd1 vssd1 vccd1 vccd1 _11538_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_305_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_7_1_wb_clk_i clkbuf_3_7_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_1_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
X_17045_ _17250_/A vssd1 vssd1 vccd1 vccd1 _17087_/S sky130_fd_sc_hd__clkbuf_2
X_11469_ _11469_/A vssd1 vssd1 vccd1 vccd1 _15616_/A sky130_fd_sc_hd__buf_8
X_14257_ _14651_/A vssd1 vssd1 vccd1 vccd1 _14351_/S sky130_fd_sc_hd__buf_2
XFILLER_172_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13208_ _13199_/A _13207_/X _11133_/A vssd1 vssd1 vccd1 vccd1 _13208_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14188_ _14196_/A _14196_/B _14713_/C _21335_/B vssd1 vssd1 vccd1 vccd1 _21555_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_112_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_313_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_286_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13139_ _13542_/A _13139_/B vssd1 vssd1 vccd1 vccd1 _15996_/A sky130_fd_sc_hd__nor2_4
X_18996_ _18996_/A vssd1 vssd1 vccd1 vccd1 _23194_/D sky130_fd_sc_hd__clkbuf_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17947_ _21220_/A vssd1 vssd1 vccd1 vccd1 _18029_/A sky130_fd_sc_hd__buf_4
XFILLER_239_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17878_ _22810_/Q input248/X _17882_/S vssd1 vssd1 vccd1 vccd1 _17879_/A sky130_fd_sc_hd__mux2_1
XFILLER_253_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19617_ _23456_/Q _19252_/A _19621_/S vssd1 vssd1 vccd1 vccd1 _19618_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16829_ _16828_/X _22525_/Q _16829_/S vssd1 vssd1 vccd1 vccd1 _16830_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_326_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19548_ _19548_/A vssd1 vssd1 vccd1 vccd1 _23425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_326_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19479_ _23395_/Q _18868_/X _19481_/S vssd1 vssd1 vccd1 vccd1 _19480_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21510_ _21522_/A _21515_/A vssd1 vssd1 vccd1 vccd1 _21511_/B sky130_fd_sc_hd__nand2_1
XFILLER_221_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22490_ _23841_/CLK _22490_/D vssd1 vssd1 vccd1 vccd1 _22490_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_142_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_349_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21441_ _21441_/A vssd1 vssd1 vccd1 vccd1 _21619_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_336_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_309_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21372_ _21372_/A _21372_/B vssd1 vssd1 vccd1 vccd1 _21373_/B sky130_fd_sc_hd__nand2_1
XFILLER_162_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23111_ _23367_/CLK _23111_/D vssd1 vssd1 vccd1 vccd1 _23111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_351_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20323_ _20323_/A _21153_/A vssd1 vssd1 vccd1 vccd1 _20323_/Y sky130_fd_sc_hd__nand2_1
XFILLER_323_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_292_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_305_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23042_ _23489_/CLK _23042_/D vssd1 vssd1 vccd1 vccd1 _23042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20254_ _20254_/A vssd1 vssd1 vccd1 vccd1 _20295_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_289_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20185_ _20146_/X _20570_/A _20184_/X _18547_/X vssd1 vssd1 vccd1 vccd1 _23655_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23944_ _23946_/CLK _23944_/D vssd1 vssd1 vccd1 vccd1 _23944_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23875_ _23876_/CLK _23875_/D vssd1 vssd1 vccd1 vccd1 _23875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_301_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22826_ _22830_/CLK _22826_/D vssd1 vssd1 vccd1 vccd1 _22826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22757_ _22789_/CLK _22757_/D vssd1 vssd1 vccd1 vccd1 _22757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_340_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12510_ _22357_/Q _22389_/Q _22678_/Q _23045_/Q _23894_/Q _23895_/Q vssd1 vssd1 vccd1
+ vccd1 _12511_/B sky130_fd_sc_hd__mux4_2
XFILLER_40_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21708_ _21708_/A _21708_/B vssd1 vssd1 vccd1 vccd1 _21709_/B sky130_fd_sc_hd__or2_1
X_13490_ _13490_/A vssd1 vssd1 vccd1 vccd1 _13490_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_201_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22688_ _23047_/CLK _22688_/D vssd1 vssd1 vccd1 vccd1 _22688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12441_ _11404_/A _13710_/A _12440_/X vssd1 vssd1 vccd1 vccd1 _12441_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21639_ _23920_/Q _21594_/A _21638_/X vssd1 vssd1 vccd1 vccd1 _21640_/B sky130_fd_sc_hd__o21ai_2
XFILLER_166_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_327_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_355_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12372_ _12344_/X _12368_/X _12370_/Y _12371_/X _11935_/B vssd1 vssd1 vccd1 vccd1
+ _14313_/A sky130_fd_sc_hd__o311ai_4
X_15160_ _15274_/C _15160_/B vssd1 vssd1 vccd1 vccd1 _15161_/B sky130_fd_sc_hd__or2_1
XFILLER_181_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_314_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14111_ _22889_/Q vssd1 vssd1 vccd1 vccd1 _14119_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11323_ _11323_/A vssd1 vssd1 vccd1 vccd1 _11365_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_180_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15091_ _15456_/A _14649_/X _14767_/X vssd1 vssd1 vccd1 vccd1 _15091_/Y sky130_fd_sc_hd__o21ai_2
X_23309_ _23565_/CLK _23309_/D vssd1 vssd1 vccd1 vccd1 _23309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_354_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14042_ _14023_/X _13786_/B _14041_/X input222/X vssd1 vssd1 vccd1 vccd1 _14042_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_69_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11254_ _12206_/A vssd1 vssd1 vccd1 vccd1 _11884_/B sky130_fd_sc_hd__buf_4
XFILLER_107_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18850_ _23133_/Q _18849_/X _18850_/S vssd1 vssd1 vccd1 vccd1 _18851_/A sky130_fd_sc_hd__mux2_1
XTAP_7164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11185_ _11493_/S vssd1 vssd1 vccd1 vccd1 _11492_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_192_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17801_ _17801_/A vssd1 vssd1 vccd1 vccd1 _22775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18781_ _18781_/A vssd1 vssd1 vccd1 vccd1 _23111_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15993_ _22940_/Q _14988_/B _15982_/X _15992_/Y _14898_/A vssd1 vssd1 vccd1 vccd1
+ _15993_/X sky130_fd_sc_hd__a221o_1
XFILLER_95_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17732_ _19164_/A _17804_/B vssd1 vssd1 vccd1 vccd1 _17789_/A sky130_fd_sc_hd__nor2_8
XTAP_5773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14944_ _13906_/A _14942_/X _14943_/Y _12600_/B vssd1 vssd1 vccd1 vccd1 _14958_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_5784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_349_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17663_ _22713_/Q _17544_/X _17671_/S vssd1 vssd1 vccd1 vccd1 _17664_/A sky130_fd_sc_hd__mux2_1
X_14875_ _23688_/Q _14494_/S _14874_/X vssd1 vssd1 vccd1 vccd1 _14875_/X sky130_fd_sc_hd__o21a_2
XFILLER_47_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19402_ _19402_/A vssd1 vssd1 vccd1 vccd1 _23360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16614_ _22456_/Q _16214_/X _16618_/S vssd1 vssd1 vccd1 vccd1 _16615_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_103 _21616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13826_ _13736_/B _13771_/X _13824_/X _13874_/B vssd1 vssd1 vccd1 vccd1 _13827_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_62_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17594_ _18820_/A vssd1 vssd1 vccd1 vccd1 _17594_/X sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_114 _20264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_125 _21386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_136 _20347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19333_ _19258_/X _23330_/Q _19333_/S vssd1 vssd1 vccd1 vccd1 _19334_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_147 _20362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16545_ _16545_/A vssd1 vssd1 vccd1 vccd1 _22425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_349_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_158 _19969_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13757_ _13757_/A vssd1 vssd1 vccd1 vccd1 _13757_/X sky130_fd_sc_hd__buf_2
XINSDIODE2_169 _17385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12708_ _12708_/A vssd1 vssd1 vccd1 vccd1 _12953_/A sky130_fd_sc_hd__buf_2
XFILLER_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19264_ _19264_/A vssd1 vssd1 vccd1 vccd1 _19264_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_189_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_349_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16476_ _15168_/X _22396_/Q _16480_/S vssd1 vssd1 vccd1 vccd1 _16477_/A sky130_fd_sc_hd__mux2_1
X_13688_ _13688_/A vssd1 vssd1 vccd1 vccd1 _14231_/A sky130_fd_sc_hd__clkbuf_2
X_18215_ _22850_/Q _18202_/X _18214_/X _18206_/X vssd1 vssd1 vccd1 vccd1 _22898_/D
+ sky130_fd_sc_hd__o211a_1
X_15427_ _15480_/A vssd1 vssd1 vccd1 vccd1 _15564_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_129_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12639_ _22470_/Q _22630_/Q _12755_/A vssd1 vssd1 vccd1 vccd1 _12639_/X sky130_fd_sc_hd__mux2_1
XPHY_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19195_ _19194_/X _23278_/Q _19195_/S vssd1 vssd1 vccd1 vccd1 _19196_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_352_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_318_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18146_ _14121_/D _22878_/Q _18158_/S vssd1 vssd1 vccd1 vccd1 _18147_/B sky130_fd_sc_hd__mux2_1
X_15358_ _23696_/Q _14494_/S _15357_/X vssd1 vssd1 vccd1 vccd1 _15358_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_156_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_356_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_306_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14309_ _13029_/B _12611_/B _14326_/S vssd1 vssd1 vccd1 vccd1 _14309_/X sky130_fd_sc_hd__mux2_1
XFILLER_305_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18077_ hold5/A _18067_/X _18068_/X _22996_/Q _18069_/X vssd1 vssd1 vccd1 vccd1 _18077_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15289_ _14720_/Y _15181_/X _15183_/X _15288_/Y vssd1 vssd1 vccd1 vccd1 _21231_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17028_ _17028_/A vssd1 vssd1 vccd1 vccd1 _17028_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_301_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18979_ _16860_/X _23187_/Q _18979_/S vssd1 vssd1 vccd1 vccd1 _18980_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21990_ _23803_/Q _21746_/X _21989_/Y _21395_/X vssd1 vssd1 vccd1 vccd1 _21990_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_273_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20941_ _21791_/A _20936_/X _20672_/B _20940_/X vssd1 vssd1 vccd1 vccd1 _20941_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_282_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23660_ _23700_/CLK _23660_/D vssd1 vssd1 vccd1 vccd1 _23660_/Q sky130_fd_sc_hd__dfxtp_1
X_20872_ _20742_/B _20864_/X _20865_/X _23775_/Q vssd1 vssd1 vccd1 vccd1 _20873_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22611_ _23552_/CLK _22611_/D vssd1 vssd1 vccd1 vccd1 _22611_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23591_ _23592_/CLK _23591_/D vssd1 vssd1 vccd1 vccd1 _23591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_329_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22542_ _23546_/CLK _22542_/D vssd1 vssd1 vccd1 vccd1 _22542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_356_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_355_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22473_ _23448_/CLK _22473_/D vssd1 vssd1 vccd1 vccd1 _22473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_309_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21424_ _21452_/A _21452_/B vssd1 vssd1 vccd1 vccd1 _21543_/B sky130_fd_sc_hd__xor2_1
XFILLER_355_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21355_ _21351_/B _21353_/Y _22091_/B vssd1 vssd1 vccd1 vccd1 _21355_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_297_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_49_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23537_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20306_ _20396_/A _20306_/B vssd1 vssd1 vccd1 vccd1 _20306_/X sky130_fd_sc_hd__or2_1
XFILLER_150_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21286_ _21379_/A _21289_/B vssd1 vssd1 vccd1 vccd1 _21287_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23025_ _23504_/CLK _23025_/D vssd1 vssd1 vccd1 vccd1 _23025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20237_ _20196_/X _20235_/X _20236_/Y _21576_/A _20200_/X vssd1 vssd1 vccd1 vccd1
+ _20615_/A sky130_fd_sc_hd__a32o_4
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20168_ _20168_/A vssd1 vssd1 vccd1 vccd1 _20169_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20099_ _20112_/C vssd1 vssd1 vccd1 vccd1 _20106_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12990_ _13051_/A _11398_/A _11403_/A _12989_/Y vssd1 vssd1 vccd1 vccd1 _13026_/A
+ sky130_fd_sc_hd__a22o_4
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23927_ _23936_/CLK _23927_/D vssd1 vssd1 vccd1 vccd1 _23927_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11941_ _13518_/B vssd1 vssd1 vccd1 vccd1 _13380_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_218_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _14359_/X _14349_/X _14660_/S vssd1 vssd1 vccd1 vccd1 _14660_/X sky130_fd_sc_hd__mux2_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _12489_/A vssd1 vssd1 vccd1 vccd1 _12387_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23858_ _23862_/CLK _23858_/D vssd1 vssd1 vccd1 vccd1 _23858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_260_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13611_ _13611_/A _13611_/B vssd1 vssd1 vccd1 vccd1 _13611_/X sky130_fd_sc_hd__or2_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22809_ _23693_/CLK _22809_/D vssd1 vssd1 vccd1 vccd1 _22809_/Q sky130_fd_sc_hd__dfxtp_2
X_14591_ _15440_/A vssd1 vssd1 vccd1 vccd1 _14592_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23789_ _23861_/CLK _23789_/D vssd1 vssd1 vccd1 vccd1 _23789_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_198_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16330_ _16330_/A vssd1 vssd1 vccd1 vccd1 _22332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13542_ _13542_/A _14274_/B vssd1 vssd1 vccd1 vccd1 _13542_/Y sky130_fd_sc_hd__nand2_1
XFILLER_347_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16261_ _16261_/A vssd1 vssd1 vccd1 vccd1 _22309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13473_ _14199_/A _13473_/B vssd1 vssd1 vccd1 vccd1 _13884_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18000_ _18029_/A vssd1 vssd1 vccd1 vccd1 _18000_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_200_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15212_ _16170_/B vssd1 vssd1 vccd1 vccd1 _15905_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_334_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12424_ _22295_/Q _23431_/Q _12424_/S vssd1 vssd1 vccd1 vccd1 _12425_/B sky130_fd_sc_hd__mux2_1
XFILLER_139_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16192_ _16005_/X _16190_/Y _16191_/Y _15574_/A vssd1 vssd1 vccd1 vccd1 _16192_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_355_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_327_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15143_ _23724_/Q _23854_/Q _15354_/S vssd1 vssd1 vccd1 vccd1 _15143_/X sky130_fd_sc_hd__mux2_1
XFILLER_354_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12355_ _22360_/Q _22392_/Q _22681_/Q _23048_/Q _11413_/A _11702_/A vssd1 vssd1 vccd1
+ vccd1 _12355_/X sky130_fd_sc_hd__mux4_2
XFILLER_315_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11306_ _11637_/A vssd1 vssd1 vccd1 vccd1 _12843_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_181_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19951_ _19977_/B _19953_/C _19950_/Y vssd1 vssd1 vccd1 vccd1 _23599_/D sky130_fd_sc_hd__o21a_1
X_15074_ _14592_/A _15065_/X _15073_/X _14748_/A vssd1 vssd1 vccd1 vccd1 _15074_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_153_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12286_ _12606_/A _12605_/A vssd1 vssd1 vccd1 vccd1 _12287_/B sky130_fd_sc_hd__nor2_1
XFILLER_316_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_302_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18902_ _18902_/A vssd1 vssd1 vccd1 vccd1 _23152_/D sky130_fd_sc_hd__clkbuf_1
X_11237_ _15826_/A _11226_/X _11236_/X vssd1 vssd1 vccd1 vccd1 _11237_/Y sky130_fd_sc_hd__o21ai_1
X_14025_ _13748_/B _14049_/A vssd1 vssd1 vccd1 vccd1 _14025_/X sky130_fd_sc_hd__and2b_1
X_19882_ _19882_/A vssd1 vssd1 vccd1 vccd1 _23573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_353_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18833_ _18833_/A vssd1 vssd1 vccd1 vccd1 _18833_/X sky130_fd_sc_hd__buf_2
XFILLER_296_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11168_ _11207_/A vssd1 vssd1 vccd1 vccd1 _11169_/A sky130_fd_sc_hd__buf_6
XTAP_6260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_295_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18764_ _18764_/A vssd1 vssd1 vccd1 vccd1 _23106_/D sky130_fd_sc_hd__clkbuf_1
X_15976_ _15976_/A vssd1 vssd1 vccd1 vccd1 _16125_/S sky130_fd_sc_hd__buf_6
XTAP_5570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11099_ _11099_/A vssd1 vssd1 vccd1 vccd1 _14521_/A sky130_fd_sc_hd__buf_8
XFILLER_110_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17715_ _22737_/Q _17623_/X _17715_/S vssd1 vssd1 vccd1 vccd1 _17716_/A sky130_fd_sc_hd__mux2_1
X_14927_ _15735_/A vssd1 vssd1 vccd1 vccd1 _16177_/S sky130_fd_sc_hd__clkbuf_2
X_18695_ _23076_/Q _17645_/X _18695_/S vssd1 vssd1 vccd1 vccd1 _18696_/A sky130_fd_sc_hd__mux2_1
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17646_ _22709_/Q _17645_/X _17646_/S vssd1 vssd1 vccd1 vccd1 _17647_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14858_ _14854_/S _14293_/X _14376_/X vssd1 vssd1 vccd1 vccd1 _14858_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13809_ _12940_/B _13808_/X _13781_/X vssd1 vssd1 vccd1 vccd1 _13809_/X sky130_fd_sc_hd__a21o_1
XFILLER_90_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17577_ _17577_/A vssd1 vssd1 vccd1 vccd1 _22687_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14789_ _14784_/Y _14787_/X _15088_/S vssd1 vssd1 vccd1 vccd1 _14789_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19316_ _19233_/X _23322_/Q _19322_/S vssd1 vssd1 vccd1 vccd1 _19317_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16528_ _16197_/X _22420_/Q _16528_/S vssd1 vssd1 vccd1 vccd1 _16529_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_338_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19247_ _19245_/X _23294_/Q _19259_/S vssd1 vssd1 vccd1 vccd1 _19248_/A sky130_fd_sc_hd__mux2_1
XFILLER_337_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16459_ _16515_/A vssd1 vssd1 vccd1 vccd1 _16528_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_192_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_337_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19178_ _19178_/A vssd1 vssd1 vccd1 vccd1 _19178_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_192_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_334_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_352_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18129_ _14119_/B _22880_/Q _18187_/A vssd1 vssd1 vccd1 vccd1 _18129_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21140_ _21158_/A vssd1 vssd1 vccd1 vccd1 _21140_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_333_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21071_ _20759_/A _21008_/A _21070_/X _21061_/X vssd1 vssd1 vccd1 vccd1 _23843_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_287_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20022_ _20041_/A _20022_/B _20034_/C vssd1 vssd1 vccd1 vccd1 _23618_/D sky130_fd_sc_hd__nor3_1
XFILLER_286_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_301_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_286_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_167_wb_clk_i _23917_/CLK vssd1 vssd1 vccd1 vccd1 _23871_/CLK sky130_fd_sc_hd__clkbuf_16
X_21973_ _23834_/Q _21972_/Y _21973_/S vssd1 vssd1 vccd1 vccd1 _21973_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23712_ _23714_/CLK _23712_/D vssd1 vssd1 vccd1 vccd1 _23712_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20924_ _23790_/Q _20911_/X _20923_/X _20920_/X vssd1 vssd1 vccd1 vccd1 _23790_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23643_ _23643_/CLK _23643_/D vssd1 vssd1 vccd1 vccd1 _23643_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20855_ _20861_/A _20855_/B vssd1 vssd1 vccd1 vccd1 _20856_/A sky130_fd_sc_hd__and2_1
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_288_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_356_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23574_ _23574_/CLK _23574_/D vssd1 vssd1 vccd1 vccd1 _23574_/Q sky130_fd_sc_hd__dfxtp_1
X_20786_ _23752_/Q _20786_/B vssd1 vssd1 vccd1 vccd1 _20786_/X sky130_fd_sc_hd__or2_1
XFILLER_288_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22525_ _23561_/CLK _22525_/D vssd1 vssd1 vccd1 vccd1 _22525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_356_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_356_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22456_ _22779_/CLK _22456_/D vssd1 vssd1 vccd1 vccd1 _22456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_339_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21407_ _21677_/A vssd1 vssd1 vccd1 vccd1 _21767_/A sky130_fd_sc_hd__buf_2
XFILLER_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22387_ _23491_/CLK _22387_/D vssd1 vssd1 vccd1 vccd1 _22387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12140_ _23473_/Q _23569_/Q _22533_/Q _22337_/Q _11745_/X _12014_/A vssd1 vssd1 vccd1
+ vccd1 _12141_/B sky130_fd_sc_hd__mux4_1
XFILLER_340_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_325_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21338_ _11084_/A _21518_/A _21382_/A vssd1 vssd1 vccd1 vccd1 _21441_/A sky130_fd_sc_hd__a21o_1
XFILLER_194_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12071_ _12071_/A _12071_/B vssd1 vssd1 vccd1 vccd1 _12071_/Y sky130_fd_sc_hd__nand2_1
X_21269_ _21269_/A _21274_/B vssd1 vssd1 vccd1 vccd1 _21269_/Y sky130_fd_sc_hd__nand2_1
XFILLER_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23008_ _23008_/CLK _23008_/D vssd1 vssd1 vccd1 vccd1 _23008_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_277_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_293_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ _15830_/A _15830_/B vssd1 vssd1 vccd1 vccd1 _15830_/Y sky130_fd_sc_hd__nand2_2
XFILLER_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_293_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _23833_/Q _14907_/A _15757_/X _15760_/X _14923_/A vssd1 vssd1 vccd1 vccd1
+ _15761_/X sky130_fd_sc_hd__a221o_1
X_12973_ _23419_/Q _23035_/Q _23387_/Q _23355_/Q _12921_/S _12749_/X vssd1 vssd1 vccd1
+ vccd1 _12973_/X sky130_fd_sc_hd__mux4_2
XFILLER_292_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_346_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17500_ _17500_/A vssd1 vssd1 vccd1 vccd1 _22657_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _23913_/Q vssd1 vssd1 vccd1 vccd1 _14713_/A sky130_fd_sc_hd__buf_6
X_18480_ _18480_/A vssd1 vssd1 vccd1 vccd1 _18480_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _11284_/A _11914_/X _11916_/X _11923_/X vssd1 vssd1 vccd1 vccd1 _11924_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_46_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _23703_/Q _15210_/X _15691_/X vssd1 vssd1 vccd1 vccd1 _15692_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_307_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17431_ _17431_/A vssd1 vssd1 vccd1 vccd1 _22627_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _14270_/X _14275_/X _14646_/S vssd1 vssd1 vccd1 vccd1 _14643_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _11834_/A _11854_/X _11230_/A vssd1 vssd1 vccd1 vccd1 _11855_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17362_ _17362_/A vssd1 vssd1 vccd1 vccd1 _22601_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14574_ input159/X input124/X _14967_/S vssd1 vssd1 vccd1 vccd1 _14574_/X sky130_fd_sc_hd__mux2_8
XFILLER_158_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11786_ _23407_/Q _23023_/Q _23375_/Q _23343_/Q _12070_/S _11163_/A vssd1 vssd1 vccd1
+ vccd1 _11786_/X sky130_fd_sc_hd__mux4_1
XFILLER_213_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19101_ _19101_/A vssd1 vssd1 vccd1 vccd1 _23240_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16313_ _16381_/S vssd1 vssd1 vccd1 vccd1 _16322_/S sky130_fd_sc_hd__buf_6
XFILLER_319_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13525_ _13525_/A _13525_/B vssd1 vssd1 vccd1 vccd1 _13526_/A sky130_fd_sc_hd__nor2_1
X_17293_ _17245_/X _17292_/X _17262_/X _17283_/X vssd1 vssd1 vccd1 vccd1 _17293_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_348_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19032_ _16831_/X _23210_/Q _19040_/S vssd1 vssd1 vccd1 vccd1 _19033_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16244_ _22304_/Q _16243_/X _16253_/S vssd1 vssd1 vccd1 vccd1 _16245_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_348_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13456_ _16679_/A _22519_/Q vssd1 vssd1 vccd1 vccd1 _13457_/A sky130_fd_sc_hd__nor2_1
XFILLER_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_328_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12407_ _22359_/Q _22391_/Q _22680_/Q _23047_/Q _11920_/X _11652_/A vssd1 vssd1 vccd1
+ vccd1 _12407_/X sky130_fd_sc_hd__mux4_2
X_16175_ _23716_/Q _15592_/A _16174_/X vssd1 vssd1 vccd1 vccd1 _16175_/X sky130_fd_sc_hd__o21a_4
X_13387_ _13387_/A _13387_/B _15580_/A _13387_/D vssd1 vssd1 vccd1 vccd1 _13395_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15126_ _20186_/A _13928_/A _15125_/X vssd1 vssd1 vccd1 vccd1 _15139_/A sky130_fd_sc_hd__a21oi_1
XFILLER_343_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12338_ _23916_/Q _12415_/S vssd1 vssd1 vccd1 vccd1 _12338_/Y sky130_fd_sc_hd__nor2_1
XFILLER_303_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_287_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19934_ _23595_/Q _19934_/B _19934_/C vssd1 vssd1 vccd1 vccd1 _19935_/C sky130_fd_sc_hd__and3_1
XFILLER_303_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15057_ input147/X input112/X _15057_/S vssd1 vssd1 vccd1 vccd1 _15057_/X sky130_fd_sc_hd__mux2_8
XFILLER_141_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_330_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12269_ _12269_/A vssd1 vssd1 vccd1 vccd1 _12269_/X sky130_fd_sc_hd__buf_4
XFILLER_330_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_287_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_296_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14008_ _14072_/C vssd1 vssd1 vccd1 vccd1 _14083_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19865_ _16236_/X _23566_/Q _19865_/S vssd1 vssd1 vccd1 vccd1 _19866_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_296_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_311_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18816_ _18816_/A vssd1 vssd1 vccd1 vccd1 _23122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19796_ _23535_/Q _19197_/A _19804_/S vssd1 vssd1 vccd1 vccd1 _19797_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18747_ _18747_/A vssd1 vssd1 vccd1 vccd1 _23098_/D sky130_fd_sc_hd__clkbuf_1
X_15959_ _23710_/Q _15592_/X _15958_/X vssd1 vssd1 vccd1 vccd1 _15959_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_237_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18678_ _23068_/Q _17620_/X _18680_/S vssd1 vssd1 vccd1 vccd1 _18679_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17629_ _17629_/A vssd1 vssd1 vccd1 vccd1 _22703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20640_ _20895_/A vssd1 vssd1 vccd1 vccd1 _20669_/B sky130_fd_sc_hd__buf_4
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20571_ _20571_/A _20936_/A vssd1 vssd1 vccd1 vccd1 _20577_/B sky130_fd_sc_hd__nor2_2
XFILLER_165_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22310_ _22695_/CLK _22310_/D vssd1 vssd1 vccd1 vccd1 _22310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23290_ _23548_/CLK _23290_/D vssd1 vssd1 vccd1 vccd1 _23290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_338_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_319_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22241_ _22025_/A _22242_/C _23844_/Q vssd1 vssd1 vccd1 vccd1 _22241_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_322_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22172_ _21712_/S _22170_/Y _22171_/Y _21767_/A vssd1 vssd1 vccd1 vccd1 _22172_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_127_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21123_ _21161_/A vssd1 vssd1 vccd1 vccd1 _21123_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_322_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21054_ _21165_/A _21064_/B vssd1 vssd1 vccd1 vccd1 _21054_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20005_ _23608_/Q _23607_/Q _20005_/C _20005_/D vssd1 vssd1 vccd1 vccd1 _20007_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_259_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_290_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_290_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_290_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21956_ _21981_/A _21956_/B vssd1 vssd1 vccd1 vccd1 _21956_/Y sky130_fd_sc_hd__nand2_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_299_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20907_ _23784_/Q _20893_/X _20905_/X _20906_/X vssd1 vssd1 vccd1 vccd1 _23784_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21887_ _21888_/A _21888_/B vssd1 vssd1 vccd1 vccd1 _21889_/A sky130_fd_sc_hd__nand2_1
XFILLER_203_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23626_ _23634_/CLK _23626_/D vssd1 vssd1 vccd1 vccd1 _23626_/Q sky130_fd_sc_hd__dfxtp_1
X_11640_ _23478_/Q _23574_/Q _22538_/Q _22342_/Q _12843_/A _12777_/A vssd1 vssd1 vccd1
+ vccd1 _11641_/B sky130_fd_sc_hd__mux4_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20838_ _20838_/A vssd1 vssd1 vccd1 vccd1 _23765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_357_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11571_ _12457_/S vssd1 vssd1 vccd1 vccd1 _12556_/A sky130_fd_sc_hd__buf_4
X_23557_ _23896_/CLK _23557_/D vssd1 vssd1 vccd1 vccd1 _23557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_357_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20769_ _23748_/Q _20628_/A _20768_/X _20763_/X vssd1 vssd1 vccd1 vccd1 _23748_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_64_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23543_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13310_ _13318_/A _13403_/B _13554_/A _13555_/A vssd1 vssd1 vccd1 vccd1 _13310_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_122_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22508_ _23693_/CLK _22508_/D vssd1 vssd1 vccd1 vccd1 _22508_/Q sky130_fd_sc_hd__dfxtp_4
X_14290_ _14290_/A vssd1 vssd1 vccd1 vccd1 _14369_/A sky130_fd_sc_hd__clkbuf_2
X_23488_ _23552_/CLK _23488_/D vssd1 vssd1 vccd1 vccd1 _23488_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_155_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13241_ _13241_/A vssd1 vssd1 vccd1 vccd1 _13242_/B sky130_fd_sc_hd__inv_2
X_22439_ _23510_/CLK _22439_/D vssd1 vssd1 vccd1 vccd1 _22439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13172_ _13229_/A _13172_/B vssd1 vssd1 vccd1 vccd1 _13172_/X sky130_fd_sc_hd__or2_1
XFILLER_182_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ _12117_/A _12118_/X _12122_/X _11131_/A vssd1 vssd1 vccd1 vccd1 _12123_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_151_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17980_ _22837_/Q _17965_/X _17978_/X _17979_/X vssd1 vssd1 vccd1 vccd1 _22837_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12054_ _11141_/A _12053_/X _11598_/X vssd1 vssd1 vccd1 vccd1 _12054_/Y sky130_fd_sc_hd__o21ai_1
X_16931_ _16950_/B vssd1 vssd1 vccd1 vccd1 _16932_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_313_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16862_ _16862_/A vssd1 vssd1 vccd1 vccd1 _22535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19650_ _19650_/A vssd1 vssd1 vccd1 vccd1 _23470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_277_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18601_ _18601_/A vssd1 vssd1 vccd1 vccd1 _23033_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_293_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15813_ _22935_/Q _14509_/A _14513_/A _22967_/Q vssd1 vssd1 vccd1 vccd1 _15813_/X
+ sky130_fd_sc_hd__o22a_1
X_19581_ _19581_/A vssd1 vssd1 vccd1 vccd1 _23439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_265_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16793_ _16793_/A vssd1 vssd1 vccd1 vccd1 _22514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_293_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_292_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18532_ _23008_/Q _18534_/B vssd1 vssd1 vccd1 vccd1 _18532_/Y sky130_fd_sc_hd__nand2_1
X_15744_ _21898_/A _15478_/X _15743_/X vssd1 vssd1 vccd1 vccd1 _15744_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12956_ _23321_/Q _23289_/Q _23257_/Q _23545_/Q _12716_/X _12717_/X vssd1 vssd1 vccd1
+ vccd1 _12956_/X sky130_fd_sc_hd__mux4_2
XFILLER_252_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _18476_/A vssd1 vssd1 vccd1 vccd1 _18463_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11907_ _11890_/A _11906_/X _11706_/X vssd1 vssd1 vccd1 vccd1 _11907_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _15865_/A _15675_/B vssd1 vssd1 vccd1 vccd1 _15675_/Y sky130_fd_sc_hd__nand2_2
XFILLER_18_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _23482_/Q _23578_/Q _22542_/Q _22346_/Q _12755_/X _12756_/X vssd1 vssd1 vccd1
+ vccd1 _12887_/X sky130_fd_sc_hd__mux4_1
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _17414_/A vssd1 vssd1 vccd1 vccd1 _22619_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _14291_/X _14381_/B _14850_/S vssd1 vssd1 vccd1 vccd1 _14626_/X sky130_fd_sc_hd__mux2_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18394_ _22959_/Q _18394_/B vssd1 vssd1 vccd1 vccd1 _18400_/C sky130_fd_sc_hd__and2_1
X_11838_ _22302_/Q _23438_/Q _12554_/S vssd1 vssd1 vccd1 vccd1 _11839_/B sky130_fd_sc_hd__mux2_1
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_348_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _22594_/Q input211/X _17347_/S vssd1 vssd1 vccd1 vccd1 _17346_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_320_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14557_ _14557_/A _14557_/B vssd1 vssd1 vccd1 vccd1 _16457_/C sky130_fd_sc_hd__nand2_1
XFILLER_147_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11769_ _11853_/A vssd1 vssd1 vccd1 vccd1 _11905_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_347_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13508_ _14313_/A _13508_/B vssd1 vssd1 vccd1 vccd1 _13508_/Y sky130_fd_sc_hd__nor2_2
X_17276_ _17276_/A vssd1 vssd1 vccd1 vccd1 _17314_/S sky130_fd_sc_hd__clkbuf_4
X_14488_ _23813_/Q _14464_/X _14472_/X _14478_/X _14487_/X vssd1 vssd1 vccd1 vccd1
+ _14488_/X sky130_fd_sc_hd__a221o_1
XFILLER_347_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19015_ _19015_/A vssd1 vssd1 vccd1 vccd1 _23203_/D sky130_fd_sc_hd__clkbuf_1
X_16227_ _18792_/A vssd1 vssd1 vccd1 vccd1 _16227_/X sky130_fd_sc_hd__clkbuf_2
X_13439_ _13439_/A vssd1 vssd1 vccd1 vccd1 _14866_/A sky130_fd_sc_hd__buf_4
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16158_ _23008_/Q _16944_/A _16085_/X input238/X vssd1 vssd1 vccd1 vccd1 _22224_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_344_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_343_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15109_ _15109_/A _15109_/B vssd1 vssd1 vccd1 vccd1 _15176_/C sky130_fd_sc_hd__nor2_1
XFILLER_303_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16089_ _19255_/A vssd1 vssd1 vccd1 vccd1 _16089_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19917_ _19915_/X _19916_/X _18423_/X vssd1 vssd1 vccd1 vccd1 _19917_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_114_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19848_ _16211_/X _23558_/Q _19854_/S vssd1 vssd1 vccd1 vccd1 _19849_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_288_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19779_ _19779_/A vssd1 vssd1 vccd1 vccd1 _23527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21810_ _21876_/A _21810_/B vssd1 vssd1 vccd1 vccd1 _21934_/A sky130_fd_sc_hd__nor2_1
XFILLER_260_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22790_ _23459_/CLK _22790_/D vssd1 vssd1 vccd1 vccd1 _22790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21741_ _21741_/A _22032_/B vssd1 vssd1 vccd1 vccd1 _21741_/Y sky130_fd_sc_hd__nor2_1
XFILLER_280_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21672_ _21673_/A _21676_/A vssd1 vssd1 vccd1 vccd1 _21674_/A sky130_fd_sc_hd__and2_1
XFILLER_339_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23411_ _23507_/CLK _23411_/D vssd1 vssd1 vccd1 vccd1 _23411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20623_ _20623_/A _20631_/B vssd1 vssd1 vccd1 vccd1 _20626_/B sky130_fd_sc_hd__nor2_4
XFILLER_138_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_327_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20554_ _21300_/B _20632_/A _20553_/X vssd1 vssd1 vccd1 vccd1 _20558_/B sky130_fd_sc_hd__o21a_1
X_23342_ _23534_/CLK _23342_/D vssd1 vssd1 vccd1 vccd1 _23342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_295_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_354_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_354_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_353_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_353_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20485_ _23713_/Q _20487_/B vssd1 vssd1 vccd1 vccd1 _20485_/X sky130_fd_sc_hd__or2_1
X_23273_ _23529_/CLK _23273_/D vssd1 vssd1 vccd1 vccd1 _23273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_313_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_307_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22224_ _22224_/A _22224_/B vssd1 vssd1 vccd1 vccd1 _22224_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_336_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22155_ _22155_/A _22155_/B _22155_/C _22155_/D vssd1 vssd1 vccd1 vccd1 _22155_/X
+ sky130_fd_sc_hd__and4_1
XTAP_6804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput460 _23885_/Q vssd1 vssd1 vccd1 vccd1 probe_opcode[6] sky130_fd_sc_hd__buf_2
XTAP_6826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21106_ _21108_/A _21106_/B vssd1 vssd1 vccd1 vccd1 _23850_/D sky130_fd_sc_hd__nor2_1
Xoutput471 _23930_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[19] sky130_fd_sc_hd__buf_2
XTAP_6837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput482 _23940_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[29] sky130_fd_sc_hd__buf_2
XTAP_6848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput493 _23945_/Q vssd1 vssd1 vccd1 vccd1 probe_state[0] sky130_fd_sc_hd__buf_2
X_22086_ _22116_/A _22116_/B vssd1 vssd1 vccd1 vccd1 _22086_/X sky130_fd_sc_hd__and2_1
XTAP_6859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_111_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _22893_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21037_ _21163_/A vssd1 vssd1 vccd1 vccd1 _21037_/X sky130_fd_sc_hd__buf_2
XFILLER_304_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12810_ _13532_/D vssd1 vssd1 vccd1 vccd1 _13629_/A sky130_fd_sc_hd__inv_2
XFILLER_170_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13790_ _13829_/B vssd1 vssd1 vccd1 vccd1 _13790_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_320_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22988_ _23009_/CLK _22988_/D vssd1 vssd1 vccd1 vccd1 _22988_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_216_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12741_ _12742_/A _12807_/A vssd1 vssd1 vccd1 vccd1 _12741_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21939_ _21812_/B _21935_/Y _22040_/A vssd1 vssd1 vccd1 vccd1 _21940_/B sky130_fd_sc_hd__o21bai_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15460_ _15460_/A _15460_/B vssd1 vssd1 vccd1 vccd1 _15460_/Y sky130_fd_sc_hd__nand2_1
X_12672_ _12672_/A vssd1 vssd1 vccd1 vccd1 _13195_/A sky130_fd_sc_hd__buf_2
XFILLER_230_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14411_ _14179_/A _14551_/A _14433_/S vssd1 vssd1 vccd1 vccd1 _14416_/B sky130_fd_sc_hd__mux2_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23609_ _23652_/CLK _23609_/D vssd1 vssd1 vccd1 vccd1 _23609_/Q sky130_fd_sc_hd__dfxtp_1
X_11623_ _11961_/A _11623_/B vssd1 vssd1 vccd1 vccd1 _11623_/X sky130_fd_sc_hd__or2_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15391_ _15391_/A _16180_/B vssd1 vssd1 vccd1 vccd1 _15391_/Y sky130_fd_sc_hd__nor2_1
XFILLER_318_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17130_ _22566_/Q _17091_/X _17083_/X _17129_/X vssd1 vssd1 vccd1 vccd1 _22566_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_169_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_357_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14342_ _12606_/B _13240_/A _15171_/A vssd1 vssd1 vccd1 vccd1 _14342_/X sky130_fd_sc_hd__mux2_1
XFILLER_329_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11554_ _16114_/A _20387_/A _13296_/B vssd1 vssd1 vccd1 vccd1 _11555_/A sky130_fd_sc_hd__mux2_2
XFILLER_318_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_317_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17061_ _17230_/A vssd1 vssd1 vccd1 vccd1 _17061_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_184_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14273_ _14288_/A vssd1 vssd1 vccd1 vccd1 _14326_/S sky130_fd_sc_hd__buf_2
X_11485_ _13295_/A _11485_/B _11485_/C vssd1 vssd1 vccd1 vccd1 _20394_/A sky130_fd_sc_hd__nor3_4
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16012_ _18856_/A vssd1 vssd1 vccd1 vccd1 _19249_/A sky130_fd_sc_hd__clkbuf_2
X_13224_ _23325_/Q _23293_/Q _23261_/Q _23549_/Q _11517_/A _11527_/A vssd1 vssd1 vccd1
+ vccd1 _13225_/B sky130_fd_sc_hd__mux4_2
XFILLER_195_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_326_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_325_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13155_ _23422_/Q _23038_/Q _23390_/Q _23358_/Q _11431_/A _13037_/A vssd1 vssd1 vccd1
+ vccd1 _13155_/X sky130_fd_sc_hd__mux4_1
XFILLER_313_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_298_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_345_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12106_ _22467_/Q _22627_/Q _22306_/Q _23442_/Q _12094_/X _11457_/B vssd1 vssd1 vccd1
+ vccd1 _12106_/X sky130_fd_sc_hd__mux4_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17963_ _18029_/A vssd1 vssd1 vccd1 vccd1 _17963_/X sky130_fd_sc_hd__clkbuf_2
X_13086_ _22803_/Q _22771_/Q _22672_/Q _22739_/Q _11205_/A _13085_/X vssd1 vssd1 vccd1
+ vccd1 _13087_/B sky130_fd_sc_hd__mux4_2
XFILLER_239_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_340_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19702_ _19163_/X _23493_/Q _19710_/S vssd1 vssd1 vccd1 vccd1 _19703_/A sky130_fd_sc_hd__mux2_1
XFILLER_300_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12037_ _12634_/A _12037_/B _12037_/C vssd1 vssd1 vccd1 vccd1 _12037_/Y sky130_fd_sc_hd__nor3_4
X_16914_ _19264_/A vssd1 vssd1 vccd1 vccd1 _16914_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_238_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17894_ _18097_/A vssd1 vssd1 vccd1 vccd1 _17894_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_266_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_293_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19633_ _19633_/A vssd1 vssd1 vccd1 vccd1 _23462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16845_ _16844_/X _22530_/Q _16845_/S vssd1 vssd1 vccd1 vccd1 _16846_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16776_ _22510_/Q _16765_/X _16766_/X input25/X vssd1 vssd1 vccd1 vccd1 _16777_/B
+ sky130_fd_sc_hd__o22a_1
X_19564_ _23432_/Q _19175_/A _19566_/S vssd1 vssd1 vccd1 vccd1 _19565_/A sky130_fd_sc_hd__mux2_1
X_13988_ _13990_/A _14082_/A vssd1 vssd1 vccd1 vccd1 _13988_/Y sky130_fd_sc_hd__nor2_8
XFILLER_19_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18515_ _23001_/Q _18518_/B vssd1 vssd1 vccd1 vccd1 _18515_/Y sky130_fd_sc_hd__nand2_1
X_15727_ _23608_/Q _14731_/A _14733_/A _23640_/Q vssd1 vssd1 vccd1 vccd1 _15727_/X
+ sky130_fd_sc_hd__o22a_4
X_12939_ _11219_/A _12929_/X _12938_/X _11124_/A vssd1 vssd1 vccd1 vccd1 _12940_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19495_ _19495_/A vssd1 vssd1 vccd1 vccd1 _23401_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18446_ _22976_/Q _18444_/B _18445_/Y vssd1 vssd1 vccd1 vccd1 _22976_/D sky130_fd_sc_hd__o21a_1
XFILLER_34_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15658_ _14822_/A _15634_/X _15657_/Y _14882_/A vssd1 vssd1 vccd1 vccd1 _15658_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14609_ _14609_/A _20409_/A vssd1 vssd1 vccd1 vccd1 _14610_/A sky130_fd_sc_hd__nor2_2
X_18377_ _22953_/Q _18377_/B vssd1 vssd1 vccd1 vccd1 _18384_/C sky130_fd_sc_hd__and2_1
X_15589_ _15589_/A vssd1 vssd1 vccd1 vccd1 _15589_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17328_ _22586_/Q _17324_/Y _17335_/S vssd1 vssd1 vccd1 vccd1 _22586_/D sky130_fd_sc_hd__a21o_1
XFILLER_239_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_336_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17259_ _23486_/Q _17230_/X _17231_/X _17181_/X _17258_/Y vssd1 vssd1 vccd1 vccd1
+ _17259_/X sky130_fd_sc_hd__a32o_1
XFILLER_146_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_335_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_351_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20270_ _20323_/A _21025_/A vssd1 vssd1 vccd1 vccd1 _20270_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_303_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_332_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22911_ _22956_/CLK _22911_/D vssd1 vssd1 vccd1 vccd1 _22911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23891_ _23893_/CLK _23891_/D vssd1 vssd1 vccd1 vccd1 _23891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22842_ _22893_/CLK _22842_/D vssd1 vssd1 vccd1 vccd1 _22842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22773_ _23073_/CLK _22773_/D vssd1 vssd1 vccd1 vccd1 _22773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_262_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21724_ _21724_/A _21724_/B vssd1 vssd1 vccd1 vccd1 _21801_/B sky130_fd_sc_hd__nor2_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21655_ _21689_/C _21694_/B vssd1 vssd1 vccd1 vccd1 _21658_/A sky130_fd_sc_hd__nor2_1
XFILLER_235_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_303_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20606_ _13440_/A _20564_/X _20598_/X vssd1 vssd1 vccd1 vccd1 _20606_/X sky130_fd_sc_hd__a21o_1
XFILLER_296_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21586_ _21564_/A _21566_/B _21563_/Y vssd1 vssd1 vccd1 vccd1 _21587_/B sky130_fd_sc_hd__o21ai_2
XFILLER_296_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23325_ _23549_/CLK _23325_/D vssd1 vssd1 vccd1 vccd1 _23325_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_opt_4_1_wb_clk_i clkbuf_opt_4_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_4_1_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_20537_ _20544_/A vssd1 vssd1 vccd1 vccd1 _21308_/B sky130_fd_sc_hd__inv_2
XFILLER_327_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23256_ _23354_/CLK _23256_/D vssd1 vssd1 vccd1 vccd1 _23256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_308_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11270_ _23942_/Q vssd1 vssd1 vccd1 vccd1 _11270_/Y sky130_fd_sc_hd__clkinv_2
X_20468_ _23706_/Q _20468_/B vssd1 vssd1 vccd1 vccd1 _20468_/X sky130_fd_sc_hd__or2_1
XTAP_7302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_7313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_307_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22207_ _22207_/A _22207_/B vssd1 vssd1 vccd1 vccd1 _22207_/Y sky130_fd_sc_hd__xnor2_4
XTAP_7324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23187_ _23507_/CLK _23187_/D vssd1 vssd1 vccd1 vccd1 _23187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20399_ _20213_/A _20759_/A _20398_/X _20392_/X vssd1 vssd1 vccd1 vccd1 _23683_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_7346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22138_ _22151_/A _22242_/B _22137_/Y _21634_/A vssd1 vssd1 vccd1 vccd1 _22146_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_7379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput290 _14094_/X vssd1 vssd1 vccd1 vccd1 addr0[5] sky130_fd_sc_hd__buf_2
XTAP_6656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14960_ input136/X input151/X _15052_/S vssd1 vssd1 vccd1 vccd1 _14960_/X sky130_fd_sc_hd__mux2_8
XTAP_6689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22069_ _21379_/X _22054_/X _22061_/Y _22068_/X _21479_/A vssd1 vssd1 vccd1 vccd1
+ _22071_/A sky130_fd_sc_hd__o2111a_1
XFILLER_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13911_ _13503_/Y _14794_/A _13902_/B _13508_/Y vssd1 vssd1 vccd1 vccd1 _13911_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_5977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14891_ _12393_/Y _14530_/X _14889_/X _21406_/A _14703_/X vssd1 vssd1 vccd1 vccd1
+ _18782_/A sky130_fd_sc_hd__a32o_4
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16630_ _16630_/A vssd1 vssd1 vccd1 vccd1 _22463_/D sky130_fd_sc_hd__clkbuf_1
X_13842_ _13842_/A _13864_/B vssd1 vssd1 vccd1 vccd1 _13842_/Y sky130_fd_sc_hd__nor2_1
XFILLER_235_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_307 _15990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16561_ _16561_/A vssd1 vssd1 vccd1 vccd1 _22432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_250_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_318 _16107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13773_ _13807_/A _14039_/C vssd1 vssd1 vccd1 vccd1 _13773_/Y sky130_fd_sc_hd__nor2_1
XINSDIODE2_329 _19987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18300_ _18317_/A _18305_/C vssd1 vssd1 vccd1 vccd1 _18300_/Y sky130_fd_sc_hd__nor2_1
X_15512_ _16144_/S _15512_/B vssd1 vssd1 vccd1 vccd1 _15512_/Y sky130_fd_sc_hd__nand2_1
X_12724_ _23224_/Q _23192_/Q _23160_/Q _23128_/Q _12716_/X _12717_/X vssd1 vssd1 vccd1
+ vccd1 _12725_/B sky130_fd_sc_hd__mux4_2
XFILLER_31_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19280_ _19337_/S vssd1 vssd1 vccd1 vccd1 _19289_/S sky130_fd_sc_hd__clkbuf_8
X_16492_ _16492_/A vssd1 vssd1 vccd1 vccd1 _22403_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_349_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18231_ _22904_/Q _18240_/B vssd1 vssd1 vccd1 vccd1 _18231_/X sky130_fd_sc_hd__or2_1
XFILLER_231_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15443_ _15729_/S vssd1 vssd1 vccd1 vccd1 _16138_/S sky130_fd_sc_hd__clkbuf_4
X_12655_ _12047_/A _12654_/X _12700_/A vssd1 vssd1 vccd1 vccd1 _12655_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_231_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_318_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18162_ _18162_/A _18178_/B vssd1 vssd1 vccd1 vccd1 _18162_/X sky130_fd_sc_hd__or2b_1
X_11606_ _12256_/A vssd1 vssd1 vccd1 vccd1 _11723_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_12_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15374_ _15374_/A vssd1 vssd1 vccd1 vccd1 _22272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12586_ _12586_/A _12586_/B vssd1 vssd1 vccd1 vccd1 _12586_/X sky130_fd_sc_hd__or2_1
X_17113_ _17230_/A vssd1 vssd1 vccd1 vccd1 _17113_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_318_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14325_ _14319_/X _14323_/Y _14850_/S vssd1 vssd1 vccd1 vccd1 _14325_/X sky130_fd_sc_hd__mux2_2
X_18093_ _22869_/Q _18081_/X _18092_/X _18090_/X vssd1 vssd1 vccd1 vccd1 _22869_/D
+ sky130_fd_sc_hd__o211a_1
X_11537_ _11537_/A vssd1 vssd1 vccd1 vccd1 _11537_/X sky130_fd_sc_hd__buf_4
XFILLER_144_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_333_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17044_ _13440_/B _17043_/X _17144_/A vssd1 vssd1 vccd1 vccd1 _17044_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_356_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_305_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14256_ _14331_/S vssd1 vssd1 vccd1 vccd1 _14651_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_333_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11468_ _11468_/A vssd1 vssd1 vccd1 vccd1 _21771_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13207_ _23421_/Q _23037_/Q _23389_/Q _23357_/Q _13090_/S _13195_/X vssd1 vssd1 vccd1
+ vccd1 _13207_/X sky130_fd_sc_hd__mux4_2
X_14187_ _14187_/A vssd1 vssd1 vccd1 vccd1 _21335_/B sky130_fd_sc_hd__buf_2
X_11399_ _14178_/A _12087_/A _11763_/B vssd1 vssd1 vccd1 vccd1 _11400_/A sky130_fd_sc_hd__a21oi_2
XFILLER_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_314_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_313_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13138_ _13542_/A _14274_/B vssd1 vssd1 vccd1 vccd1 _13491_/A sky130_fd_sc_hd__and2_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _16883_/X _23194_/Q _19001_/S vssd1 vssd1 vccd1 vccd1 _18996_/A sky130_fd_sc_hd__mux2_1
XFILLER_313_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_286_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _13131_/A _13069_/B vssd1 vssd1 vccd1 vccd1 _13069_/Y sky130_fd_sc_hd__nor2_1
X_17946_ _20808_/A vssd1 vssd1 vccd1 vccd1 _21220_/A sky130_fd_sc_hd__buf_8
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17877_ _17877_/A vssd1 vssd1 vccd1 vccd1 _22809_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_254_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19616_ _19616_/A vssd1 vssd1 vccd1 vccd1 _23455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_253_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16828_ _19178_/A vssd1 vssd1 vccd1 vccd1 _16828_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_281_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19547_ _19255_/X _23425_/Q _19549_/S vssd1 vssd1 vccd1 vccd1 _19548_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16759_ _16759_/A _16759_/B vssd1 vssd1 vccd1 vccd1 _16760_/A sky130_fd_sc_hd__or2_1
XFILLER_326_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19478_ _19478_/A vssd1 vssd1 vccd1 vccd1 _23394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_250_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18429_ _22971_/Q _18429_/B vssd1 vssd1 vccd1 vccd1 _18435_/C sky130_fd_sc_hd__and2_1
XFILLER_222_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21440_ _21431_/A _21366_/X _21419_/X _21439_/Y _21175_/X vssd1 vssd1 vccd1 vccd1
+ _23915_/D sky130_fd_sc_hd__o221a_1
XFILLER_119_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_309_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21371_ _23816_/Q _23750_/Q vssd1 vssd1 vccd1 vccd1 _21372_/B sky130_fd_sc_hd__or2_1
XFILLER_336_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_308_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23110_ _23526_/CLK _23110_/D vssd1 vssd1 vccd1 vccd1 _23110_/Q sky130_fd_sc_hd__dfxtp_1
X_20322_ _20226_/X _21920_/A _20321_/X vssd1 vssd1 vccd1 vccd1 _21153_/A sky130_fd_sc_hd__a21oi_4
XFILLER_162_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_351_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_317_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_305_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23041_ _23451_/CLK _23041_/D vssd1 vssd1 vccd1 vccd1 _23041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20253_ _20213_/X _20630_/A _20252_/X _20246_/X vssd1 vssd1 vccd1 vccd1 _23663_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_190_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_288_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_333_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20184_ _23655_/Q _20223_/B vssd1 vssd1 vccd1 vccd1 _20184_/X sky130_fd_sc_hd__or2_1
XFILLER_289_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_331_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_292_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23943_ _23946_/CLK _23943_/D vssd1 vssd1 vccd1 vccd1 _23943_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23874_ _23874_/CLK _23874_/D vssd1 vssd1 vccd1 vccd1 _23874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22825_ _22830_/CLK _22825_/D vssd1 vssd1 vccd1 vccd1 _22825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_272_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22756_ _23578_/CLK _22756_/D vssd1 vssd1 vccd1 vccd1 _22756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_358_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21707_ _21708_/A _21708_/B vssd1 vssd1 vccd1 vccd1 _21709_/A sky130_fd_sc_hd__nand2_1
XFILLER_347_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22687_ _23054_/CLK _22687_/D vssd1 vssd1 vccd1 vccd1 _22687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_358_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12440_ _23888_/Q _13472_/A _12344_/X vssd1 vssd1 vccd1 vccd1 _12440_/X sky130_fd_sc_hd__a21o_1
X_21638_ _23920_/Q _15280_/A _21593_/B vssd1 vssd1 vccd1 vccd1 _21638_/X sky130_fd_sc_hd__a21o_1
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12371_ _12371_/A _12371_/B vssd1 vssd1 vccd1 vccd1 _12371_/X sky130_fd_sc_hd__or2_1
X_21569_ _22171_/B vssd1 vssd1 vccd1 vccd1 _21569_/X sky130_fd_sc_hd__buf_2
XFILLER_165_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14110_ _22888_/Q _14110_/B _22887_/Q _14121_/D vssd1 vssd1 vccd1 vccd1 _18198_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_315_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11322_ _11527_/A vssd1 vssd1 vccd1 vccd1 _11323_/A sky130_fd_sc_hd__buf_6
X_23308_ _23500_/CLK _23308_/D vssd1 vssd1 vccd1 vccd1 _23308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_299_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15090_ _15090_/A _15090_/B vssd1 vssd1 vccd1 vccd1 _15090_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14041_ _14041_/A vssd1 vssd1 vccd1 vccd1 _14041_/X sky130_fd_sc_hd__clkbuf_2
XTAP_7110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23239_ _23559_/CLK _23239_/D vssd1 vssd1 vccd1 vccd1 _23239_/Q sky130_fd_sc_hd__dfxtp_1
X_11253_ _14172_/C _11382_/B _14815_/C vssd1 vssd1 vccd1 vccd1 _12206_/A sky130_fd_sc_hd__and3_1
XTAP_7121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11184_ _13268_/A vssd1 vssd1 vccd1 vccd1 _11424_/A sky130_fd_sc_hd__buf_2
XFILLER_133_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17800_ _22775_/Q _17642_/X _17802_/S vssd1 vssd1 vccd1 vccd1 _17801_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15992_ _16109_/A _15992_/B vssd1 vssd1 vccd1 vccd1 _15992_/Y sky130_fd_sc_hd__nand2_1
X_18780_ _23111_/Q _18779_/X _18786_/S vssd1 vssd1 vccd1 vccd1 _18781_/A sky130_fd_sc_hd__mux2_1
XTAP_6475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17731_ _17731_/A vssd1 vssd1 vccd1 vccd1 _22744_/D sky130_fd_sc_hd__clkbuf_1
X_14943_ _12600_/A _14254_/X _14761_/X vssd1 vssd1 vccd1 vccd1 _14943_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_294_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14874_ _23816_/Q _14464_/X _14870_/X _14873_/X _14612_/X vssd1 vssd1 vccd1 vccd1
+ _14874_/X sky130_fd_sc_hd__a221o_1
X_17662_ _17730_/S vssd1 vssd1 vccd1 vccd1 _17671_/S sky130_fd_sc_hd__buf_6
XFILLER_224_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19401_ _23360_/Q _18859_/X _19405_/S vssd1 vssd1 vccd1 vccd1 _19402_/A sky130_fd_sc_hd__mux2_1
XFILLER_251_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13825_ _15576_/A _14021_/C vssd1 vssd1 vccd1 vccd1 _13874_/B sky130_fd_sc_hd__or2_1
X_16613_ _16613_/A vssd1 vssd1 vccd1 vccd1 _22455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_291_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17593_ _17593_/A vssd1 vssd1 vccd1 vccd1 _22692_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_104 _21596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_115 _20264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_126 _21340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19332_ _19332_/A vssd1 vssd1 vccd1 vccd1 _23329_/D sky130_fd_sc_hd__clkbuf_1
X_16544_ _14893_/X _22425_/Q _16546_/S vssd1 vssd1 vccd1 vccd1 _16545_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_137 _20334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_349_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_148 _13836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13756_ _13786_/A _13756_/B vssd1 vssd1 vccd1 vccd1 _13757_/A sky130_fd_sc_hd__and2_1
XINSDIODE2_159 _19969_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12707_ _12707_/A vssd1 vssd1 vccd1 vccd1 _12707_/X sky130_fd_sc_hd__buf_2
XFILLER_231_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19263_ _19263_/A vssd1 vssd1 vccd1 vccd1 _23299_/D sky130_fd_sc_hd__clkbuf_1
X_16475_ _16475_/A vssd1 vssd1 vccd1 vccd1 _22395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_338_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13687_ _14204_/A vssd1 vssd1 vccd1 vccd1 _13688_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_349_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18214_ _22898_/Q _18214_/B vssd1 vssd1 vccd1 vccd1 _18214_/X sky130_fd_sc_hd__or2_1
X_15426_ _15565_/A vssd1 vssd1 vccd1 vccd1 _15480_/A sky130_fd_sc_hd__clkbuf_2
X_12638_ _22309_/Q _23445_/Q _12978_/S vssd1 vssd1 vccd1 vccd1 _12638_/X sky130_fd_sc_hd__mux2_1
XPHY_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19194_ _19194_/A vssd1 vssd1 vccd1 vccd1 _19194_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18145_ _18164_/A _18144_/Y _18018_/A vssd1 vssd1 vccd1 vccd1 _18158_/S sky130_fd_sc_hd__o21a_2
X_15357_ _23824_/Q _14464_/X _15353_/X _15356_/X _14612_/X vssd1 vssd1 vccd1 vccd1
+ _15357_/X sky130_fd_sc_hd__a221o_2
XFILLER_356_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12569_ _23305_/Q _23273_/Q _23241_/Q _23529_/Q _11699_/A _11840_/A vssd1 vssd1 vccd1
+ vccd1 _12570_/B sky130_fd_sc_hd__mux4_1
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_318_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14308_ _14317_/S _13525_/B _14307_/X vssd1 vssd1 vccd1 vccd1 _14308_/Y sky130_fd_sc_hd__o21ai_1
X_18076_ hold5/A _18066_/X _18074_/X _18075_/X vssd1 vssd1 vccd1 vccd1 _22863_/D sky130_fd_sc_hd__o211a_1
XFILLER_172_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15288_ _13739_/A _15675_/B _15287_/Y _13875_/C vssd1 vssd1 vccd1 vccd1 _15288_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17027_ _22556_/Q _16922_/X _16973_/X _17026_/X vssd1 vssd1 vccd1 vccd1 _22556_/D
+ sky130_fd_sc_hd__a211o_1
X_14239_ _15033_/S vssd1 vssd1 vccd1 vccd1 _15052_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_171_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_320_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_286_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_314_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18978_ _18978_/A vssd1 vssd1 vccd1 vccd1 _23186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17929_ _22821_/Q _17922_/X _17918_/X input262/X _17915_/X vssd1 vssd1 vccd1 vccd1
+ _17929_/X sky130_fd_sc_hd__a221o_1
XFILLER_227_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20940_ _20970_/A vssd1 vssd1 vccd1 vccd1 _20940_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_281_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20871_ _20871_/A vssd1 vssd1 vccd1 vccd1 _23774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_281_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22610_ _23646_/CLK _22610_/D vssd1 vssd1 vccd1 vccd1 _22610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23590_ _23592_/CLK _23590_/D vssd1 vssd1 vccd1 vccd1 _23590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22541_ _23100_/CLK _22541_/D vssd1 vssd1 vccd1 vccd1 _22541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22472_ _22632_/CLK _22472_/D vssd1 vssd1 vccd1 vccd1 _22472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_337_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_309_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21423_ _21431_/A _21441_/A _21421_/Y _20502_/A _21422_/X vssd1 vssd1 vccd1 vccd1
+ _21452_/B sky130_fd_sc_hd__a221o_1
XFILLER_136_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_324_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21354_ _21575_/A vssd1 vssd1 vccd1 vccd1 _22091_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_135_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_351_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20305_ _20305_/A vssd1 vssd1 vccd1 vccd1 _20396_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_312_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21285_ _21285_/A vssd1 vssd1 vccd1 vccd1 _21379_/A sky130_fd_sc_hd__buf_4
XFILLER_146_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_351_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23024_ _23504_/CLK _23024_/D vssd1 vssd1 vccd1 vccd1 _23024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20236_ _20236_/A _20236_/B vssd1 vssd1 vccd1 vccd1 _20236_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_89_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23073_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20167_ _20404_/B vssd1 vssd1 vccd1 vccd1 _20177_/A sky130_fd_sc_hd__buf_2
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23367_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20098_ _23640_/Q _23639_/Q _20098_/C _20098_/D vssd1 vssd1 vccd1 vccd1 _20112_/C
+ sky130_fd_sc_hd__and4_1
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23926_ _23926_/CLK _23926_/D vssd1 vssd1 vccd1 vccd1 _23926_/Q sky130_fd_sc_hd__dfxtp_2
X_11940_ _11940_/A _13528_/B vssd1 vssd1 vccd1 vccd1 _13518_/B sky130_fd_sc_hd__nor2_1
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_291_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_273_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11871_ _11926_/A _11871_/B vssd1 vssd1 vccd1 vccd1 _11871_/X sky130_fd_sc_hd__or2_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23857_ _23862_/CLK _23857_/D vssd1 vssd1 vccd1 vccd1 _23857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13610_ _13619_/A _13531_/X _12005_/Y vssd1 vssd1 vccd1 vccd1 _13611_/B sky130_fd_sc_hd__o21a_1
XFILLER_38_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22808_ _23588_/CLK _22808_/D vssd1 vssd1 vccd1 vccd1 _22808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _22915_/Q _15259_/B vssd1 vssd1 vccd1 vccd1 _14590_/X sky130_fd_sc_hd__and2_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_343_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23788_ _23911_/CLK _23788_/D vssd1 vssd1 vccd1 vccd1 _23788_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13541_ _13492_/X _13540_/A _13632_/B _13540_/X _13579_/A vssd1 vssd1 vccd1 vccd1
+ _13573_/B sky130_fd_sc_hd__o221a_1
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22739_ _23583_/CLK _22739_/D vssd1 vssd1 vccd1 vccd1 _22739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16260_ _22309_/Q _16259_/X _16269_/S vssd1 vssd1 vccd1 vccd1 _16261_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ _13472_/A _13472_/B vssd1 vssd1 vccd1 vccd1 _14199_/A sky130_fd_sc_hd__nor2_1
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15211_ _15211_/A vssd1 vssd1 vccd1 vccd1 _15211_/X sky130_fd_sc_hd__clkbuf_2
X_12423_ _12423_/A _12423_/B vssd1 vssd1 vccd1 vccd1 _12423_/Y sky130_fd_sc_hd__nand2_1
XFILLER_200_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16191_ _16191_/A _16191_/B vssd1 vssd1 vccd1 vccd1 _16191_/Y sky130_fd_sc_hd__nand2_1
XFILLER_328_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_327_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15142_ _23660_/Q _15353_/B vssd1 vssd1 vccd1 vccd1 _15142_/X sky130_fd_sc_hd__or2_1
XFILLER_355_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_337_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12354_ _23208_/Q _23176_/Q _23144_/Q _23112_/Q _11113_/A _12199_/X vssd1 vssd1 vccd1
+ vccd1 _12354_/X sky130_fd_sc_hd__mux4_2
XFILLER_342_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_315_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_299_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11305_ _11305_/A vssd1 vssd1 vccd1 vccd1 _11637_/A sky130_fd_sc_hd__buf_6
XFILLER_126_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_343_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19950_ _19950_/A _19950_/B vssd1 vssd1 vccd1 vccd1 _19950_/Y sky130_fd_sc_hd__nor2_1
X_15073_ _23846_/Q _14737_/X _15072_/X vssd1 vssd1 vccd1 vccd1 _15073_/X sky130_fd_sc_hd__o21a_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12285_ _12606_/A _12605_/A vssd1 vssd1 vccd1 vccd1 _12287_/A sky130_fd_sc_hd__and2_2
XFILLER_107_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18901_ _23152_/Q _18808_/X _18907_/S vssd1 vssd1 vccd1 vccd1 _18902_/A sky130_fd_sc_hd__mux2_1
X_14024_ _14023_/X _13741_/B _14013_/X input245/X vssd1 vssd1 vccd1 vccd1 _14024_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_316_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11236_ _11236_/A vssd1 vssd1 vccd1 vccd1 _11236_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19881_ _16259_/X _23573_/Q _19887_/S vssd1 vssd1 vccd1 vccd1 _19882_/A sky130_fd_sc_hd__mux2_1
XFILLER_316_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_296_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18832_ _18832_/A vssd1 vssd1 vccd1 vccd1 _23127_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_295_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11167_ _13096_/A vssd1 vssd1 vccd1 vccd1 _11207_/A sky130_fd_sc_hd__buf_4
XFILLER_310_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_353_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_311_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18763_ _16908_/X _23106_/Q _18763_/S vssd1 vssd1 vccd1 vccd1 _18764_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15975_ _19245_/A vssd1 vssd1 vccd1 vccd1 _15975_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11098_ _15775_/A vssd1 vssd1 vccd1 vccd1 _11099_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17714_ _17714_/A vssd1 vssd1 vccd1 vccd1 _22736_/D sky130_fd_sc_hd__clkbuf_1
X_14926_ _15346_/A _14903_/X _14925_/X _14748_/X vssd1 vssd1 vccd1 vccd1 _14926_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_236_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18694_ _18694_/A vssd1 vssd1 vccd1 vccd1 _23075_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17645_ _18871_/A vssd1 vssd1 vccd1 vccd1 _17645_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14857_ _14843_/X _14849_/Y _14856_/Y _15292_/S vssd1 vssd1 vccd1 vccd1 _16057_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_91_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ _13808_/A vssd1 vssd1 vccd1 vccd1 _13808_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14788_ _14855_/A vssd1 vssd1 vccd1 vccd1 _15088_/S sky130_fd_sc_hd__clkbuf_2
X_17576_ _22687_/Q _17575_/X _17576_/S vssd1 vssd1 vccd1 vccd1 _17577_/A sky130_fd_sc_hd__mux2_1
X_19315_ _19315_/A vssd1 vssd1 vccd1 vccd1 _23321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_251_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13739_ _13739_/A vssd1 vssd1 vccd1 vccd1 _13739_/X sky130_fd_sc_hd__buf_2
X_16527_ _16527_/A vssd1 vssd1 vccd1 vccd1 _22419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19246_ _19246_/A vssd1 vssd1 vccd1 vccd1 _19259_/S sky130_fd_sc_hd__buf_4
X_16458_ _18625_/B _19843_/B vssd1 vssd1 vccd1 vccd1 _16515_/A sky130_fd_sc_hd__or2_4
XFILLER_32_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15409_ _14800_/A _15393_/X _15408_/Y _14586_/A vssd1 vssd1 vccd1 vccd1 _15409_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_19177_ _19177_/A vssd1 vssd1 vccd1 vccd1 _23272_/D sky130_fd_sc_hd__clkbuf_1
X_16389_ _16389_/A vssd1 vssd1 vccd1 vccd1 _22357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_334_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18128_ _18116_/Y _18126_/X _18127_/X _18121_/X vssd1 vssd1 vccd1 vccd1 _22880_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18059_ hold6/A _18052_/X _18053_/X _22990_/Q _18054_/X vssd1 vssd1 vccd1 vccd1 _18059_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_160_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21070_ _23843_/Q _21072_/B vssd1 vssd1 vccd1 vccd1 _21070_/X sky130_fd_sc_hd__or2_1
XFILLER_259_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20021_ _23616_/Q _23615_/Q _20021_/C _20031_/D vssd1 vssd1 vccd1 vccd1 _20034_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_141_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_287_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_286_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21972_ _21972_/A _21972_/B vssd1 vssd1 vccd1 vccd1 _21972_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23711_ _23714_/CLK _23711_/D vssd1 vssd1 vccd1 vccd1 _23711_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20923_ _13945_/B _20922_/X _20626_/B _20912_/X vssd1 vssd1 vccd1 vccd1 _20923_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_227_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23642_ _23643_/CLK _23642_/D vssd1 vssd1 vccd1 vccd1 _23642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20854_ _20711_/B _20846_/X _20847_/X _23770_/Q vssd1 vssd1 vccd1 vccd1 _20855_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23573_ _23573_/CLK _23573_/D vssd1 vssd1 vccd1 vccd1 _23573_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_136_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _22968_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20785_ _13454_/Y _20773_/Y _20583_/B _21148_/A vssd1 vssd1 vccd1 vccd1 _20785_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_148_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_490 _13967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_356_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_329_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22524_ _23368_/CLK _22524_/D vssd1 vssd1 vccd1 vccd1 _22524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22455_ _23558_/CLK _22455_/D vssd1 vssd1 vccd1 vccd1 _22455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_315_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_339_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21406_ _21406_/A _22224_/B vssd1 vssd1 vccd1 vccd1 _21406_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22386_ _23522_/CLK _22386_/D vssd1 vssd1 vccd1 vccd1 _22386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_352_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21337_ _15826_/A _15631_/A _21336_/X _23888_/Q vssd1 vssd1 vccd1 vccd1 _21342_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_324_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_352_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_297_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12070_ _22467_/Q _22627_/Q _12070_/S vssd1 vssd1 vccd1 vccd1 _12071_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21268_ _15929_/X _21242_/X _21267_/Y _21236_/X vssd1 vssd1 vccd1 vccd1 _23903_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23007_ _23009_/CLK _23007_/D vssd1 vssd1 vccd1 vccd1 _23007_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_132_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20219_ _20305_/A vssd1 vssd1 vccd1 vccd1 _20275_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_320_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21199_ _21199_/A _21199_/B vssd1 vssd1 vccd1 vccd1 _21199_/Y sky130_fd_sc_hd__nand2_1
XFILLER_293_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15760_ _23769_/Q _14911_/A _14913_/A _15758_/X _15759_/X vssd1 vssd1 vccd1 vccd1
+ _15760_/X sky130_fd_sc_hd__a221o_1
X_12972_ _13091_/A _12972_/B vssd1 vssd1 vccd1 vccd1 _12972_/Y sky130_fd_sc_hd__nor2_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _23912_/Q _14814_/C _23913_/Q vssd1 vssd1 vccd1 vccd1 _21339_/B sky130_fd_sc_hd__o21ai_2
X_11923_ _12144_/A _11917_/X _11922_/X _11348_/A vssd1 vssd1 vccd1 vccd1 _11923_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_346_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23909_ _23945_/CLK _23909_/D vssd1 vssd1 vccd1 vccd1 _23909_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15691_ _23831_/Q _15211_/X _15687_/X _15690_/X _15222_/X vssd1 vssd1 vccd1 vccd1
+ _15691_/X sky130_fd_sc_hd__a221o_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _22627_/Q _16249_/X _17432_/S vssd1 vssd1 vccd1 vccd1 _17431_/A sky130_fd_sc_hd__mux2_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14642_ _14636_/X _14640_/X _14852_/S vssd1 vssd1 vccd1 vccd1 _14642_/X sky130_fd_sc_hd__mux2_2
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ _23470_/Q _23566_/Q _22530_/Q _22334_/Q _11770_/A _12246_/A vssd1 vssd1 vccd1
+ vccd1 _11854_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14573_ _15114_/S vssd1 vssd1 vccd1 vccd1 _14967_/S sky130_fd_sc_hd__clkbuf_4
X_17361_ _22601_/Q input195/X _17369_/S vssd1 vssd1 vccd1 vccd1 _17362_/A sky130_fd_sc_hd__mux2_1
XFILLER_260_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11785_ _11905_/A _11785_/B vssd1 vssd1 vccd1 vccd1 _11785_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19100_ _23240_/Q _18782_/X _19102_/S vssd1 vssd1 vccd1 vccd1 _19101_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16312_ _16368_/A vssd1 vssd1 vccd1 vccd1 _16381_/S sky130_fd_sc_hd__buf_6
X_13524_ _13524_/A vssd1 vssd1 vccd1 vccd1 _13524_/Y sky130_fd_sc_hd__inv_2
X_17292_ _22166_/A _17291_/X _17292_/S vssd1 vssd1 vccd1 vccd1 _17292_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16243_ _18808_/A vssd1 vssd1 vccd1 vccd1 _16243_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19031_ _19088_/S vssd1 vssd1 vccd1 vccd1 _19040_/S sky130_fd_sc_hd__clkbuf_8
X_13455_ _13455_/A _13455_/B _13455_/C vssd1 vssd1 vccd1 vccd1 _13455_/Y sky130_fd_sc_hd__nor3_4
XFILLER_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12406_ _12406_/A _12406_/B vssd1 vssd1 vccd1 vccd1 _12406_/Y sky130_fd_sc_hd__nor2_1
X_16174_ _23844_/Q _15593_/A _16170_/X _16173_/X _14922_/A vssd1 vssd1 vccd1 vccd1
+ _16174_/X sky130_fd_sc_hd__a221o_1
XFILLER_12_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13386_ _13386_/A _13386_/B _13383_/X _13385_/Y vssd1 vssd1 vccd1 vccd1 _13387_/D
+ sky130_fd_sc_hd__or4bb_4
XFILLER_126_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_315_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15125_ _12234_/X _14254_/X _14761_/X _12236_/B _14837_/X vssd1 vssd1 vccd1 vccd1
+ _15125_/X sky130_fd_sc_hd__a221o_1
XFILLER_115_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12337_ _11683_/A _12323_/X _12336_/X _12594_/A vssd1 vssd1 vccd1 vccd1 _21444_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_303_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_342_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19933_ _19934_/B _19934_/C _23595_/Q vssd1 vssd1 vccd1 vccd1 _19935_/B sky130_fd_sc_hd__a21oi_1
XFILLER_287_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15056_ _15056_/A _15056_/B vssd1 vssd1 vccd1 vccd1 _15484_/A sky130_fd_sc_hd__nand2_2
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12268_ _12410_/A _12268_/B vssd1 vssd1 vccd1 vccd1 _12268_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14007_ input215/X _14004_/X _14006_/X vssd1 vssd1 vccd1 vccd1 _14007_/X sky130_fd_sc_hd__a21o_4
X_11219_ _11219_/A vssd1 vssd1 vccd1 vccd1 _15929_/A sky130_fd_sc_hd__buf_8
X_19864_ _19864_/A vssd1 vssd1 vccd1 vccd1 _23565_/D sky130_fd_sc_hd__clkbuf_1
X_12199_ _12458_/A vssd1 vssd1 vccd1 vccd1 _12199_/X sky130_fd_sc_hd__buf_4
XFILLER_295_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18815_ _23122_/Q _18814_/X _18818_/S vssd1 vssd1 vccd1 vccd1 _18816_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19795_ _19841_/S vssd1 vssd1 vccd1 vccd1 _19804_/S sky130_fd_sc_hd__buf_4
XFILLER_95_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18746_ _16883_/X _23098_/Q _18752_/S vssd1 vssd1 vccd1 vccd1 _18747_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15958_ _23838_/Q _15593_/X _15954_/X _15957_/X _14738_/X vssd1 vssd1 vccd1 vccd1
+ _15958_/X sky130_fd_sc_hd__a221o_1
XFILLER_255_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput190 localMemory_wb_adr_i[0] vssd1 vssd1 vccd1 vccd1 input190/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14909_ _23657_/Q _15985_/B vssd1 vssd1 vccd1 vccd1 _14909_/X sky130_fd_sc_hd__or2_1
X_18677_ _18677_/A vssd1 vssd1 vccd1 vccd1 _23067_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15889_ _15872_/X _15888_/Y _16188_/A vssd1 vssd1 vccd1 vccd1 _15889_/X sky130_fd_sc_hd__o21a_1
X_17628_ _22703_/Q _17626_/X _17640_/S vssd1 vssd1 vccd1 vccd1 _17629_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17559_ _18785_/A vssd1 vssd1 vccd1 vccd1 _17559_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_211_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20570_ _20570_/A vssd1 vssd1 vccd1 vccd1 _20571_/A sky130_fd_sc_hd__inv_2
XFILLER_20_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19229_ _19229_/A vssd1 vssd1 vccd1 vccd1 _19229_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22240_ _23778_/Q _22240_/B vssd1 vssd1 vccd1 vccd1 _22242_/C sky130_fd_sc_hd__xnor2_1
XFILLER_353_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_307_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22171_ _22171_/A _22171_/B vssd1 vssd1 vccd1 vccd1 _22171_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21122_ _21122_/A vssd1 vssd1 vccd1 vccd1 _21134_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_274_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21053_ _20713_/A _21047_/X _21052_/X _21049_/X vssd1 vssd1 vccd1 vccd1 _23835_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20004_ _23613_/Q _20014_/C _23614_/Q vssd1 vssd1 vccd1 vccd1 _20008_/B sky130_fd_sc_hd__a21oi_1
XFILLER_274_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_290_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_286_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21955_ _21569_/X _21953_/X _21954_/Y _21577_/X vssd1 vssd1 vccd1 vccd1 _21956_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_55_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_299_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20906_ _20948_/A vssd1 vssd1 vccd1 vccd1 _20906_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21886_ _23831_/Q _21885_/X _21973_/S vssd1 vssd1 vccd1 vccd1 _21886_/X sky130_fd_sc_hd__mux2_2
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23625_ _23634_/CLK _23625_/D vssd1 vssd1 vccd1 vccd1 _23625_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_74_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_306_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20837_ _20843_/A _20837_/B vssd1 vssd1 vccd1 vccd1 _20838_/A sky130_fd_sc_hd__and2_1
XFILLER_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_329_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11570_ _12985_/A _11570_/B vssd1 vssd1 vccd1 vccd1 _11570_/Y sky130_fd_sc_hd__nor2_1
X_23556_ _23556_/CLK _23556_/D vssd1 vssd1 vccd1 vccd1 _23556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20768_ _20768_/A _20888_/B _20768_/C vssd1 vssd1 vccd1 vccd1 _20768_/X sky130_fd_sc_hd__or3_1
XFILLER_195_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22507_ _23693_/CLK _22507_/D vssd1 vssd1 vccd1 vccd1 _22507_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_52_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23487_ _23551_/CLK _23487_/D vssd1 vssd1 vccd1 vccd1 _23487_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_344_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20699_ _20759_/B vssd1 vssd1 vccd1 vccd1 _20731_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_318_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13240_ _13240_/A vssd1 vssd1 vccd1 vccd1 _13240_/Y sky130_fd_sc_hd__inv_2
X_22438_ _23541_/CLK _22438_/D vssd1 vssd1 vccd1 vccd1 _22438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13171_ _23422_/Q _23038_/Q _23390_/Q _23358_/Q _13114_/A _13127_/A vssd1 vssd1 vccd1
+ vccd1 _13172_/B sky130_fd_sc_hd__mux4_1
XFILLER_170_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22369_ _23571_/CLK _22369_/D vssd1 vssd1 vccd1 vccd1 _22369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_353_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_325_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_313_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12122_ _12071_/A _12119_/X _12121_/X vssd1 vssd1 vccd1 vccd1 _12122_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_33_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23580_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_324_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_297_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12053_ _23411_/Q _23027_/Q _23379_/Q _23347_/Q _12675_/A _12746_/A vssd1 vssd1 vccd1
+ vccd1 _12053_/X sky130_fd_sc_hd__mux4_1
X_16930_ _22809_/Q _17244_/B vssd1 vssd1 vccd1 vccd1 _16950_/B sky130_fd_sc_hd__and2_1
XFILLER_313_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_293_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16861_ _16860_/X _22535_/Q _16861_/S vssd1 vssd1 vccd1 vccd1 _16862_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18600_ _16879_/X _23033_/Q _18608_/S vssd1 vssd1 vccd1 vccd1 _18601_/A sky130_fd_sc_hd__mux2_1
XFILLER_281_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15812_ _22967_/Q _15811_/X _15982_/B vssd1 vssd1 vccd1 vccd1 _15812_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19580_ _23439_/Q _19197_/A _19588_/S vssd1 vssd1 vccd1 vccd1 _19581_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16792_ _16795_/A _16792_/B vssd1 vssd1 vccd1 vccd1 _16793_/A sky130_fd_sc_hd__or2_1
XFILLER_77_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18531_ _18520_/X _18530_/Y _18264_/A vssd1 vssd1 vccd1 vccd1 _23007_/D sky130_fd_sc_hd__a21oi_1
XFILLER_292_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12955_ _12995_/A _12955_/B vssd1 vssd1 vccd1 vccd1 _12955_/X sky130_fd_sc_hd__or2_1
XFILLER_246_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15743_ _15480_/X _13599_/X _15663_/X _15742_/X vssd1 vssd1 vccd1 vccd1 _15743_/X
+ sky130_fd_sc_hd__o211a_2
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11906_ _23469_/Q _23565_/Q _22529_/Q _22333_/Q _11574_/A _11696_/X vssd1 vssd1 vccd1
+ vccd1 _11906_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18462_ _22981_/Q _18465_/B vssd1 vssd1 vccd1 vccd1 _18462_/Y sky130_fd_sc_hd__nand2_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _12886_/A _12886_/B vssd1 vssd1 vccd1 vccd1 _12886_/Y sky130_fd_sc_hd__nor2_1
XFILLER_179_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _15674_/A vssd1 vssd1 vccd1 vccd1 _15674_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_233_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17413_ _22619_/Q _16223_/X _17421_/S vssd1 vssd1 vccd1 vccd1 _17414_/A sky130_fd_sc_hd__mux2_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14625_ _14949_/S vssd1 vssd1 vccd1 vccd1 _14854_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_11837_ _11837_/A _11837_/B vssd1 vssd1 vccd1 vccd1 _11837_/Y sky130_fd_sc_hd__nand2_1
X_18393_ _18401_/A _18393_/B _18394_/B vssd1 vssd1 vccd1 vccd1 _22958_/D sky130_fd_sc_hd__nor3_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17344_ _17344_/A vssd1 vssd1 vccd1 vccd1 _22593_/D sky130_fd_sc_hd__clkbuf_1
X_14556_ _16530_/A _21294_/A _16953_/B _14556_/D vssd1 vssd1 vccd1 vccd1 _14557_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11768_ _12567_/A vssd1 vssd1 vccd1 vccd1 _11853_/A sky130_fd_sc_hd__buf_2
XFILLER_320_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13507_ _14791_/A _12443_/A _13505_/X _13464_/B _13506_/X vssd1 vssd1 vccd1 vccd1
+ _13902_/B sky130_fd_sc_hd__a221o_2
XFILLER_347_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17275_ _22579_/Q _17255_/X _17240_/X _17274_/X vssd1 vssd1 vccd1 vccd1 _22579_/D
+ sky130_fd_sc_hd__a211o_1
X_14487_ _23749_/Q _14482_/X _14486_/X _23653_/Q vssd1 vssd1 vccd1 vccd1 _14487_/X
+ sky130_fd_sc_hd__a22o_1
X_11699_ _11699_/A vssd1 vssd1 vccd1 vccd1 _11700_/A sky130_fd_sc_hd__buf_8
XFILLER_228_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19014_ _16911_/X _23203_/Q _19016_/S vssd1 vssd1 vccd1 vccd1 _19015_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16226_ _16226_/A vssd1 vssd1 vccd1 vccd1 _22298_/D sky130_fd_sc_hd__clkbuf_1
X_13438_ _20532_/A vssd1 vssd1 vccd1 vccd1 _13439_/A sky130_fd_sc_hd__buf_2
XFILLER_335_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16157_ _14175_/A _15478_/X _16195_/S vssd1 vssd1 vccd1 vccd1 _16157_/X sky130_fd_sc_hd__a21o_1
XFILLER_350_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13369_ _13913_/A _13369_/B vssd1 vssd1 vccd1 vccd1 _13370_/D sky130_fd_sc_hd__xnor2_1
XFILLER_303_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_331_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_288_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15108_ _15187_/A _14246_/B _15107_/X _13688_/A _22518_/Q vssd1 vssd1 vccd1 vccd1
+ _15109_/B sky130_fd_sc_hd__o32ai_4
XFILLER_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16088_ _18862_/A vssd1 vssd1 vccd1 vccd1 _19255_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_288_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19916_ _19922_/D vssd1 vssd1 vccd1 vccd1 _19916_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15039_ _14819_/X _15036_/X _15038_/Y _14698_/X vssd1 vssd1 vccd1 vccd1 _15039_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_331_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_296_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19847_ _19847_/A vssd1 vssd1 vccd1 vccd1 _23557_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19778_ _23527_/Q _19172_/A _19782_/S vssd1 vssd1 vccd1 vccd1 _19779_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_329_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18729_ _18729_/A vssd1 vssd1 vccd1 vccd1 _23090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21740_ _21740_/A _21740_/B vssd1 vssd1 vccd1 vccd1 _21740_/X sky130_fd_sc_hd__xor2_1
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21671_ _21640_/A _21640_/B _21637_/A vssd1 vssd1 vccd1 vccd1 _21675_/A sky130_fd_sc_hd__o21ai_1
XFILLER_225_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23410_ _23474_/CLK _23410_/D vssd1 vssd1 vccd1 vccd1 _23410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20622_ _20622_/A vssd1 vssd1 vccd1 vccd1 _20623_/A sky130_fd_sc_hd__inv_2
XFILLER_189_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23341_ _23407_/CLK _23341_/D vssd1 vssd1 vccd1 vccd1 _23341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_338_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_327_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20553_ _11069_/D _20642_/A _20733_/A vssd1 vssd1 vccd1 vccd1 _20553_/X sky130_fd_sc_hd__a21o_1
XFILLER_354_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23272_ _23496_/CLK _23272_/D vssd1 vssd1 vccd1 vccd1 _23272_/Q sky130_fd_sc_hd__dfxtp_1
X_20484_ _23712_/Q _20416_/B _20482_/Y _20483_/X vssd1 vssd1 vccd1 vccd1 _23712_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_307_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_1_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
X_22223_ _22223_/A _22223_/B vssd1 vssd1 vccd1 vccd1 _22223_/X sky130_fd_sc_hd__or2_1
XFILLER_98_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_307_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22154_ _23841_/Q _22153_/Y _22190_/B vssd1 vssd1 vccd1 vccd1 _22154_/X sky130_fd_sc_hd__mux2_1
XFILLER_306_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput450 _22886_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[1] sky130_fd_sc_hd__buf_2
XFILLER_105_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_350_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput461 _23911_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[0] sky130_fd_sc_hd__buf_2
XTAP_6827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21105_ _23850_/Q _21096_/X _21098_/X _20580_/A vssd1 vssd1 vccd1 vccd1 _21106_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput472 _23912_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[1] sky130_fd_sc_hd__buf_2
XTAP_6838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput483 _23913_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[2] sky130_fd_sc_hd__buf_2
X_22085_ _22085_/A _22085_/B vssd1 vssd1 vccd1 vccd1 _22085_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_303_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput494 _23946_/Q vssd1 vssd1 vccd1 vccd1 probe_state[1] sky130_fd_sc_hd__buf_2
XFILLER_99_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21036_ _21185_/A vssd1 vssd1 vccd1 vccd1 _21163_/A sky130_fd_sc_hd__buf_4
XFILLER_102_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_151_wb_clk_i _23945_/CLK vssd1 vssd1 vccd1 vccd1 _23861_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_290_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22987_ _23009_/CLK _22987_/D vssd1 vssd1 vccd1 vccd1 _22987_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_234_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ _21899_/A _21900_/A _13500_/A vssd1 vssd1 vccd1 vccd1 _12807_/A sky130_fd_sc_hd__mux2_2
XFILLER_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21938_ _21877_/Y _21876_/X _21934_/C _21936_/X _21937_/Y vssd1 vssd1 vccd1 vccd1
+ _22040_/A sky130_fd_sc_hd__a311o_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12671_ _12671_/A vssd1 vssd1 vccd1 vccd1 _12672_/A sky130_fd_sc_hd__buf_4
XFILLER_242_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21869_ _13432_/B _21336_/B _21868_/X vssd1 vssd1 vccd1 vccd1 _21869_/X sky130_fd_sc_hd__a21o_1
XFILLER_70_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _22905_/Q _14153_/X _14151_/X _22598_/Q vssd1 vssd1 vccd1 vccd1 _14551_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_230_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23608_ _23637_/CLK _23608_/D vssd1 vssd1 vccd1 vccd1 _23608_/Q sky130_fd_sc_hd__dfxtp_2
X_11622_ _23318_/Q _23286_/Q _23254_/Q _23542_/Q _11893_/S _11621_/X vssd1 vssd1 vccd1
+ vccd1 _11623_/B sky130_fd_sc_hd__mux4_1
XFILLER_231_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _15455_/A _15387_/X _15389_/X vssd1 vssd1 vccd1 vccd1 _15390_/X sky130_fd_sc_hd__o21a_1
XFILLER_179_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_357_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14341_ _14339_/X _14340_/X _14351_/S vssd1 vssd1 vccd1 vccd1 _14341_/X sky130_fd_sc_hd__mux2_1
X_23539_ _23572_/CLK _23539_/D vssd1 vssd1 vccd1 vccd1 _23539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11553_ _13234_/S vssd1 vssd1 vccd1 vccd1 _13296_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_329_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_357_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17060_ input75/X input104/X _17084_/S vssd1 vssd1 vccd1 vccd1 _17060_/X sky130_fd_sc_hd__mux2_8
XFILLER_345_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_317_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14272_ _14268_/X _14270_/X _14310_/S vssd1 vssd1 vccd1 vccd1 _14272_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11484_ _11476_/Y _11478_/Y _11480_/Y _11482_/Y _11483_/X vssd1 vssd1 vccd1 vccd1
+ _11485_/C sky130_fd_sc_hd__o221a_1
XFILLER_7_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_344_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16011_ _16007_/X _16009_/Y _22119_/A _15321_/X vssd1 vssd1 vccd1 vccd1 _18856_/A
+ sky130_fd_sc_hd__a2bb2o_4
X_13223_ _12745_/X _13216_/X _13218_/X _13222_/X vssd1 vssd1 vccd1 vccd1 _13223_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_195_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_298_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_298_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_325_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13154_ _13158_/A _13154_/B vssd1 vssd1 vccd1 vccd1 _13154_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_345_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_297_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12105_ _12105_/A _12105_/B vssd1 vssd1 vccd1 vccd1 _12105_/X sky130_fd_sc_hd__or2_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _22831_/Q _17956_/X _17959_/X input277/X _17951_/X vssd1 vssd1 vccd1 vccd1
+ _17962_/X sky130_fd_sc_hd__a221o_1
X_13085_ _13096_/A vssd1 vssd1 vccd1 vccd1 _13085_/X sky130_fd_sc_hd__clkbuf_4
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_297_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19701_ _19769_/S vssd1 vssd1 vccd1 vccd1 _19710_/S sky130_fd_sc_hd__buf_6
X_12036_ _12027_/Y _12031_/Y _12033_/Y _12035_/Y _11657_/X vssd1 vssd1 vccd1 vccd1
+ _12037_/C sky130_fd_sc_hd__o221a_1
X_16913_ _16913_/A vssd1 vssd1 vccd1 vccd1 _22551_/D sky130_fd_sc_hd__clkbuf_1
X_17893_ _17971_/A vssd1 vssd1 vccd1 vccd1 _18097_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19632_ _19169_/X _23462_/Q _19638_/S vssd1 vssd1 vccd1 vccd1 _19633_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16844_ _19194_/A vssd1 vssd1 vccd1 vccd1 _16844_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_293_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_293_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19563_ _19563_/A vssd1 vssd1 vccd1 vccd1 _23431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_281_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16775_ _16775_/A vssd1 vssd1 vccd1 vccd1 _22509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13987_ _14220_/A _13993_/A vssd1 vssd1 vccd1 vccd1 _13990_/A sky130_fd_sc_hd__or2_4
XFILLER_93_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18514_ _18507_/X _18513_/Y _18503_/X vssd1 vssd1 vccd1 vccd1 _23000_/D sky130_fd_sc_hd__a21oi_1
XFILLER_230_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15726_ _22965_/Q _15726_/B vssd1 vssd1 vccd1 vccd1 _15726_/X sky130_fd_sc_hd__or2_1
XFILLER_34_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _12931_/Y _12933_/Y _12935_/Y _12937_/Y _11246_/A vssd1 vssd1 vccd1 vccd1
+ _12938_/X sky130_fd_sc_hd__o221a_1
XFILLER_230_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19494_ _19178_/X _23401_/Q _19494_/S vssd1 vssd1 vccd1 vccd1 _19495_/A sky130_fd_sc_hd__mux2_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18445_ _19950_/A _18445_/B vssd1 vssd1 vccd1 vccd1 _18445_/Y sky130_fd_sc_hd__nor2_1
XFILLER_234_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15657_ _15345_/A _15641_/X _15656_/Y _15697_/A vssd1 vssd1 vccd1 vccd1 _15657_/Y
+ sky130_fd_sc_hd__o22ai_1
X_12869_ _13492_/A vssd1 vssd1 vccd1 vccd1 _13592_/A sky130_fd_sc_hd__buf_4
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14608_ _23750_/Q _14482_/X _14478_/X _14600_/X _14607_/X vssd1 vssd1 vccd1 vccd1
+ _14608_/X sky130_fd_sc_hd__a221o_1
X_18376_ _18401_/A _18376_/B _18377_/B vssd1 vssd1 vccd1 vccd1 _22952_/D sky130_fd_sc_hd__nor3_1
XFILLER_15_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15588_ _22930_/Q vssd1 vssd1 vccd1 vccd1 _18314_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_221_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17327_ _17371_/A vssd1 vssd1 vccd1 vccd1 _17335_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_202_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14539_ _14538_/X _22249_/D _14539_/S vssd1 vssd1 vccd1 vccd1 _18770_/A sky130_fd_sc_hd__mux2_2
XFILLER_30_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17258_ _17258_/A vssd1 vssd1 vccd1 vccd1 _17258_/Y sky130_fd_sc_hd__inv_2
XFILLER_336_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_335_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16209_ _22293_/Q _16200_/X _16221_/S vssd1 vssd1 vccd1 vccd1 _16210_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_351_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17189_ _22571_/Q _17141_/X _17131_/X _17188_/X vssd1 vssd1 vccd1 vccd1 _22571_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_289_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_303_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22910_ _22923_/CLK _22910_/D vssd1 vssd1 vccd1 vccd1 _22910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23890_ _23907_/CLK _23890_/D vssd1 vssd1 vccd1 vccd1 _23890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22841_ _22893_/CLK _22841_/D vssd1 vssd1 vccd1 vccd1 _22841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22772_ _23391_/CLK _22772_/D vssd1 vssd1 vccd1 vccd1 _22772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21723_ _21721_/X _21720_/X _21719_/Y _21718_/Y vssd1 vssd1 vccd1 vccd1 _21724_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_80_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_303_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21654_ _21653_/B _21653_/C _21653_/A vssd1 vssd1 vccd1 vccd1 _21694_/B sky130_fd_sc_hd__a21oi_2
X_20605_ _20605_/A _20631_/B vssd1 vssd1 vccd1 vccd1 _20608_/B sky130_fd_sc_hd__nor2_2
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21585_ _21585_/A _21585_/B vssd1 vssd1 vccd1 vccd1 _21587_/A sky130_fd_sc_hd__nand2_1
XFILLER_138_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_326_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23324_ _23419_/CLK _23324_/D vssd1 vssd1 vccd1 vccd1 _23324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_296_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20536_ _20781_/A _20536_/B _20779_/A vssd1 vssd1 vccd1 vccd1 _20544_/A sky130_fd_sc_hd__or3_2
XFILLER_137_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_315_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23255_ _23543_/CLK _23255_/D vssd1 vssd1 vccd1 vccd1 _23255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_342_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20467_ _20467_/A vssd1 vssd1 vccd1 vccd1 _20467_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_307_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22206_ _22206_/A _22206_/B vssd1 vssd1 vccd1 vccd1 _22207_/B sky130_fd_sc_hd__nand2_2
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23186_ _23538_/CLK _23186_/D vssd1 vssd1 vccd1 vccd1 _23186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20398_ _23683_/Q _20404_/B vssd1 vssd1 vccd1 vccd1 _20398_/X sky130_fd_sc_hd__or2_1
XTAP_6602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22137_ _22242_/B _22137_/B vssd1 vssd1 vccd1 vccd1 _22137_/Y sky130_fd_sc_hd__nand2_1
XTAP_7369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput291 _14096_/X vssd1 vssd1 vccd1 vccd1 addr0[6] sky130_fd_sc_hd__buf_2
XTAP_5923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22068_ _21594_/B _22066_/X _22067_/Y _21677_/X vssd1 vssd1 vccd1 vccd1 _22068_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_6679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13910_ _15037_/A vssd1 vssd1 vccd1 vccd1 _13910_/X sky130_fd_sc_hd__buf_6
X_21019_ _20622_/A _21008_/X _21018_/X _21010_/X vssd1 vssd1 vccd1 vccd1 _23822_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14890_ _22981_/Q _14137_/A _14980_/A input240/X vssd1 vssd1 vccd1 vccd1 _21406_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_331_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13841_ _13874_/C vssd1 vssd1 vccd1 vccd1 _13864_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_262_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_308 _18856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13772_ _14021_/C _13739_/A _13771_/X _13730_/X vssd1 vssd1 vccd1 vccd1 _14039_/C
+ sky130_fd_sc_hd__a22oi_4
X_16560_ _15324_/X _22432_/Q _16568_/S vssd1 vssd1 vccd1 vccd1 _16561_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_319 _16107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15511_ _15440_/X _15504_/X _15510_/Y _15150_/A vssd1 vssd1 vccd1 vccd1 _15512_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_12723_ _12707_/X _12712_/X _12715_/X _12722_/X _11378_/A vssd1 vssd1 vccd1 vccd1
+ _12738_/B sky130_fd_sc_hd__a311o_2
X_16491_ _15523_/X _22403_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _16492_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18230_ _18243_/A vssd1 vssd1 vccd1 vccd1 _18240_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_349_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12654_ _23477_/Q _23573_/Q _22537_/Q _22341_/Q _12680_/A _12041_/A vssd1 vssd1 vccd1
+ vccd1 _12654_/X sky130_fd_sc_hd__mux4_2
X_15442_ _23666_/Q _15905_/B vssd1 vssd1 vccd1 vccd1 _15442_/X sky130_fd_sc_hd__or2_1
XFILLER_188_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11605_ _12365_/A vssd1 vssd1 vccd1 vccd1 _12256_/A sky130_fd_sc_hd__buf_6
X_18161_ _22891_/Q vssd1 vssd1 vccd1 vccd1 _18162_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_230_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15373_ _15372_/X _22272_/Q _15524_/S vssd1 vssd1 vccd1 vccd1 _15374_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12585_ _22361_/Q _22393_/Q _22682_/Q _23049_/Q _11799_/A _12329_/X vssd1 vssd1 vccd1
+ vccd1 _12586_/B sky130_fd_sc_hd__mux4_2
XFILLER_318_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17112_ input81/X input46/X _17132_/S vssd1 vssd1 vccd1 vccd1 _17112_/X sky130_fd_sc_hd__mux2_8
XFILLER_156_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11536_ _13180_/A _11536_/B vssd1 vssd1 vccd1 vccd1 _11536_/X sky130_fd_sc_hd__or2_1
X_14324_ _14635_/A vssd1 vssd1 vccd1 vccd1 _14850_/S sky130_fd_sc_hd__buf_2
X_18092_ _22868_/Q _18082_/X _18083_/X _23001_/Q _18084_/X vssd1 vssd1 vccd1 vccd1
+ _18092_/X sky130_fd_sc_hd__a221o_1
XFILLER_318_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_317_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17043_ _23466_/Q _16987_/X _16988_/X _17042_/X _15005_/B vssd1 vssd1 vccd1 vccd1
+ _17043_/X sky130_fd_sc_hd__a32o_1
XFILLER_184_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14255_ _14290_/A vssd1 vssd1 vccd1 vccd1 _14331_/S sky130_fd_sc_hd__clkbuf_2
X_11467_ _15630_/A _11466_/X _11288_/X vssd1 vssd1 vccd1 vccd1 _11467_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_333_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_298_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13206_ _13206_/A _13206_/B vssd1 vssd1 vccd1 vccd1 _13206_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14186_ _14814_/C vssd1 vssd1 vccd1 vccd1 _14713_/C sky130_fd_sc_hd__buf_4
X_11398_ _11398_/A vssd1 vssd1 vccd1 vccd1 _16005_/A sky130_fd_sc_hd__buf_4
XFILLER_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13137_ _13139_/B vssd1 vssd1 vccd1 vccd1 _14274_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_97_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_341_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18994_ _18994_/A vssd1 vssd1 vccd1 vccd1 _23193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_313_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_297_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _22826_/Q _17938_/X _17896_/X _17944_/X _17933_/X vssd1 vssd1 vccd1 vccd1
+ _17945_/X sky130_fd_sc_hd__a221o_1
XFILLER_300_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13068_ _23232_/Q _23200_/Q _23168_/Q _23136_/Q _13275_/A _11527_/X vssd1 vssd1 vccd1
+ vccd1 _13069_/B sky130_fd_sc_hd__mux4_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12019_ _12949_/A _12019_/B vssd1 vssd1 vccd1 vccd1 _12019_/Y sky130_fd_sc_hd__nor2_1
XFILLER_239_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17876_ _22809_/Q input247/X _17882_/S vssd1 vssd1 vccd1 vccd1 _17877_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_294_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19615_ _23455_/Q _19249_/A _19621_/S vssd1 vssd1 vccd1 vccd1 _19616_/A sky130_fd_sc_hd__mux2_1
XFILLER_254_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16827_ _16827_/A vssd1 vssd1 vccd1 vccd1 _22524_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19546_ _19546_/A vssd1 vssd1 vccd1 vccd1 _23424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16758_ _22505_/Q _16747_/X _16748_/X input19/X vssd1 vssd1 vccd1 vccd1 _16759_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_253_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_326_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15709_ _18830_/A vssd1 vssd1 vccd1 vccd1 _19223_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19477_ _23394_/Q _18865_/X _19477_/S vssd1 vssd1 vccd1 vccd1 _19478_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16689_ _16729_/A vssd1 vssd1 vccd1 vccd1 _16689_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18428_ _19923_/A _18428_/B _18429_/B vssd1 vssd1 vccd1 vccd1 _22970_/D sky130_fd_sc_hd__nor3_1
XFILLER_250_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18359_ _22947_/Q _18359_/B vssd1 vssd1 vccd1 vccd1 _18366_/C sky130_fd_sc_hd__and2_1
XFILLER_222_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21370_ _23816_/Q _23750_/Q vssd1 vssd1 vccd1 vccd1 _21372_/A sky130_fd_sc_hd__nand2_1
XFILLER_175_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_336_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20321_ _20376_/A _20318_/X _20319_/Y _20320_/X vssd1 vssd1 vccd1 vccd1 _20321_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_323_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23040_ _23264_/CLK _23040_/D vssd1 vssd1 vccd1 vccd1 _23040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_289_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20252_ _23663_/Q _20277_/B vssd1 vssd1 vccd1 vccd1 _20252_/X sky130_fd_sc_hd__or2_1
XFILLER_171_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_288_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20183_ _20404_/B vssd1 vssd1 vccd1 vccd1 _20223_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_249_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23942_ _23942_/CLK _23942_/D vssd1 vssd1 vccd1 vccd1 _23942_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_285_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23873_ _23874_/CLK _23873_/D vssd1 vssd1 vccd1 vccd1 _23873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22824_ _23583_/CLK _22824_/D vssd1 vssd1 vccd1 vccd1 _22824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22755_ _23459_/CLK _22755_/D vssd1 vssd1 vccd1 vccd1 _22755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_345_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21706_ _23825_/Q _21705_/Y _22019_/A vssd1 vssd1 vccd1 vccd1 _21706_/X sky130_fd_sc_hd__mux2_1
X_22686_ _23367_/CLK _22686_/D vssd1 vssd1 vccd1 vccd1 _22686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_358_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21637_ _21637_/A _21637_/B vssd1 vssd1 vccd1 vccd1 _21640_/A sky130_fd_sc_hd__nand2_1
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12370_ _12370_/A _13763_/A vssd1 vssd1 vccd1 vccd1 _12370_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21568_ _23821_/Q _21838_/A _21567_/Y _21377_/A vssd1 vssd1 vccd1 vccd1 _21568_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_197_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11321_ _11533_/A vssd1 vssd1 vccd1 vccd1 _11527_/A sky130_fd_sc_hd__clkbuf_4
X_23307_ _23467_/CLK _23307_/D vssd1 vssd1 vccd1 vccd1 _23307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_355_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20519_ _23707_/Q _20524_/B _20519_/C vssd1 vssd1 vccd1 vccd1 _20520_/D sky130_fd_sc_hd__and3_1
XFILLER_154_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_314_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21499_ _21500_/A _21500_/B vssd1 vssd1 vccd1 vccd1 _21513_/A sky130_fd_sc_hd__nor2_1
XFILLER_299_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14040_ input221/X _14038_/X _14039_/X vssd1 vssd1 vccd1 vccd1 _14040_/X sky130_fd_sc_hd__a21bo_4
XTAP_7100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23238_ _23526_/CLK _23238_/D vssd1 vssd1 vccd1 vccd1 _23238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11252_ _11382_/C vssd1 vssd1 vccd1 vccd1 _14815_/C sky130_fd_sc_hd__clkbuf_4
XTAP_7111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23169_ _23451_/CLK _23169_/D vssd1 vssd1 vccd1 vccd1 _23169_/Q sky130_fd_sc_hd__dfxtp_1
X_11183_ _13051_/A vssd1 vssd1 vccd1 vccd1 _13268_/A sky130_fd_sc_hd__buf_2
XFILLER_350_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ _14516_/A _15984_/X _15990_/Y _15652_/X vssd1 vssd1 vccd1 vccd1 _15992_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17730_ _22744_/Q _17645_/X _17730_/S vssd1 vssd1 vccd1 vccd1 _17731_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14942_ _14942_/A vssd1 vssd1 vccd1 vccd1 _14942_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_342_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17661_ _17717_/A vssd1 vssd1 vccd1 vccd1 _17730_/S sky130_fd_sc_hd__buf_6
XFILLER_349_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14873_ _23752_/Q _14482_/X _14478_/X _14871_/X _14872_/X vssd1 vssd1 vccd1 vccd1
+ _14873_/X sky130_fd_sc_hd__a221o_1
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19400_ _19400_/A vssd1 vssd1 vccd1 vccd1 _23359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16612_ _22455_/Q _16211_/X _16618_/S vssd1 vssd1 vccd1 vccd1 _16613_/A sky130_fd_sc_hd__mux2_1
XFILLER_263_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13824_ _12839_/B _13808_/X _13781_/X vssd1 vssd1 vccd1 vccd1 _13824_/X sky130_fd_sc_hd__a21o_1
XFILLER_29_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17592_ _22692_/Q _17591_/X _17592_/S vssd1 vssd1 vccd1 vccd1 _17593_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_105 _21596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_116 _12424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19331_ _19255_/X _23329_/Q _19333_/S vssd1 vssd1 vccd1 vccd1 _19332_/A sky130_fd_sc_hd__mux2_1
XFILLER_251_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_127 _21340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16543_ _16543_/A vssd1 vssd1 vccd1 vccd1 _22424_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_138 _13022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13755_ _13803_/A _13730_/X _13771_/B _13739_/X _14015_/C vssd1 vssd1 vccd1 vccd1
+ _13756_/B sky130_fd_sc_hd__a32o_2
XFILLER_204_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_149 _13242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_349_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19262_ _19261_/X _23299_/Q _19265_/S vssd1 vssd1 vccd1 vccd1 _19263_/A sky130_fd_sc_hd__mux2_1
X_12706_ _23930_/Q vssd1 vssd1 vccd1 vccd1 _21899_/A sky130_fd_sc_hd__inv_2
XFILLER_43_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16474_ _15104_/X _22395_/Q _16480_/S vssd1 vssd1 vccd1 vccd1 _16475_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13686_ _13686_/A _13686_/B _13583_/A vssd1 vssd1 vccd1 vccd1 _14204_/A sky130_fd_sc_hd__or3b_4
X_18213_ _22849_/Q _18202_/X _18212_/X _18206_/X vssd1 vssd1 vccd1 vccd1 _22897_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_176_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15425_ _15425_/A vssd1 vssd1 vccd1 vccd1 _21720_/A sky130_fd_sc_hd__buf_8
XPHY_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12637_ _12685_/A vssd1 vssd1 vccd1 vccd1 _12637_/X sky130_fd_sc_hd__buf_6
X_19193_ _19193_/A vssd1 vssd1 vccd1 vccd1 _23277_/D sky130_fd_sc_hd__clkbuf_1
XPHY_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_318_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18144_ _18163_/B _18144_/B vssd1 vssd1 vccd1 vccd1 _18144_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12568_ _23401_/Q _23017_/Q _23369_/Q _23337_/Q _11148_/A _11840_/X vssd1 vssd1 vccd1
+ vccd1 _12568_/X sky130_fd_sc_hd__mux4_1
X_15356_ _23760_/Q _14482_/X _14478_/X _15354_/X _15355_/X vssd1 vssd1 vccd1 vccd1
+ _15356_/X sky130_fd_sc_hd__a221o_2
XFILLER_8_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11519_ _11519_/A vssd1 vssd1 vccd1 vccd1 _11519_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_172_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14307_ _14330_/S _14307_/B vssd1 vssd1 vccd1 vccd1 _14307_/X sky130_fd_sc_hd__or2_1
XFILLER_7_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18075_ _18105_/A vssd1 vssd1 vccd1 vccd1 _18075_/X sky130_fd_sc_hd__buf_2
XFILLER_305_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15287_ _15287_/A _15432_/B vssd1 vssd1 vccd1 vccd1 _15287_/Y sky130_fd_sc_hd__nand2_2
X_12499_ _22261_/Q _23077_/Q _23493_/Q _22422_/Q _23894_/Q _23895_/Q vssd1 vssd1 vccd1
+ vccd1 _12500_/B sky130_fd_sc_hd__mux4_1
XFILLER_144_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17026_ _17000_/X _17015_/X _17025_/X _17012_/X vssd1 vssd1 vccd1 vccd1 _17026_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_236_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14238_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14238_/X sky130_fd_sc_hd__buf_4
XFILLER_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_302_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_302_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_299_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14169_ _14609_/A vssd1 vssd1 vccd1 vccd1 _15066_/B sky130_fd_sc_hd__buf_2
XFILLER_124_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_286_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18977_ _16857_/X _23186_/Q _18979_/S vssd1 vssd1 vccd1 vccd1 _18978_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17928_ _22821_/Q _17914_/X _17927_/X _17912_/X vssd1 vssd1 vccd1 vccd1 _22821_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_267_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17859_ _22801_/Q _17623_/X _17859_/S vssd1 vssd1 vccd1 vccd1 _17860_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_332_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20870_ _20879_/A _20870_/B vssd1 vssd1 vccd1 vccd1 _20871_/A sky130_fd_sc_hd__and2_1
XFILLER_81_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19529_ _19540_/A vssd1 vssd1 vccd1 vccd1 _19538_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_223_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22540_ _23544_/CLK _22540_/D vssd1 vssd1 vccd1 vccd1 _22540_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_223_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22471_ _23480_/CLK _22471_/D vssd1 vssd1 vccd1 vccd1 _22471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_337_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21422_ _21422_/A _21615_/A vssd1 vssd1 vccd1 vccd1 _21422_/X sky130_fd_sc_hd__and2_1
XFILLER_337_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_337_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21353_ _21353_/A _21353_/B vssd1 vssd1 vccd1 vccd1 _21353_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_324_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20304_ _15656_/Y _20295_/X _20306_/B vssd1 vssd1 vccd1 vccd1 _20304_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_324_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21284_ _21079_/A _21199_/B _21283_/Y _21281_/X vssd1 vssd1 vccd1 vccd1 _23910_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_293_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23023_ _23535_/CLK _23023_/D vssd1 vssd1 vccd1 vccd1 _23023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_293_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20235_ _15230_/X _20169_/A _20236_/B vssd1 vssd1 vccd1 vccd1 _20235_/X sky130_fd_sc_hd__a21o_1
XFILLER_304_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20166_ _20344_/A vssd1 vssd1 vccd1 vccd1 _20404_/B sky130_fd_sc_hd__buf_2
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_292_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20097_ _23640_/Q _20110_/C vssd1 vssd1 vccd1 vccd1 _20100_/B sky130_fd_sc_hd__nor2_1
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23925_ _23936_/CLK _23925_/D vssd1 vssd1 vccd1 vccd1 _23925_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_58_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23510_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _22366_/Q _22398_/Q _22687_/Q _23054_/Q _12094_/A _11869_/X vssd1 vssd1 vccd1
+ vccd1 _11871_/B sky130_fd_sc_hd__mux4_1
XFILLER_233_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23856_ _23856_/CLK _23856_/D vssd1 vssd1 vccd1 vccd1 _23856_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_309_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22807_ _23893_/CLK _22807_/D vssd1 vssd1 vccd1 vccd1 _22807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23787_ _23862_/CLK _23787_/D vssd1 vssd1 vccd1 vccd1 _23787_/Q sky130_fd_sc_hd__dfxtp_4
X_20999_ _21072_/B vssd1 vssd1 vccd1 vccd1 _21009_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13540_ _13540_/A _13632_/C vssd1 vssd1 vccd1 vccd1 _13540_/X sky130_fd_sc_hd__or2_1
X_22738_ _23549_/CLK _22738_/D vssd1 vssd1 vccd1 vccd1 _22738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_347_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ _13471_/A _23945_/Q vssd1 vssd1 vccd1 vccd1 _13603_/A sky130_fd_sc_hd__or2_4
X_22669_ _23580_/CLK _22669_/D vssd1 vssd1 vccd1 vccd1 _22669_/Q sky130_fd_sc_hd__dfxtp_1
X_15210_ _15210_/A vssd1 vssd1 vccd1 vccd1 _15210_/X sky130_fd_sc_hd__buf_4
XFILLER_40_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12422_ _22456_/Q _22616_/Q _12424_/S vssd1 vssd1 vccd1 vccd1 _12423_/B sky130_fd_sc_hd__mux2_1
X_16190_ _14568_/A _16165_/Y _16189_/X vssd1 vssd1 vccd1 vccd1 _16190_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_343_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_328_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15141_ _23596_/Q _14450_/X _14455_/X _23628_/Q vssd1 vssd1 vccd1 vccd1 _15141_/X
+ sky130_fd_sc_hd__o22a_2
X_12353_ _11138_/A _12348_/Y _12350_/Y _12352_/Y vssd1 vssd1 vccd1 vccd1 _12353_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_153_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_337_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_342_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11304_ _11821_/A vssd1 vssd1 vccd1 vccd1 _11305_/A sky130_fd_sc_hd__buf_6
X_15072_ _23691_/Q _15222_/A _15066_/X _15071_/X _14745_/Y vssd1 vssd1 vccd1 vccd1
+ _15072_/X sky130_fd_sc_hd__a221o_1
XFILLER_303_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12284_ _11884_/B _20217_/A _12283_/X vssd1 vssd1 vccd1 vccd1 _12605_/A sky130_fd_sc_hd__o21a_4
XFILLER_114_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14023_ _14083_/A vssd1 vssd1 vccd1 vccd1 _14023_/X sky130_fd_sc_hd__buf_2
X_18900_ _18900_/A vssd1 vssd1 vccd1 vccd1 _23151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_330_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11235_ _11235_/A vssd1 vssd1 vccd1 vccd1 _11236_/A sky130_fd_sc_hd__buf_6
XFILLER_181_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19880_ _19880_/A vssd1 vssd1 vccd1 vccd1 _23572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18831_ _23127_/Q _18830_/X _18834_/S vssd1 vssd1 vccd1 vccd1 _18832_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_353_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11166_ _11166_/A vssd1 vssd1 vccd1 vccd1 _13096_/A sky130_fd_sc_hd__buf_4
XTAP_6240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_14_0_wb_clk_i clkbuf_3_7_1_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_14_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_310_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18762_ _18762_/A vssd1 vssd1 vccd1 vccd1 _23105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15974_ _18852_/A vssd1 vssd1 vccd1 vccd1 _19245_/A sky130_fd_sc_hd__clkbuf_2
XTAP_6295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11097_ _13472_/B vssd1 vssd1 vccd1 vccd1 _15775_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17713_ _22736_/Q _17620_/X _17715_/S vssd1 vssd1 vccd1 vccd1 _17714_/A sky130_fd_sc_hd__mux2_1
XTAP_5583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14925_ _23689_/Q _14905_/X _14924_/X vssd1 vssd1 vccd1 vccd1 _14925_/X sky130_fd_sc_hd__o21a_2
XTAP_5594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18693_ _23075_/Q _17642_/X _18695_/S vssd1 vssd1 vccd1 vccd1 _18694_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ _17644_/A vssd1 vssd1 vccd1 vccd1 _22708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_291_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14856_ _15490_/S _14852_/X _14855_/X vssd1 vssd1 vccd1 vccd1 _14856_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_64_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13807_ _13807_/A _14046_/C vssd1 vssd1 vccd1 vccd1 _13807_/Y sky130_fd_sc_hd__nor2_1
XFILLER_302_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17575_ _18801_/A vssd1 vssd1 vccd1 vccd1 _17575_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14787_ _14785_/X _15086_/A _15018_/S vssd1 vssd1 vccd1 vccd1 _14787_/X sky130_fd_sc_hd__mux2_1
XFILLER_302_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11999_ _22469_/Q _22629_/Q _22308_/Q _23444_/Q _12733_/A _12844_/A vssd1 vssd1 vccd1
+ vccd1 _11999_/X sky130_fd_sc_hd__mux4_1
X_19314_ _19229_/X _23321_/Q _19322_/S vssd1 vssd1 vccd1 vccd1 _19315_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16526_ _16161_/X _22419_/Q _16528_/S vssd1 vssd1 vccd1 vccd1 _16527_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13738_ _13738_/A vssd1 vssd1 vccd1 vccd1 _13739_/A sky130_fd_sc_hd__buf_2
XFILLER_149_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19245_ _19245_/A vssd1 vssd1 vccd1 vccd1 _19245_/X sky130_fd_sc_hd__clkbuf_2
X_16457_ _16203_/B _16457_/B _16457_/C vssd1 vssd1 vccd1 vccd1 _19843_/B sky130_fd_sc_hd__nand3b_2
X_13669_ _13669_/A _16927_/A vssd1 vssd1 vccd1 vccd1 _14147_/B sky130_fd_sc_hd__nor2_1
XFILLER_337_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15408_ _15408_/A vssd1 vssd1 vccd1 vccd1 _15408_/Y sky130_fd_sc_hd__inv_2
XFILLER_319_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_318_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19176_ _19175_/X _23272_/Q _19179_/S vssd1 vssd1 vccd1 vccd1 _19177_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16388_ _14534_/X _22357_/Q _16396_/S vssd1 vssd1 vccd1 vccd1 _16389_/A sky130_fd_sc_hd__mux2_1
XFILLER_319_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18127_ _18116_/A _14107_/X _22880_/Q vssd1 vssd1 vccd1 vccd1 _18127_/X sky130_fd_sc_hd__a21o_1
XFILLER_157_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15339_ _14847_/X _14852_/X _15339_/S vssd1 vssd1 vccd1 vccd1 _15340_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18058_ hold6/A _18051_/X _18057_/X _18045_/X vssd1 vssd1 vccd1 vccd1 _22857_/D sky130_fd_sc_hd__o211a_1
XFILLER_306_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17009_ _14196_/B _17008_/X _17009_/S vssd1 vssd1 vccd1 vccd1 _17009_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_327_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20020_ _23618_/Q _23617_/Q vssd1 vssd1 vccd1 vccd1 _20031_/D sky130_fd_sc_hd__and2_1
XFILLER_286_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21971_ _21971_/A _21971_/B vssd1 vssd1 vccd1 vccd1 _21972_/B sky130_fd_sc_hd__nor2_1
XFILLER_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23710_ _23714_/CLK _23710_/D vssd1 vssd1 vccd1 vccd1 _23710_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20922_ _20936_/A vssd1 vssd1 vccd1 vccd1 _20922_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_270_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_281_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23641_ _23643_/CLK _23641_/D vssd1 vssd1 vccd1 vccd1 _23641_/Q sky130_fd_sc_hd__dfxtp_1
X_20853_ _20853_/A vssd1 vssd1 vccd1 vccd1 _23769_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23572_ _23572_/CLK _23572_/D vssd1 vssd1 vccd1 vccd1 _23572_/Q sky130_fd_sc_hd__dfxtp_1
X_20784_ _21357_/C vssd1 vssd1 vccd1 vccd1 _21148_/A sky130_fd_sc_hd__buf_4
XFILLER_22_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_480 _20327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_491 _13972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22523_ _23367_/CLK _22523_/D vssd1 vssd1 vccd1 vccd1 _22523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_298_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22454_ _23896_/CLK _22454_/D vssd1 vssd1 vccd1 vccd1 _22454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_356_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_176_wb_clk_i _23931_/CLK vssd1 vssd1 vccd1 vccd1 _23810_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21405_ _21712_/S vssd1 vssd1 vccd1 vccd1 _22224_/B sky130_fd_sc_hd__buf_2
XFILLER_148_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_105_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23423_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22385_ _23553_/CLK _22385_/D vssd1 vssd1 vccd1 vccd1 _22385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_325_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_309_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21336_ _21336_/A _21336_/B vssd1 vssd1 vccd1 vccd1 _21336_/X sky130_fd_sc_hd__and2_2
XFILLER_151_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_352_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21267_ _21267_/A _21274_/B vssd1 vssd1 vccd1 vccd1 _21267_/Y sky130_fd_sc_hd__nand2_1
XFILLER_340_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23006_ _23009_/CLK _23006_/D vssd1 vssd1 vccd1 vccd1 _23006_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_289_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20218_ _17052_/A _20215_/X _20217_/Y vssd1 vssd1 vccd1 vccd1 _20218_/Y sky130_fd_sc_hd__o21ai_1
X_21198_ _21243_/A vssd1 vssd1 vccd1 vccd1 _21199_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20149_ _20250_/A vssd1 vssd1 vccd1 vccd1 _20236_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12971_ _23323_/Q _23291_/Q _23259_/Q _23547_/Q _12921_/S _12749_/X vssd1 vssd1 vccd1
+ vccd1 _12972_/B sky130_fd_sc_hd__mux4_2
XFILLER_292_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _21350_/B vssd1 vssd1 vccd1 vccd1 _21351_/B sky130_fd_sc_hd__buf_6
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23908_ _23910_/CLK _23908_/D vssd1 vssd1 vccd1 vccd1 _23908_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11922_ _12397_/A _11922_/B vssd1 vssd1 vccd1 vccd1 _11922_/X sky130_fd_sc_hd__or2_1
XFILLER_218_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15690_ _23767_/Q _15215_/X _15216_/X _15688_/X _15689_/X vssd1 vssd1 vccd1 vccd1
+ _15690_/X sky130_fd_sc_hd__a221o_4
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _14949_/S vssd1 vssd1 vccd1 vccd1 _14852_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23839_ _23876_/CLK _23839_/D vssd1 vssd1 vccd1 vccd1 _23839_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _11853_/A _11853_/B vssd1 vssd1 vccd1 vccd1 _11853_/Y sky130_fd_sc_hd__nor2_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17360_ _17371_/A vssd1 vssd1 vccd1 vccd1 _17369_/S sky130_fd_sc_hd__buf_2
XFILLER_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14572_ _22488_/Q _14232_/X _14247_/A _14571_/X _14071_/A vssd1 vssd1 vccd1 vccd1
+ _14572_/X sky130_fd_sc_hd__o221a_1
X_11784_ _23311_/Q _23279_/Q _23247_/Q _23535_/Q _11708_/S _11621_/X vssd1 vssd1 vccd1
+ vccd1 _11785_/B sky130_fd_sc_hd__mux4_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16311_ _19843_/A _19771_/A vssd1 vssd1 vccd1 vccd1 _16368_/A sky130_fd_sc_hd__or2_4
X_13523_ _13525_/A _13523_/B vssd1 vssd1 vccd1 vccd1 _13524_/A sky130_fd_sc_hd__and2_1
X_17291_ _21605_/A _17290_/X _17291_/S vssd1 vssd1 vccd1 vccd1 _17291_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_347_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19030_ _19030_/A vssd1 vssd1 vccd1 vccd1 _23209_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_347_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16242_ _16242_/A vssd1 vssd1 vccd1 vccd1 _22303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_335_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13454_ _13454_/A _13455_/B _13455_/C vssd1 vssd1 vccd1 vccd1 _13454_/Y sky130_fd_sc_hd__nor3_4
XFILLER_201_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_356_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12405_ _23207_/Q _23175_/Q _23143_/Q _23111_/Q _11455_/A _11733_/A vssd1 vssd1 vccd1
+ vccd1 _12406_/B sky130_fd_sc_hd__mux4_1
X_16173_ _23780_/Q _15595_/A _15596_/A _16171_/X _16172_/X vssd1 vssd1 vccd1 vccd1
+ _16173_/X sky130_fd_sc_hd__a221o_1
X_13385_ _13623_/A _13385_/B vssd1 vssd1 vccd1 vccd1 _13385_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_328_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_327_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15124_ _15122_/X _14940_/B _15123_/Y _15010_/A vssd1 vssd1 vccd1 vccd1 _15124_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_353_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12336_ _11819_/X _12327_/X _12331_/X _12335_/X _11375_/A vssd1 vssd1 vccd1 vccd1
+ _12336_/X sky130_fd_sc_hd__a311o_1
XFILLER_342_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_331_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19932_ _19932_/A vssd1 vssd1 vccd1 vccd1 _20008_/A sky130_fd_sc_hd__buf_2
X_15055_ _22517_/Q _14231_/A _14238_/A _15054_/X vssd1 vssd1 vccd1 vccd1 _15056_/B
+ sky130_fd_sc_hd__o22a_1
X_12267_ _23467_/Q _23563_/Q _22527_/Q _22331_/Q _11455_/A _11733_/A vssd1 vssd1 vccd1
+ vccd1 _12268_/B sky130_fd_sc_hd__mux4_1
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11218_ _11218_/A vssd1 vssd1 vccd1 vccd1 _11219_/A sky130_fd_sc_hd__buf_6
XFILLER_268_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14006_ _14015_/A _14036_/B _14006_/C vssd1 vssd1 vccd1 vccd1 _14006_/X sky130_fd_sc_hd__and3_1
X_19863_ _16233_/X _23565_/Q _19865_/S vssd1 vssd1 vccd1 vccd1 _19864_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12198_ _12196_/X _12197_/X _11706_/A vssd1 vssd1 vccd1 vccd1 _12198_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_311_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18814_ _18814_/A vssd1 vssd1 vccd1 vccd1 _18814_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11149_ _11770_/A vssd1 vssd1 vccd1 vccd1 _11708_/S sky130_fd_sc_hd__buf_4
XTAP_6070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19794_ _19794_/A vssd1 vssd1 vccd1 vccd1 _23534_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18745_ _18745_/A vssd1 vssd1 vccd1 vccd1 _23097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15957_ _23774_/Q _15595_/X _15596_/X _15955_/X _15956_/X vssd1 vssd1 vccd1 vccd1
+ _15957_/X sky130_fd_sc_hd__a221o_2
XTAP_5391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput180 irq[3] vssd1 vssd1 vccd1 vccd1 _20511_/C sky130_fd_sc_hd__clkbuf_4
Xinput191 localMemory_wb_adr_i[10] vssd1 vssd1 vccd1 vccd1 input191/X sky130_fd_sc_hd__clkbuf_1
X_14908_ _16137_/B vssd1 vssd1 vccd1 vccd1 _15985_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_18676_ _23067_/Q _17617_/X _18680_/S vssd1 vssd1 vccd1 vccd1 _18677_/A sky130_fd_sc_hd__mux2_1
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15888_ _15964_/A _17232_/A vssd1 vssd1 vccd1 vccd1 _15888_/Y sky130_fd_sc_hd__nor2_1
XFILLER_251_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17627_ _17627_/A vssd1 vssd1 vccd1 vccd1 _17640_/S sky130_fd_sc_hd__buf_6
XFILLER_36_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14839_ _14839_/A vssd1 vssd1 vccd1 vccd1 _14839_/X sky130_fd_sc_hd__buf_2
XFILLER_52_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17558_ _17558_/A vssd1 vssd1 vccd1 vccd1 _22681_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23531_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16509_ _15861_/X _22411_/Q _16513_/S vssd1 vssd1 vccd1 vccd1 _16510_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_339_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17489_ _17489_/A vssd1 vssd1 vccd1 vccd1 _22652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19228_ _19228_/A vssd1 vssd1 vccd1 vccd1 _23288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_347_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19159_ _23267_/Q _18868_/X _19161_/S vssd1 vssd1 vccd1 vccd1 _19160_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22170_ _22170_/A _22170_/B vssd1 vssd1 vccd1 vccd1 _22170_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_307_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_322_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21121_ _21121_/A _21121_/B vssd1 vssd1 vccd1 vccd1 _23856_/D sky130_fd_sc_hd__nor2_1
XFILLER_133_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21052_ _23835_/Q _21068_/B vssd1 vssd1 vccd1 vccd1 _21052_/X sky130_fd_sc_hd__or2_1
XFILLER_28_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_330_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20003_ _23612_/Q _23611_/Q _20003_/C _20005_/D vssd1 vssd1 vccd1 vccd1 _20014_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_98_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_290_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21954_ _21954_/A _22032_/B vssd1 vssd1 vccd1 vccd1 _21954_/Y sky130_fd_sc_hd__nor2_1
XFILLER_243_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20905_ _21400_/A _20894_/X _20583_/B _20897_/X vssd1 vssd1 vccd1 vccd1 _20905_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21885_ _21885_/A _21885_/B vssd1 vssd1 vccd1 vccd1 _21885_/X sky130_fd_sc_hd__xor2_1
XFILLER_203_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23624_ _23624_/CLK _23624_/D vssd1 vssd1 vccd1 vccd1 _23624_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20836_ _20678_/B _20828_/X _20829_/X _23765_/Q vssd1 vssd1 vccd1 vccd1 _20837_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_306_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23555_ _23555_/CLK _23555_/D vssd1 vssd1 vccd1 vccd1 _23555_/Q sky130_fd_sc_hd__dfxtp_1
X_20767_ _11270_/Y _20732_/X _20766_/Y vssd1 vssd1 vccd1 vccd1 _20768_/C sky130_fd_sc_hd__a21oi_2
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_356_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_329_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22506_ _23700_/CLK _22506_/D vssd1 vssd1 vccd1 vccd1 _22506_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_317_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23486_ _23582_/CLK _23486_/D vssd1 vssd1 vccd1 vccd1 _23486_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_195_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20698_ _20730_/A vssd1 vssd1 vccd1 vccd1 _20727_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_168_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_356_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22437_ _23510_/CLK _22437_/D vssd1 vssd1 vccd1 vccd1 _22437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_353_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13170_ _23326_/Q _23294_/Q _23262_/Q _23550_/Q _11532_/X _11544_/A vssd1 vssd1 vccd1
+ vccd1 _13170_/X sky130_fd_sc_hd__mux4_1
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22368_ _23440_/CLK _22368_/D vssd1 vssd1 vccd1 vccd1 _22368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_313_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12121_ _12073_/A _12120_/X _12082_/A vssd1 vssd1 vccd1 vccd1 _12121_/X sky130_fd_sc_hd__a21o_1
XFILLER_325_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21319_ _21319_/A _21319_/B vssd1 vssd1 vccd1 vccd1 _21319_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_340_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22299_ _23563_/CLK _22299_/D vssd1 vssd1 vccd1 vccd1 _22299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12052_ _12056_/A _12052_/B vssd1 vssd1 vccd1 vccd1 _12052_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23420_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_266_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16860_ _19210_/A vssd1 vssd1 vccd1 vccd1 _16860_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15811_ _14592_/A _15804_/X _15810_/X _14748_/A vssd1 vssd1 vccd1 vccd1 _15811_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_120_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16791_ _22514_/Q _16783_/X _16784_/X input29/X vssd1 vssd1 vccd1 vccd1 _16792_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18530_ _23007_/Q _18530_/B vssd1 vssd1 vccd1 vccd1 _18530_/Y sky130_fd_sc_hd__nand2_1
XFILLER_281_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15742_ _14568_/A _15716_/X _15741_/Y _16191_/A vssd1 vssd1 vccd1 vccd1 _15742_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _23481_/Q _23577_/Q _22541_/Q _22345_/Q _12709_/X _12710_/X vssd1 vssd1 vccd1
+ vccd1 _12955_/B sky130_fd_sc_hd__mux4_1
XFILLER_206_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _18451_/X _18460_/Y _22260_/A vssd1 vssd1 vccd1 vccd1 _22980_/D sky130_fd_sc_hd__a21oi_1
X_11905_ _11905_/A _11905_/B vssd1 vssd1 vccd1 vccd1 _11905_/Y sky130_fd_sc_hd__nor2_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15673_ _15673_/A vssd1 vssd1 vccd1 vccd1 _15891_/A sky130_fd_sc_hd__buf_4
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _22282_/Q _23098_/Q _23514_/Q _22443_/Q _12692_/X _11594_/A vssd1 vssd1 vccd1
+ vccd1 _12886_/B sky130_fd_sc_hd__mux4_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _17469_/S vssd1 vssd1 vccd1 vccd1 _17421_/S sky130_fd_sc_hd__buf_4
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14624_ _15249_/S vssd1 vssd1 vccd1 vccd1 _15339_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18392_ _22957_/Q _22958_/Q _18392_/C vssd1 vssd1 vccd1 vccd1 _18394_/B sky130_fd_sc_hd__and3_1
XFILLER_61_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11836_ _22463_/Q _22623_/Q _12554_/S vssd1 vssd1 vccd1 vccd1 _11837_/B sky130_fd_sc_hd__mux2_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _22593_/Q input210/X _17347_/S vssd1 vssd1 vccd1 vccd1 _17344_/A sky130_fd_sc_hd__mux2_1
X_14555_ _21677_/A _21293_/A vssd1 vssd1 vccd1 vccd1 _14556_/D sky130_fd_sc_hd__or2_2
XFILLER_14_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _12532_/A vssd1 vssd1 vccd1 vccd1 _12567_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13506_ _14292_/A _13506_/B vssd1 vssd1 vccd1 vccd1 _13506_/X sky130_fd_sc_hd__and2_1
X_17274_ _17242_/X _17266_/X _17273_/X _17237_/X vssd1 vssd1 vccd1 vccd1 _17274_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_159_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14486_ _14606_/A vssd1 vssd1 vccd1 vccd1 _14486_/X sky130_fd_sc_hd__clkbuf_4
X_11698_ _11698_/A _11698_/B vssd1 vssd1 vccd1 vccd1 _11698_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_347_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_307_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19013_ _19013_/A vssd1 vssd1 vccd1 vccd1 _23202_/D sky130_fd_sc_hd__clkbuf_1
X_16225_ _22298_/Q _16223_/X _16237_/S vssd1 vssd1 vccd1 vccd1 _16226_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13437_ _14177_/A vssd1 vssd1 vccd1 vccd1 _20532_/A sky130_fd_sc_hd__buf_2
XFILLER_316_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16156_ _15564_/A _16131_/A _15672_/X _16155_/X vssd1 vssd1 vccd1 vccd1 _16156_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_344_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13368_ _13356_/A _13355_/A _12602_/X vssd1 vssd1 vccd1 vccd1 _13369_/B sky130_fd_sc_hd__o21ai_1
XFILLER_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_331_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15107_ input166/X input131/X _15110_/S vssd1 vssd1 vccd1 vccd1 _15107_/X sky130_fd_sc_hd__mux2_8
XFILLER_288_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12319_ _22782_/Q _22750_/Q _22651_/Q _22718_/Q _11814_/X _11815_/X vssd1 vssd1 vccd1
+ vccd1 _12319_/X sky130_fd_sc_hd__mux4_2
X_16087_ _16083_/X _22171_/A _16195_/S vssd1 vssd1 vccd1 vccd1 _18862_/A sky130_fd_sc_hd__mux2_8
X_13299_ _13319_/A _13300_/B vssd1 vssd1 vccd1 vccd1 _13301_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19915_ _23589_/Q vssd1 vssd1 vccd1 vccd1 _19915_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_269_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15038_ _15161_/A _21442_/B vssd1 vssd1 vccd1 vccd1 _15038_/Y sky130_fd_sc_hd__nor2_1
XFILLER_269_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19846_ _16200_/X _23557_/Q _19854_/S vssd1 vssd1 vccd1 vccd1 _19847_/A sky130_fd_sc_hd__mux2_1
XFILLER_296_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16989_ _17042_/A vssd1 vssd1 vccd1 vccd1 _16989_/X sky130_fd_sc_hd__buf_2
X_19777_ _19777_/A vssd1 vssd1 vccd1 vccd1 _23526_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18728_ _16857_/X _23090_/Q _18730_/S vssd1 vssd1 vccd1 vccd1 _18729_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18659_ _18659_/A vssd1 vssd1 vccd1 vccd1 _23059_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21670_ _23824_/Q _21669_/Y _22083_/A vssd1 vssd1 vccd1 vccd1 _21670_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20621_ _23725_/Q _20593_/X _20620_/X _20602_/X vssd1 vssd1 vccd1 vccd1 _23725_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23340_ _23950_/A _23340_/D vssd1 vssd1 vccd1 vccd1 _23340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_338_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20552_ _20662_/A vssd1 vssd1 vccd1 vccd1 _20733_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23271_ _23527_/CLK _23271_/D vssd1 vssd1 vccd1 vccd1 _23271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20483_ _20602_/A vssd1 vssd1 vccd1 vccd1 _20483_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22222_ _22222_/A _22222_/B vssd1 vssd1 vccd1 vccd1 _22223_/B sky130_fd_sc_hd__and2_1
XFILLER_341_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22153_ _22153_/A _22153_/B vssd1 vssd1 vccd1 vccd1 _22153_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_322_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput440 _22586_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_stall_o sky130_fd_sc_hd__buf_2
XFILLER_161_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21104_ _21108_/A _21104_/B vssd1 vssd1 vccd1 vccd1 _23849_/D sky130_fd_sc_hd__nor2_1
Xoutput451 _22887_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[2] sky130_fd_sc_hd__buf_2
XTAP_6817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput462 _23921_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[10] sky130_fd_sc_hd__buf_2
XFILLER_105_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_350_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22084_ _23838_/Q _22190_/B _22083_/Y _21377_/A vssd1 vssd1 vccd1 vccd1 _22084_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput473 _23931_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[20] sky130_fd_sc_hd__buf_2
XFILLER_78_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput484 _23941_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[30] sky130_fd_sc_hd__buf_2
XFILLER_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput495 _13433_/X vssd1 vssd1 vccd1 vccd1 probe_takeBranch sky130_fd_sc_hd__buf_2
X_21035_ _23829_/Q _21048_/B vssd1 vssd1 vccd1 vccd1 _21035_/X sky130_fd_sc_hd__or2_1
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_304_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22986_ _23009_/CLK _22986_/D vssd1 vssd1 vccd1 vccd1 _22986_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_262_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21937_ _21937_/A vssd1 vssd1 vccd1 vccd1 _21937_/Y sky130_fd_sc_hd__inv_2
XFILLER_271_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12670_ _12818_/A _12670_/B vssd1 vssd1 vccd1 vccd1 _12670_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_191_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23397_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21868_ _21868_/A _21868_/B _21868_/C vssd1 vssd1 vccd1 vccd1 _21868_/X sky130_fd_sc_hd__or3_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23607_ _23637_/CLK _23607_/D vssd1 vssd1 vccd1 vccd1 _23607_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11621_/A vssd1 vssd1 vccd1 vccd1 _11621_/X sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_120_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23634_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_230_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20819_ _20825_/A _20819_/B vssd1 vssd1 vccd1 vccd1 _20820_/A sky130_fd_sc_hd__and2_1
XFILLER_196_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21799_ _21799_/A _21799_/B vssd1 vssd1 vccd1 vccd1 _21799_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_329_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14340_ _12340_/B _14274_/B _15171_/A vssd1 vssd1 vccd1 vccd1 _14340_/X sky130_fd_sc_hd__mux2_1
X_11552_ _20532_/B _11552_/B _11552_/C vssd1 vssd1 vccd1 vccd1 _20387_/A sky130_fd_sc_hd__nand3_4
X_23538_ _23538_/CLK _23538_/D vssd1 vssd1 vccd1 vccd1 _23538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_357_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11483_ _11483_/A vssd1 vssd1 vccd1 vccd1 _11483_/X sky130_fd_sc_hd__buf_6
X_14271_ _14290_/A vssd1 vssd1 vccd1 vccd1 _14310_/S sky130_fd_sc_hd__clkbuf_2
X_23469_ _23565_/CLK _23469_/D vssd1 vssd1 vccd1 vccd1 _23469_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16010_ _23004_/Q _16084_/A _16085_/A input233/X vssd1 vssd1 vccd1 vccd1 _22119_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_137_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13222_ _13218_/A _13219_/X _13221_/X _11537_/A vssd1 vssd1 vccd1 vccd1 _13222_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_353_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_341_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_325_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13153_ _23326_/Q _23294_/Q _23262_/Q _23550_/Q _11205_/A _13085_/X vssd1 vssd1 vccd1
+ vccd1 _13154_/B sky130_fd_sc_hd__mux4_1
XFILLER_151_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_312_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_345_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12104_ _22790_/Q _22758_/Q _22659_/Q _22726_/Q _12094_/X _11457_/B vssd1 vssd1 vccd1
+ vccd1 _12105_/B sky130_fd_sc_hd__mux4_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17961_ _22831_/Q _17950_/X _17960_/X _17948_/X vssd1 vssd1 vccd1 vccd1 _22831_/D
+ sky130_fd_sc_hd__o211a_1
X_13084_ _13084_/A vssd1 vssd1 vccd1 vccd1 _13149_/A sky130_fd_sc_hd__clkbuf_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12035_ _12949_/A _12034_/X _12721_/A vssd1 vssd1 vccd1 vccd1 _12035_/Y sky130_fd_sc_hd__o21ai_1
X_19700_ _19756_/A vssd1 vssd1 vccd1 vccd1 _19769_/S sky130_fd_sc_hd__buf_6
X_16912_ _16911_/X _22551_/Q _16915_/S vssd1 vssd1 vccd1 vccd1 _16913_/A sky130_fd_sc_hd__mux2_1
X_17892_ _18018_/A _18191_/A vssd1 vssd1 vccd1 vccd1 _17971_/A sky130_fd_sc_hd__nand2_1
XFILLER_266_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19631_ _19631_/A vssd1 vssd1 vccd1 vccd1 _23461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16843_ _16843_/A vssd1 vssd1 vccd1 vccd1 _22529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19562_ _23431_/Q _19172_/A _19566_/S vssd1 vssd1 vccd1 vccd1 _19563_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16774_ _16777_/A _16774_/B vssd1 vssd1 vccd1 vccd1 _16775_/A sky130_fd_sc_hd__or2_1
XFILLER_81_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13986_ _13986_/A vssd1 vssd1 vccd1 vccd1 _13986_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_281_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18513_ _23000_/Q _18518_/B vssd1 vssd1 vccd1 vccd1 _18513_/Y sky130_fd_sc_hd__nand2_1
XFILLER_234_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15725_ _15724_/X _14931_/A _14933_/A _22965_/Q vssd1 vssd1 vccd1 vccd1 _15725_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12937_ _12968_/A _12937_/B vssd1 vssd1 vccd1 vccd1 _12937_/Y sky130_fd_sc_hd__nor2_1
XFILLER_262_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19493_ _19493_/A vssd1 vssd1 vccd1 vccd1 _23400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18444_ _22976_/Q _18444_/B vssd1 vssd1 vccd1 vccd1 _18445_/B sky130_fd_sc_hd__and2_1
XFILLER_234_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15656_ _14755_/X _15643_/X _15655_/X vssd1 vssd1 vccd1 vccd1 _15656_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_179_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12868_ _12868_/A _13495_/A vssd1 vssd1 vccd1 vccd1 _13492_/A sky130_fd_sc_hd__nor2_1
XFILLER_222_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14607_ _23782_/Q _14605_/X _14606_/X vssd1 vssd1 vccd1 vccd1 _14607_/X sky130_fd_sc_hd__a21o_1
XFILLER_18_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18375_ _22951_/Q _22952_/Q _18375_/C vssd1 vssd1 vccd1 vccd1 _18377_/B sky130_fd_sc_hd__and3_1
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11819_ _11819_/A vssd1 vssd1 vccd1 vccd1 _11819_/X sky130_fd_sc_hd__buf_4
XFILLER_310_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15587_ _22930_/Q _14509_/X _14513_/X _22962_/Q vssd1 vssd1 vccd1 vccd1 _15587_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12799_ _12789_/Y _12791_/Y _12795_/Y _12798_/Y _11657_/X vssd1 vssd1 vccd1 vccd1
+ _12800_/C sky130_fd_sc_hd__o221a_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17326_ _17326_/A _17326_/B _17326_/C vssd1 vssd1 vccd1 vccd1 _17371_/A sky130_fd_sc_hd__and3_4
X_14538_ _23889_/Q vssd1 vssd1 vccd1 vccd1 _14538_/X sky130_fd_sc_hd__buf_4
XFILLER_174_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_336_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_335_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17257_ _22087_/A vssd1 vssd1 vccd1 vccd1 _22116_/A sky130_fd_sc_hd__clkbuf_16
X_14469_ _15729_/S vssd1 vssd1 vccd1 vccd1 _16171_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_317_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16208_ _16307_/S vssd1 vssd1 vccd1 vccd1 _16221_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17188_ _17167_/X _17179_/X _17187_/X _17176_/X vssd1 vssd1 vccd1 vccd1 _17188_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_316_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16139_ _23811_/Q _14916_/A _15067_/A vssd1 vssd1 vccd1 vccd1 _16139_/X sky130_fd_sc_hd__a21o_1
XFILLER_303_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_288_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_303_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_303_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19829_ _23550_/Q _19245_/A _19837_/S vssd1 vssd1 vccd1 vccd1 _19830_/A sky130_fd_sc_hd__mux2_1
XFILLER_257_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22840_ _22893_/CLK _22840_/D vssd1 vssd1 vccd1 vccd1 _22840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22771_ _23583_/CLK _22771_/D vssd1 vssd1 vccd1 vccd1 _22771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21722_ _21718_/Y _21719_/Y _21720_/X _21721_/X vssd1 vssd1 vccd1 vccd1 _21724_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_224_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21653_ _21653_/A _21653_/B _21653_/C vssd1 vssd1 vccd1 vccd1 _21689_/C sky130_fd_sc_hd__and3_1
XFILLER_40_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_339_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20604_ _20604_/A vssd1 vssd1 vccd1 vccd1 _20605_/A sky130_fd_sc_hd__inv_2
X_21584_ _21630_/A _23756_/Q vssd1 vssd1 vccd1 vccd1 _21585_/B sky130_fd_sc_hd__nand2_1
XFILLER_177_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23323_ _23547_/CLK _23323_/D vssd1 vssd1 vccd1 vccd1 _23323_/Q sky130_fd_sc_hd__dfxtp_1
X_20535_ _21093_/A _20535_/B vssd1 vssd1 vccd1 vccd1 _20779_/A sky130_fd_sc_hd__and2_1
XFILLER_166_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_326_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_308_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_354_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23254_ _23541_/CLK _23254_/D vssd1 vssd1 vccd1 vccd1 _23254_/Q sky130_fd_sc_hd__dfxtp_1
X_20466_ _20700_/A _20447_/X _20465_/X _20459_/X vssd1 vssd1 vccd1 vccd1 _23705_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_307_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22205_ _22205_/A _22205_/B vssd1 vssd1 vccd1 vccd1 _22206_/B sky130_fd_sc_hd__or2_1
XFILLER_341_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23185_ _23507_/CLK _23185_/D vssd1 vssd1 vccd1 vccd1 _23185_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_7315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20397_ _20320_/X _20395_/Y _20396_/X _22224_/A _20294_/X vssd1 vssd1 vccd1 vccd1
+ _20759_/A sky130_fd_sc_hd__a32o_4
XTAP_7326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22136_ _22136_/A _22136_/B vssd1 vssd1 vccd1 vccd1 _22137_/B sky130_fd_sc_hd__xnor2_1
XTAP_7359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_323_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_322_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_322_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput292 _14098_/X vssd1 vssd1 vccd1 vccd1 addr0[7] sky130_fd_sc_hd__buf_2
XTAP_6658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_288_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22067_ _22067_/A _22197_/B vssd1 vssd1 vccd1 vccd1 _22067_/Y sky130_fd_sc_hd__nor2_1
XTAP_6669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21018_ _21630_/A _21028_/B vssd1 vssd1 vccd1 vccd1 _21018_/X sky130_fd_sc_hd__or2_1
XTAP_5957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_331_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13840_ _13840_/A _13863_/B vssd1 vssd1 vccd1 vccd1 _13840_/Y sky130_fd_sc_hd__nor2_1
XFILLER_262_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_290_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13771_ _13875_/A _13771_/B vssd1 vssd1 vccd1 vccd1 _13771_/X sky130_fd_sc_hd__and2_1
XINSDIODE2_309 _18856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22969_ _22971_/CLK _22969_/D vssd1 vssd1 vccd1 vccd1 _22969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15510_ _23699_/Q _14905_/A _15509_/X vssd1 vssd1 vccd1 vccd1 _15510_/Y sky130_fd_sc_hd__o21ai_4
X_12722_ _12953_/A _12718_/X _12720_/X _12721_/X vssd1 vssd1 vccd1 vccd1 _12722_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16490_ _16490_/A vssd1 vssd1 vccd1 vccd1 _22402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15441_ _23602_/Q _15589_/A _15590_/A _23634_/Q vssd1 vssd1 vccd1 vccd1 _15441_/X
+ sky130_fd_sc_hd__o22a_2
X_12653_ _12047_/A _12652_/X _11598_/X vssd1 vssd1 vccd1 vccd1 _12653_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_188_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18160_ _18160_/A vssd1 vssd1 vccd1 vccd1 _22889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11604_ _12463_/A vssd1 vssd1 vccd1 vccd1 _12365_/A sky130_fd_sc_hd__clkbuf_4
X_15372_ _19201_/A vssd1 vssd1 vccd1 vccd1 _15372_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_358_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12584_ _12577_/X _12579_/X _12581_/X _12583_/X _11375_/A vssd1 vssd1 vccd1 vccd1
+ _12594_/B sky130_fd_sc_hd__a221o_1
XFILLER_357_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17111_ _22564_/Q _17091_/X _17083_/X _17110_/X vssd1 vssd1 vccd1 vccd1 _22564_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_184_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14323_ _14323_/A vssd1 vssd1 vccd1 vccd1 _14323_/Y sky130_fd_sc_hd__inv_2
X_18091_ _22868_/Q _18081_/X _18089_/X _18090_/X vssd1 vssd1 vccd1 vccd1 _22868_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_317_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11535_ _23426_/Q _23042_/Q _23394_/Q _23362_/Q _11532_/X _11544_/A vssd1 vssd1 vccd1
+ vccd1 _11536_/B sky130_fd_sc_hd__mux4_1
XFILLER_209_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17042_ _17042_/A vssd1 vssd1 vccd1 vccd1 _17042_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14254_ _15582_/B vssd1 vssd1 vccd1 vccd1 _14254_/X sky130_fd_sc_hd__buf_2
XFILLER_333_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11466_ _23491_/Q _23587_/Q _22551_/Q _22355_/Q _11461_/X _11462_/X vssd1 vssd1 vccd1
+ vccd1 _11466_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13205_ _23325_/Q _23293_/Q _23261_/Q _23549_/Q _11431_/A _13037_/A vssd1 vssd1 vccd1
+ vccd1 _13206_/B sky130_fd_sc_hd__mux4_2
XFILLER_332_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14185_ _23881_/Q vssd1 vssd1 vccd1 vccd1 _14196_/B sky130_fd_sc_hd__buf_6
XFILLER_171_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11397_ _23909_/Q vssd1 vssd1 vccd1 vccd1 _14175_/A sky130_fd_sc_hd__clkinv_2
XFILLER_174_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13136_ _16003_/A _20368_/A _13185_/S vssd1 vssd1 vccd1 vccd1 _13139_/B sky130_fd_sc_hd__mux2_1
XFILLER_98_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_297_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18993_ _16879_/X _23193_/Q _19001_/S vssd1 vssd1 vccd1 vccd1 _18994_/A sky130_fd_sc_hd__mux2_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17944_ _17944_/A _17987_/S vssd1 vssd1 vccd1 vccd1 _17944_/X sky130_fd_sc_hd__or2b_1
XFILLER_279_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13067_ _11353_/A _13060_/Y _13062_/Y _13064_/Y _13066_/Y vssd1 vssd1 vccd1 vccd1
+ _13067_/X sky130_fd_sc_hd__o32a_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_300_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12018_ _23315_/Q _23283_/Q _23251_/Q _23539_/Q _12008_/X _12734_/A vssd1 vssd1 vccd1
+ vccd1 _12019_/B sky130_fd_sc_hd__mux4_1
XFILLER_94_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17875_ _17875_/A vssd1 vssd1 vccd1 vccd1 _22808_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19614_ _19614_/A vssd1 vssd1 vccd1 vccd1 _23454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_254_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16826_ _16825_/X _22524_/Q _16829_/S vssd1 vssd1 vccd1 vccd1 _16827_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19545_ _19252_/X _23424_/Q _19549_/S vssd1 vssd1 vccd1 vccd1 _19546_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16757_ _16757_/A vssd1 vssd1 vccd1 vccd1 _22504_/D sky130_fd_sc_hd__clkbuf_1
X_13969_ _13969_/A vssd1 vssd1 vccd1 vccd1 _13979_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15708_ _15706_/X _21888_/B _15708_/S vssd1 vssd1 vccd1 vccd1 _18830_/A sky130_fd_sc_hd__mux2_8
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19476_ _19476_/A vssd1 vssd1 vccd1 vccd1 _23393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_262_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16688_ _16783_/A vssd1 vssd1 vccd1 vccd1 _16729_/A sky130_fd_sc_hd__buf_6
XFILLER_61_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18427_ _18427_/A _22970_/Q _18427_/C vssd1 vssd1 vccd1 vccd1 _18429_/B sky130_fd_sc_hd__and3_1
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ _13532_/A _14674_/X _15638_/X vssd1 vssd1 vccd1 vccd1 _15639_/X sky130_fd_sc_hd__a21o_2
XFILLER_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18358_ _18358_/A _18358_/B _18359_/B vssd1 vssd1 vccd1 vccd1 _22946_/D sky130_fd_sc_hd__nor3_1
XFILLER_203_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17309_ _21079_/B _17308_/X _17317_/S vssd1 vssd1 vccd1 vccd1 _17309_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18289_ _18298_/D vssd1 vssd1 vccd1 vccd1 _18296_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_175_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20320_ _20320_/A vssd1 vssd1 vccd1 vccd1 _20320_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_336_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_317_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20251_ _20187_/X _20249_/X _20250_/Y _21641_/A _20200_/X vssd1 vssd1 vccd1 vccd1
+ _20630_/A sky130_fd_sc_hd__a32o_4
XFILLER_351_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20182_ _20147_/X _21351_/B _20181_/X vssd1 vssd1 vccd1 vccd1 _20570_/A sky130_fd_sc_hd__o21ai_4
XFILLER_277_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_320_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23941_ _23942_/CLK _23941_/D vssd1 vssd1 vccd1 vccd1 _23941_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23872_ _23876_/CLK _23872_/D vssd1 vssd1 vccd1 vccd1 _23872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_272_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22823_ _22830_/CLK _22823_/D vssd1 vssd1 vccd1 vccd1 _22823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22754_ _23054_/CLK _22754_/D vssd1 vssd1 vccd1 vccd1 _22754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_358_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21705_ _21705_/A _21705_/B vssd1 vssd1 vccd1 vccd1 _21705_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22685_ _23564_/CLK _22685_/D vssd1 vssd1 vccd1 vccd1 _22685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_338_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_358_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21636_ _21636_/A _21641_/A vssd1 vssd1 vccd1 vccd1 _21637_/B sky130_fd_sc_hd__or2_1
XFILLER_339_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21567_ _22025_/A _21567_/B vssd1 vssd1 vccd1 vccd1 _21567_/Y sky130_fd_sc_hd__nand2_1
XFILLER_355_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11320_ _11320_/A vssd1 vssd1 vccd1 vccd1 _11533_/A sky130_fd_sc_hd__buf_2
X_23306_ _23466_/CLK _23306_/D vssd1 vssd1 vccd1 vccd1 _23306_/Q sky130_fd_sc_hd__dfxtp_1
X_20518_ _23715_/Q _20523_/B _20518_/C vssd1 vssd1 vccd1 vccd1 _20520_/C sky130_fd_sc_hd__and3_1
XFILLER_138_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_315_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21498_ _23819_/Q _21496_/Y _22083_/A vssd1 vssd1 vccd1 vccd1 _21498_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_314_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11251_ _23882_/Q _23881_/Q _14814_/C vssd1 vssd1 vccd1 vccd1 _11382_/C sky130_fd_sc_hd__and3b_1
XFILLER_326_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20449_ _20654_/A _20447_/X _20448_/X _20445_/X vssd1 vssd1 vccd1 vccd1 _23698_/D
+ sky130_fd_sc_hd__o211a_1
X_23237_ _23525_/CLK _23237_/D vssd1 vssd1 vccd1 vccd1 _23237_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_7101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11182_ _13158_/A vssd1 vssd1 vccd1 vccd1 _13051_/A sky130_fd_sc_hd__buf_4
XFILLER_134_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23168_ _23264_/CLK _23168_/D vssd1 vssd1 vccd1 vccd1 _23168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22119_ _22119_/A _22224_/B vssd1 vssd1 vccd1 vccd1 _22119_/Y sky130_fd_sc_hd__nor2_1
XTAP_7189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23099_ _23515_/CLK _23099_/D vssd1 vssd1 vccd1 vccd1 _23099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_294_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15990_ _23711_/Q _15592_/X _15989_/X vssd1 vssd1 vccd1 vccd1 _15990_/Y sky130_fd_sc_hd__o21ai_4
XTAP_6455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14941_ _13906_/Y _14940_/B _14940_/Y _14682_/X vssd1 vssd1 vccd1 vccd1 _14941_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17660_ _19555_/B _17804_/B vssd1 vssd1 vccd1 vccd1 _17717_/A sky130_fd_sc_hd__nor2_8
XFILLER_75_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14872_ _23784_/Q _14605_/X _14486_/X vssd1 vssd1 vccd1 vccd1 _14872_/X sky130_fd_sc_hd__a21o_1
XFILLER_275_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16611_ _16611_/A vssd1 vssd1 vccd1 vccd1 _22454_/D sky130_fd_sc_hd__clkbuf_1
X_13823_ _13861_/A _14052_/C vssd1 vssd1 vccd1 vccd1 _13823_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17591_ _18817_/A vssd1 vssd1 vccd1 vccd1 _17591_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_106 _21601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19330_ _19330_/A vssd1 vssd1 vccd1 vccd1 _23328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16542_ _14811_/X _22424_/Q _16546_/S vssd1 vssd1 vccd1 vccd1 _16543_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_117 _20217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_128 _14292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13754_ _13974_/B _13754_/B vssd1 vssd1 vccd1 vccd1 _13754_/Y sky130_fd_sc_hd__nor2_1
XINSDIODE2_139 _13022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12705_ _11277_/A _12667_/X _11402_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _12742_/A
+ sky130_fd_sc_hd__a22o_4
X_19261_ _19261_/A vssd1 vssd1 vccd1 vccd1 _19261_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_349_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16473_ _16473_/A vssd1 vssd1 vccd1 vccd1 _22394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13685_ _14072_/B vssd1 vssd1 vccd1 vccd1 _13715_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_232_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18212_ _22897_/Q _18214_/B vssd1 vssd1 vccd1 vccd1 _18212_/X sky130_fd_sc_hd__or2_1
XFILLER_204_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15424_ _15424_/A vssd1 vssd1 vccd1 vccd1 _22273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_349_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12636_ _12636_/A vssd1 vssd1 vccd1 vccd1 _12636_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19192_ _19191_/X _23277_/Q _19195_/S vssd1 vssd1 vccd1 vccd1 _19193_/A sky130_fd_sc_hd__mux2_1
XPHY_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18143_ _18172_/A vssd1 vssd1 vccd1 vccd1 _18144_/B sky130_fd_sc_hd__clkbuf_2
XPHY_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15355_ _23792_/Q _14605_/X _14486_/X vssd1 vssd1 vccd1 vccd1 _15355_/X sky130_fd_sc_hd__a21o_1
X_12567_ _12567_/A _12567_/B vssd1 vssd1 vccd1 vccd1 _12567_/X sky130_fd_sc_hd__or2_1
XFILLER_345_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14306_ _14304_/X _14305_/X _14369_/A vssd1 vssd1 vccd1 vccd1 _14306_/X sky130_fd_sc_hd__mux2_1
X_18074_ _22862_/Q _18067_/X _18068_/X _22995_/Q _18069_/X vssd1 vssd1 vccd1 vccd1
+ _18074_/X sky130_fd_sc_hd__a221o_1
X_11518_ _11533_/A vssd1 vssd1 vccd1 vccd1 _11519_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_356_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_333_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15286_ _15286_/A _15433_/B vssd1 vssd1 vccd1 vccd1 _15675_/B sky130_fd_sc_hd__nand2_1
XFILLER_184_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_305_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12498_ _11561_/A _11404_/B _12520_/S vssd1 vssd1 vccd1 vccd1 _12546_/A sky130_fd_sc_hd__o21ai_1
XFILLER_345_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17025_ _13454_/Y _17648_/B _16947_/X _17021_/X _17024_/X vssd1 vssd1 vccd1 vccd1
+ _17025_/X sky130_fd_sc_hd__a311o_1
XFILLER_236_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14237_ _22503_/Q _14232_/X _13888_/B _14236_/X vssd1 vssd1 vccd1 vccd1 _15186_/A
+ sky130_fd_sc_hd__o211ai_2
X_11449_ _11236_/A _11446_/X _11448_/X _11247_/A vssd1 vssd1 vccd1 vccd1 _11449_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_291_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14168_ _20533_/C _14128_/Y _14133_/X _14167_/X vssd1 vssd1 vccd1 vccd1 _14609_/A
+ sky130_fd_sc_hd__o31a_4
XFILLER_301_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_341_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_286_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13119_ _13180_/A _13119_/B vssd1 vssd1 vccd1 vccd1 _13119_/Y sky130_fd_sc_hd__nor2_1
XFILLER_298_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_302_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18976_ _18976_/A vssd1 vssd1 vccd1 vccd1 _23185_/D sky130_fd_sc_hd__clkbuf_1
X_14099_ _14099_/A vssd1 vssd1 vccd1 vccd1 _14099_/Y sky130_fd_sc_hd__inv_2
XFILLER_286_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17927_ _22820_/Q _17922_/X _17896_/X _17926_/X _17915_/X vssd1 vssd1 vccd1 vccd1
+ _17927_/X sky130_fd_sc_hd__a221o_1
XFILLER_285_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_294_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17858_ _17858_/A vssd1 vssd1 vccd1 vccd1 _22800_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16809_ _16809_/A vssd1 vssd1 vccd1 vccd1 _22519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17789_ _17789_/A vssd1 vssd1 vccd1 vccd1 _17798_/S sky130_fd_sc_hd__buf_6
XFILLER_214_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19528_ _19528_/A vssd1 vssd1 vccd1 vccd1 _23416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19459_ _19459_/A vssd1 vssd1 vccd1 vccd1 _23385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_328_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22470_ _23575_/CLK _22470_/D vssd1 vssd1 vccd1 vccd1 _22470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_349_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21421_ _21520_/A _21421_/B vssd1 vssd1 vccd1 vccd1 _21421_/Y sky130_fd_sc_hd__nor2_1
XFILLER_348_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21352_ _21403_/A _21352_/B vssd1 vssd1 vccd1 vccd1 _21353_/B sky130_fd_sc_hd__nor2_1
XFILLER_163_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20303_ _20303_/A _20340_/B vssd1 vssd1 vccd1 vccd1 _20306_/B sky130_fd_sc_hd__or2_1
XFILLER_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21283_ _21283_/A _21283_/B vssd1 vssd1 vccd1 vccd1 _21283_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23022_ _23502_/CLK _23022_/D vssd1 vssd1 vccd1 vccd1 _23022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20234_ _20234_/A _20340_/B vssd1 vssd1 vccd1 vccd1 _20236_/B sky130_fd_sc_hd__nor2_1
XFILLER_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20165_ _20379_/A vssd1 vssd1 vccd1 vccd1 _20165_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_320_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20096_ _20120_/A _20096_/B _20110_/C vssd1 vssd1 vccd1 vccd1 _23639_/D sky130_fd_sc_hd__nor3_1
XFILLER_292_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23924_ _23926_/CLK _23924_/D vssd1 vssd1 vccd1 vccd1 _23924_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_291_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23855_ _23856_/CLK _23855_/D vssd1 vssd1 vccd1 vccd1 _23855_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6_1_wb_clk_i clkbuf_3_6_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_1_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22806_ _23585_/CLK _22806_/D vssd1 vssd1 vccd1 vccd1 _22806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23786_ _23862_/CLK _23786_/D vssd1 vssd1 vccd1 vccd1 _23786_/Q sky130_fd_sc_hd__dfxtp_4
X_20998_ _23814_/Q _20993_/X _20996_/Y _20997_/X vssd1 vssd1 vccd1 vccd1 _23814_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_225_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_98_wb_clk_i _22899_/CLK vssd1 vssd1 vccd1 vccd1 _23426_/CLK sky130_fd_sc_hd__clkbuf_16
X_22737_ _23451_/CLK _22737_/D vssd1 vssd1 vccd1 vccd1 _22737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_347_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13470_ _13470_/A _21335_/C vssd1 vssd1 vccd1 vccd1 _13470_/X sky130_fd_sc_hd__or2_4
XFILLER_125_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23895_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22668_ _22801_/CLK _22668_/D vssd1 vssd1 vccd1 vccd1 _22668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_346_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_329_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12421_ _12421_/A _12421_/B vssd1 vssd1 vccd1 vccd1 _12421_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21619_ _21636_/A _21619_/B vssd1 vssd1 vccd1 vccd1 _21619_/X sky130_fd_sc_hd__and2_1
X_22599_ _22600_/CLK _22599_/D vssd1 vssd1 vccd1 vccd1 _22599_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_337_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15140_ _22921_/Q _15259_/B vssd1 vssd1 vccd1 vccd1 _15140_/X sky130_fd_sc_hd__and2_1
XFILLER_343_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12352_ _11138_/A _12351_/X _11780_/A vssd1 vssd1 vccd1 vccd1 _12352_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_126_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_299_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11303_ _12324_/A vssd1 vssd1 vccd1 vccd1 _11821_/A sky130_fd_sc_hd__clkbuf_4
X_15071_ _23659_/Q _15067_/X _15068_/X _15070_/X _15593_/A vssd1 vssd1 vccd1 vccd1
+ _15071_/X sky130_fd_sc_hd__a221o_2
X_12283_ _23917_/Q _12283_/B vssd1 vssd1 vccd1 vccd1 _12283_/X sky130_fd_sc_hd__or2_1
X_14022_ input244/X _14004_/X _14021_/X vssd1 vssd1 vccd1 vccd1 _14022_/X sky130_fd_sc_hd__a21o_4
X_11234_ _12816_/A vssd1 vssd1 vccd1 vccd1 _11235_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_296_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18830_ _18830_/A vssd1 vssd1 vccd1 vccd1 _18830_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_268_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11165_ _12685_/A vssd1 vssd1 vccd1 vccd1 _11166_/A sky130_fd_sc_hd__buf_4
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_353_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_310_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18761_ _16905_/X _23105_/Q _18763_/S vssd1 vssd1 vccd1 vccd1 _18762_/A sky130_fd_sc_hd__mux2_1
X_15973_ _15968_/X _15970_/Y _22116_/B _15321_/X vssd1 vssd1 vccd1 vccd1 _18852_/A
+ sky130_fd_sc_hd__a2bb2o_4
X_11096_ _13459_/A vssd1 vssd1 vccd1 vccd1 _13472_/B sky130_fd_sc_hd__inv_2
XTAP_6285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17712_ _17712_/A vssd1 vssd1 vccd1 vccd1 _22735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14924_ _23817_/Q _14907_/X _14909_/X _14921_/X _14923_/X vssd1 vssd1 vccd1 vccd1
+ _14924_/X sky130_fd_sc_hd__a221o_4
XFILLER_282_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18692_ _18692_/A vssd1 vssd1 vccd1 vccd1 _23074_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17643_ _22708_/Q _17642_/X _17646_/S vssd1 vssd1 vccd1 vccd1 _17644_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14855_ _14855_/A _14855_/B vssd1 vssd1 vccd1 vccd1 _14855_/X sky130_fd_sc_hd__or2_1
XFILLER_251_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_291_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13806_ _13790_/X _13852_/A _13804_/Y _13851_/A vssd1 vssd1 vccd1 vccd1 _14046_/C
+ sky130_fd_sc_hd__a211o_4
XFILLER_91_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17574_ _17574_/A vssd1 vssd1 vccd1 vccd1 _22686_/D sky130_fd_sc_hd__clkbuf_1
X_14786_ _14345_/X _14319_/X _14845_/S vssd1 vssd1 vccd1 vccd1 _15086_/A sky130_fd_sc_hd__mux2_2
X_11998_ _12024_/A vssd1 vssd1 vccd1 vccd1 _12733_/A sky130_fd_sc_hd__buf_6
XFILLER_205_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_323_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19313_ _19324_/A vssd1 vssd1 vccd1 vccd1 _19322_/S sky130_fd_sc_hd__clkbuf_4
X_16525_ _16525_/A vssd1 vssd1 vccd1 vccd1 _22418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13737_ _13737_/A vssd1 vssd1 vccd1 vccd1 _13738_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_189_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19244_ _19244_/A vssd1 vssd1 vccd1 vccd1 _23293_/D sky130_fd_sc_hd__clkbuf_1
X_16456_ _16456_/A vssd1 vssd1 vccd1 vccd1 _22388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_319_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13668_ _22612_/Q vssd1 vssd1 vccd1 vccd1 _16927_/A sky130_fd_sc_hd__buf_2
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15407_ _14516_/A _15394_/X _15406_/X vssd1 vssd1 vccd1 vccd1 _15408_/A sky130_fd_sc_hd__o21ai_4
X_12619_ _12780_/A vssd1 vssd1 vccd1 vccd1 _12958_/A sky130_fd_sc_hd__buf_2
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19175_ _19175_/A vssd1 vssd1 vccd1 vccd1 _19175_/X sky130_fd_sc_hd__clkbuf_2
X_16387_ _16455_/S vssd1 vssd1 vccd1 vccd1 _16396_/S sky130_fd_sc_hd__buf_8
X_13599_ _13599_/A _13599_/B vssd1 vssd1 vccd1 vccd1 _13599_/X sky130_fd_sc_hd__xor2_4
XFILLER_318_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18126_ _14119_/C _22879_/Q _18126_/S vssd1 vssd1 vccd1 vccd1 _18126_/X sky130_fd_sc_hd__mux2_1
XFILLER_352_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15338_ _15338_/A _15338_/B vssd1 vssd1 vccd1 vccd1 _15338_/X sky130_fd_sc_hd__or2_2
XFILLER_200_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_334_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18057_ hold4/A _18052_/X _18053_/X _22989_/Q _18054_/X vssd1 vssd1 vccd1 vccd1 _18057_/X
+ sky130_fd_sc_hd__a221o_1
X_15269_ _22955_/Q _15268_/X _16028_/A vssd1 vssd1 vccd1 vccd1 _15269_/X sky130_fd_sc_hd__mux2_1
X_17008_ _23463_/Q _16987_/X _16988_/X _16989_/X _14756_/X vssd1 vssd1 vccd1 vccd1
+ _17008_/X sky130_fd_sc_hd__a32o_1
XFILLER_299_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_299_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_286_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18959_ _19016_/S vssd1 vssd1 vccd1 vccd1 _18968_/S sky130_fd_sc_hd__buf_4
XFILLER_6_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21970_ _23834_/Q _23768_/Q vssd1 vssd1 vccd1 vccd1 _21971_/B sky130_fd_sc_hd__nor2_1
XFILLER_239_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20921_ _23789_/Q _20911_/X _20919_/X _20920_/X vssd1 vssd1 vccd1 vccd1 _23789_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_255_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23640_ _23643_/CLK _23640_/D vssd1 vssd1 vccd1 vccd1 _23640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20852_ _20861_/A _20852_/B vssd1 vssd1 vccd1 vccd1 _20853_/A sky130_fd_sc_hd__and2_1
XFILLER_81_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23571_ _23571_/CLK _23571_/D vssd1 vssd1 vccd1 vccd1 _23571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20783_ _23751_/Q _20786_/B _20782_/X _20763_/X vssd1 vssd1 vccd1 vccd1 _23751_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_223_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_470 _15671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_481 _19969_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22522_ _23558_/CLK _22522_/D vssd1 vssd1 vccd1 vccd1 _22522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_329_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_328_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_492 _13651_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22453_ _23556_/CLK _22453_/D vssd1 vssd1 vccd1 vccd1 _22453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21404_ _21404_/A _21404_/B vssd1 vssd1 vccd1 vccd1 _21404_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_136_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22384_ _23584_/CLK _22384_/D vssd1 vssd1 vccd1 vccd1 _22384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21335_ _21335_/A _21335_/B _21335_/C vssd1 vssd1 vccd1 vccd1 _21336_/B sky130_fd_sc_hd__and3_2
XFILLER_108_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_145_wb_clk_i _22899_/CLK vssd1 vssd1 vccd1 vccd1 _22908_/CLK sky130_fd_sc_hd__clkbuf_16
X_21266_ _15864_/X _21196_/X _21265_/X vssd1 vssd1 vccd1 vccd1 _23902_/D sky130_fd_sc_hd__o21ba_2
XFILLER_89_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23005_ _23005_/CLK _23005_/D vssd1 vssd1 vccd1 vccd1 _23005_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20217_ _20217_/A _20279_/B vssd1 vssd1 vccd1 vccd1 _20217_/Y sky130_fd_sc_hd__nand2_1
XFILLER_235_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21197_ _21260_/S vssd1 vssd1 vccd1 vccd1 _21243_/A sky130_fd_sc_hd__buf_2
XFILLER_289_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20148_ _20148_/A vssd1 vssd1 vccd1 vccd1 _20250_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_320_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20079_ _23632_/Q _20079_/B _20079_/C _20085_/D vssd1 vssd1 vccd1 vccd1 _20090_/D
+ sky130_fd_sc_hd__and4_1
X_12970_ _12926_/A _12969_/X _11233_/A vssd1 vssd1 vccd1 vccd1 _12970_/Y sky130_fd_sc_hd__o21ai_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23907_ _23907_/CLK _23907_/D vssd1 vssd1 vccd1 vccd1 _23907_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _22462_/Q _22622_/Q _22301_/Q _23437_/Q _11920_/X _11652_/A vssd1 vssd1 vccd1
+ vccd1 _11922_/B sky130_fd_sc_hd__mux4_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _14637_/X _14638_/X _14853_/S vssd1 vssd1 vccd1 vccd1 _14640_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23838_ _23841_/CLK _23838_/D vssd1 vssd1 vccd1 vccd1 _23838_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11852_ _22270_/Q _23086_/Q _23502_/Q _22431_/Q _11595_/A _11621_/A vssd1 vssd1 vccd1
+ vccd1 _11853_/B sky130_fd_sc_hd__mux4_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ input133/X input118/X _15033_/S vssd1 vssd1 vccd1 vccd1 _14571_/X sky130_fd_sc_hd__mux2_8
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11783_ _12371_/A _11772_/Y _11774_/Y _11782_/X _11216_/A vssd1 vssd1 vccd1 vccd1
+ _11793_/B sky130_fd_sc_hd__o311a_1
X_23769_ _23776_/CLK _23769_/D vssd1 vssd1 vccd1 vccd1 _23769_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16310_ _16310_/A _16457_/B vssd1 vssd1 vccd1 vccd1 _19771_/A sky130_fd_sc_hd__or2b_4
XFILLER_82_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13522_ _13522_/A vssd1 vssd1 vccd1 vccd1 _13525_/A sky130_fd_sc_hd__inv_2
XFILLER_242_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17290_ _23489_/Q _17016_/X _17017_/X _17268_/X _17289_/Y vssd1 vssd1 vccd1 vccd1
+ _17290_/X sky130_fd_sc_hd__a32o_1
XFILLER_186_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16241_ _22303_/Q _16239_/X _16253_/S vssd1 vssd1 vccd1 vccd1 _16242_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13453_ _21079_/B _14175_/B _20533_/B _21285_/A vssd1 vssd1 vccd1 vccd1 _13455_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12404_ _12397_/Y _12399_/Y _12401_/Y _12403_/Y _11273_/A vssd1 vssd1 vccd1 vccd1
+ _12414_/B sky130_fd_sc_hd__o221a_1
XFILLER_127_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_316_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16172_ _23812_/Q _14916_/A _15067_/A vssd1 vssd1 vccd1 vccd1 _16172_/X sky130_fd_sc_hd__a21o_1
XFILLER_356_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13384_ _12159_/A _12163_/Y _13345_/X vssd1 vssd1 vccd1 vccd1 _13385_/B sky130_fd_sc_hd__a21oi_1
XFILLER_315_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15123_ _15123_/A _15335_/B vssd1 vssd1 vccd1 vccd1 _15123_/Y sky130_fd_sc_hd__nor2_1
X_12335_ _12316_/A _12332_/X _12334_/X _11679_/A vssd1 vssd1 vccd1 vccd1 _12335_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_343_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_315_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_330_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19931_ _19934_/B _19934_/C _19930_/Y vssd1 vssd1 vccd1 vccd1 _23594_/D sky130_fd_sc_hd__o21a_1
X_15054_ input165/X input130/X _15114_/S vssd1 vssd1 vccd1 vccd1 _15054_/X sky130_fd_sc_hd__mux2_8
XFILLER_147_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12266_ _12406_/A _12265_/X _11347_/A vssd1 vssd1 vccd1 vccd1 _12266_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_324_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_342_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14005_ _14072_/C vssd1 vssd1 vccd1 vccd1 _14036_/B sky130_fd_sc_hd__clkbuf_1
X_11217_ _11217_/A vssd1 vssd1 vccd1 vccd1 _11218_/A sky130_fd_sc_hd__buf_4
X_19862_ _19862_/A vssd1 vssd1 vccd1 vccd1 _23564_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_268_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12197_ _23468_/Q _23564_/Q _22528_/Q _22332_/Q _11148_/A _11840_/X vssd1 vssd1 vccd1
+ vccd1 _12197_/X sky130_fd_sc_hd__mux4_2
XFILLER_122_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18813_ _18813_/A vssd1 vssd1 vccd1 vccd1 _23121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11148_ _11148_/A vssd1 vssd1 vccd1 vccd1 _11770_/A sky130_fd_sc_hd__buf_4
XTAP_6071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19793_ _23534_/Q _19194_/A _19793_/S vssd1 vssd1 vccd1 vccd1 _19794_/A sky130_fd_sc_hd__mux2_1
XTAP_6082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18744_ _16879_/X _23097_/Q _18752_/S vssd1 vssd1 vccd1 vccd1 _18745_/A sky130_fd_sc_hd__mux2_1
XFILLER_283_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11079_ _23893_/Q vssd1 vssd1 vccd1 vccd1 _11080_/A sky130_fd_sc_hd__inv_2
X_15956_ _23806_/Q _14742_/X _14606_/A vssd1 vssd1 vccd1 vccd1 _15956_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput170 dout1[9] vssd1 vssd1 vccd1 vccd1 input170/X sky130_fd_sc_hd__clkbuf_1
XFILLER_255_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput181 irq[4] vssd1 vssd1 vccd1 vccd1 _20508_/C sky130_fd_sc_hd__buf_2
Xinput192 localMemory_wb_adr_i[11] vssd1 vssd1 vccd1 vccd1 input192/X sky130_fd_sc_hd__clkbuf_1
X_14907_ _14907_/A vssd1 vssd1 vccd1 vccd1 _14907_/X sky130_fd_sc_hd__buf_2
XFILLER_292_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15887_ _15003_/X _15874_/X _15886_/X vssd1 vssd1 vccd1 vccd1 _17232_/A sky130_fd_sc_hd__o21ai_4
XFILLER_236_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18675_ _18675_/A vssd1 vssd1 vccd1 vccd1 _23066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17626_ _18852_/A vssd1 vssd1 vccd1 vccd1 _17626_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14838_ _13508_/Y _14254_/X _14761_/X _13503_/Y _14837_/X vssd1 vssd1 vccd1 vccd1
+ _14838_/X sky130_fd_sc_hd__a221o_1
XFILLER_252_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17557_ _22681_/Q _17556_/X _17560_/S vssd1 vssd1 vccd1 vccd1 _17558_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14769_ _15341_/S _14768_/Y _14630_/X vssd1 vssd1 vccd1 vccd1 _16097_/B sky130_fd_sc_hd__a21o_1
XFILLER_205_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16508_ _16508_/A vssd1 vssd1 vccd1 vccd1 _22410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17488_ _22652_/Q _16227_/X _17494_/S vssd1 vssd1 vccd1 vccd1 _17489_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19227_ _19226_/X _23288_/Q _19227_/S vssd1 vssd1 vccd1 vccd1 _19228_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16439_ _16439_/A vssd1 vssd1 vccd1 vccd1 _22380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19158_ _19158_/A vssd1 vssd1 vccd1 vccd1 _23266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18109_ _22874_/Q _18097_/X _18098_/X _23007_/Q _18099_/X vssd1 vssd1 vccd1 vccd1
+ _18109_/X sky130_fd_sc_hd__a221o_1
XFILLER_258_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19089_ _19089_/A vssd1 vssd1 vccd1 vccd1 _23236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_306_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_333_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21120_ _23856_/Q _21110_/X _21111_/X _20623_/A vssd1 vssd1 vccd1 vccd1 _21121_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_322_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21051_ _21051_/A vssd1 vssd1 vccd1 vccd1 _21068_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_259_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20002_ _23610_/Q _23609_/Q vssd1 vssd1 vccd1 vccd1 _20005_/D sky130_fd_sc_hd__and2_1
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_330_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21953_ _21953_/A _21953_/B vssd1 vssd1 vccd1 vccd1 _21953_/X sky130_fd_sc_hd__xor2_1
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20904_ _23914_/Q vssd1 vssd1 vccd1 vccd1 _21400_/A sky130_fd_sc_hd__buf_6
XFILLER_282_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21884_ _21884_/A _21883_/Y vssd1 vssd1 vccd1 vccd1 _21885_/B sky130_fd_sc_hd__or2b_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23623_ _23634_/CLK _23623_/D vssd1 vssd1 vccd1 vccd1 _23623_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20835_ _20835_/A vssd1 vssd1 vccd1 vccd1 _23764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23554_ _23554_/CLK _23554_/D vssd1 vssd1 vccd1 vccd1 _23554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20766_ _21079_/A _20564_/X _20733_/X vssd1 vssd1 vccd1 vccd1 _20766_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_168_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22505_ _23684_/CLK _22505_/D vssd1 vssd1 vccd1 vccd1 _22505_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_356_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23485_ _23547_/CLK _23485_/D vssd1 vssd1 vccd1 vccd1 _23485_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_156_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20697_ _20729_/A vssd1 vssd1 vccd1 vccd1 _20697_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_356_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22436_ _23505_/CLK _22436_/D vssd1 vssd1 vccd1 vccd1 _22436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_338_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22367_ _23567_/CLK _22367_/D vssd1 vssd1 vccd1 vccd1 _22367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12120_ _22305_/Q _23441_/Q _12120_/S vssd1 vssd1 vccd1 vccd1 _12120_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21318_ _21318_/A _21318_/B vssd1 vssd1 vccd1 vccd1 _21319_/B sky130_fd_sc_hd__nand2_1
XFILLER_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22298_ _23564_/CLK _22298_/D vssd1 vssd1 vccd1 vccd1 _22298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_324_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12051_ _23315_/Q _23283_/Q _23251_/Q _23539_/Q _11972_/X _12756_/A vssd1 vssd1 vccd1
+ vccd1 _12052_/B sky130_fd_sc_hd__mux4_1
XFILLER_278_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21249_ _17172_/A _15634_/X _21257_/S vssd1 vssd1 vccd1 vccd1 _21250_/B sky130_fd_sc_hd__mux2_1
XFILLER_117_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15810_ _23706_/Q _15210_/A _15809_/X vssd1 vssd1 vccd1 vccd1 _15810_/X sky130_fd_sc_hd__o21a_2
X_16790_ _16790_/A vssd1 vssd1 vccd1 vccd1 _22513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_350_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15741_ _14822_/A _15717_/X _15740_/X vssd1 vssd1 vccd1 vccd1 _15741_/Y sky130_fd_sc_hd__a21oi_2
X_12953_ _12953_/A _12953_/B vssd1 vssd1 vccd1 vccd1 _12953_/X sky130_fd_sc_hd__or2_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ _22269_/Q _23085_/Q _23501_/Q _22430_/Q _12070_/S _11613_/A vssd1 vssd1 vccd1
+ vccd1 _11905_/B sky130_fd_sc_hd__mux4_1
X_18460_ _22980_/Q _18465_/B vssd1 vssd1 vccd1 vccd1 _18460_/Y sky130_fd_sc_hd__nand2_1
XFILLER_261_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_42_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23570_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15672_ _15672_/A vssd1 vssd1 vccd1 vccd1 _15672_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _12871_/A _12883_/X _11132_/A vssd1 vssd1 vccd1 vccd1 _12884_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_245_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17411_ _17411_/A vssd1 vssd1 vccd1 vccd1 _22618_/D sky130_fd_sc_hd__clkbuf_1
X_14623_ _15387_/S vssd1 vssd1 vccd1 vccd1 _15292_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18391_ _15351_/A _18392_/C _22958_/Q vssd1 vssd1 vccd1 vccd1 _18393_/B sky130_fd_sc_hd__a21oi_1
XFILLER_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11835_ _12556_/A vssd1 vssd1 vccd1 vccd1 _12554_/S sky130_fd_sc_hd__buf_4
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17342_/A vssd1 vssd1 vccd1 vccd1 _22592_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14554_ _23946_/Q vssd1 vssd1 vccd1 vccd1 _21677_/A sky130_fd_sc_hd__buf_2
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _13337_/A vssd1 vssd1 vccd1 vccd1 _13343_/B sky130_fd_sc_hd__inv_2
XFILLER_202_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13505_ _13505_/A _13506_/B vssd1 vssd1 vccd1 vccd1 _13505_/X sky130_fd_sc_hd__or2_2
X_17273_ _17245_/X _17272_/X _17262_/X _17215_/X vssd1 vssd1 vccd1 vccd1 _17273_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_9_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14485_ _15067_/A vssd1 vssd1 vccd1 vccd1 _14606_/A sky130_fd_sc_hd__clkbuf_4
X_11697_ _23216_/Q _23184_/Q _23152_/Q _23120_/Q _11574_/A _11696_/X vssd1 vssd1 vccd1
+ vccd1 _11698_/B sky130_fd_sc_hd__mux4_1
XFILLER_202_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19012_ _16908_/X _23202_/Q _19012_/S vssd1 vssd1 vccd1 vccd1 _19013_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16224_ _16307_/S vssd1 vssd1 vccd1 vccd1 _16237_/S sky130_fd_sc_hd__buf_4
XFILLER_201_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13436_ _13436_/A _14250_/A vssd1 vssd1 vccd1 vccd1 _14177_/A sky130_fd_sc_hd__nand2_1
XFILLER_127_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_316_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16155_ _15752_/X _16148_/X _16154_/Y _16005_/X vssd1 vssd1 vccd1 vccd1 _16155_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13367_ _13367_/A _14759_/A _13367_/C _13367_/D vssd1 vssd1 vccd1 vccd1 _13370_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ _15106_/A vssd1 vssd1 vccd1 vccd1 _22267_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12318_ _12318_/A _12318_/B vssd1 vssd1 vccd1 vccd1 _12318_/X sky130_fd_sc_hd__or2_1
XFILLER_316_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16086_ _23006_/Q _16944_/A _16085_/X input235/X vssd1 vssd1 vccd1 vccd1 _22171_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_182_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_343_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_308_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_303_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13298_ _13319_/B vssd1 vssd1 vccd1 vccd1 _13300_/B sky130_fd_sc_hd__inv_2
XFILLER_330_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19914_ _19914_/A vssd1 vssd1 vccd1 vccd1 _23588_/D sky130_fd_sc_hd__clkbuf_1
X_15037_ _15037_/A _15049_/C vssd1 vssd1 vccd1 vccd1 _21442_/B sky130_fd_sc_hd__xnor2_1
XFILLER_130_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12249_ _12196_/X _12243_/Y _12246_/Y _12248_/Y vssd1 vssd1 vccd1 vccd1 _12249_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_69_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19845_ _19913_/S vssd1 vssd1 vccd1 vccd1 _19854_/S sky130_fd_sc_hd__buf_4
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_288_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19776_ _23526_/Q _19169_/A _19782_/S vssd1 vssd1 vccd1 vccd1 _19777_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16988_ _17231_/A vssd1 vssd1 vccd1 vccd1 _16988_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18727_ _18727_/A vssd1 vssd1 vccd1 vccd1 _23089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15939_ _22087_/A _15940_/B vssd1 vssd1 vccd1 vccd1 _16039_/C sky130_fd_sc_hd__and2_2
XFILLER_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_329_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18658_ _23059_/Q _17591_/X _18658_/S vssd1 vssd1 vccd1 vccd1 _18659_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17609_ _17609_/A vssd1 vssd1 vccd1 vccd1 _22697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18589_ _16863_/X _23028_/Q _18597_/S vssd1 vssd1 vccd1 vccd1 _18590_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20620_ _20626_/A _20620_/B _20620_/C vssd1 vssd1 vccd1 vccd1 _20620_/X sky130_fd_sc_hd__or3_1
XFILLER_269_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20551_ _14970_/S _13481_/B _13455_/Y vssd1 vssd1 vccd1 vccd1 _20662_/A sky130_fd_sc_hd__a21o_1
XFILLER_164_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23270_ _23494_/CLK _23270_/D vssd1 vssd1 vccd1 vccd1 _23270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_319_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20482_ _21177_/A _20482_/B vssd1 vssd1 vccd1 vccd1 _20482_/Y sky130_fd_sc_hd__nand2_1
XFILLER_335_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_319_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22221_ _22222_/A _22222_/B vssd1 vssd1 vccd1 vccd1 _22223_/A sky130_fd_sc_hd__nor2_1
XFILLER_336_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_307_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_335_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22152_ _22151_/X _22136_/B _22134_/B vssd1 vssd1 vccd1 vccd1 _22153_/B sky130_fd_sc_hd__a21oi_1
XFILLER_336_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput430 _22555_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[2] sky130_fd_sc_hd__buf_2
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_306_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput441 output441/A vssd1 vssd1 vccd1 vccd1 probe_env[0] sky130_fd_sc_hd__buf_2
XFILLER_105_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21103_ _23849_/Q _21096_/X _21098_/X _20571_/A vssd1 vssd1 vccd1 vccd1 _21104_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_160_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput452 _22888_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[3] sky130_fd_sc_hd__buf_2
XTAP_6818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22083_ _22083_/A _22083_/B vssd1 vssd1 vccd1 vccd1 _22083_/Y sky130_fd_sc_hd__nand2_1
Xoutput463 _23922_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[11] sky130_fd_sc_hd__buf_2
XFILLER_102_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput474 _23932_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[21] sky130_fd_sc_hd__buf_2
XFILLER_321_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput485 _23942_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[31] sky130_fd_sc_hd__buf_2
Xoutput496 _13666_/X vssd1 vssd1 vccd1 vccd1 web0 sky130_fd_sc_hd__buf_2
XFILLER_287_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21034_ _23828_/Q _20993_/X _21033_/Y _21023_/X vssd1 vssd1 vccd1 vccd1 _23828_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_304_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22985_ _23424_/CLK _22985_/D vssd1 vssd1 vccd1 vccd1 _22985_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_103_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21936_ _21936_/A _21936_/B _21936_/C vssd1 vssd1 vccd1 vccd1 _21936_/X sky130_fd_sc_hd__and3_1
XFILLER_320_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21867_ _21867_/A vssd1 vssd1 vccd1 vccd1 _21867_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23606_ _23637_/CLK _23606_/D vssd1 vssd1 vccd1 vccd1 _23606_/Q sky130_fd_sc_hd__dfxtp_1
X_11620_ _23414_/Q _23030_/Q _23382_/Q _23350_/Q _11561_/A _11568_/A vssd1 vssd1 vccd1
+ vccd1 _11620_/X sky130_fd_sc_hd__mux4_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20818_ _20645_/B _20810_/X _20811_/X _23760_/Q vssd1 vssd1 vccd1 vccd1 _20819_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21798_ _21725_/X _21724_/A _21724_/B vssd1 vssd1 vccd1 vccd1 _21798_/X sky130_fd_sc_hd__o21ba_1
XFILLER_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_329_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11551_ _11541_/X _11546_/X _11548_/X _11550_/X _11278_/A vssd1 vssd1 vccd1 vccd1
+ _11552_/C sky130_fd_sc_hd__a221o_1
X_23537_ _23537_/CLK _23537_/D vssd1 vssd1 vccd1 vccd1 _23537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20749_ _20749_/A _20759_/B vssd1 vssd1 vccd1 vccd1 _20752_/B sky130_fd_sc_hd__and2_1
XFILLER_156_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_345_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_345_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14270_ _12605_/A _13240_/Y _14329_/S vssd1 vssd1 vccd1 vccd1 _14270_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11482_ _21848_/A _11481_/X _15671_/A vssd1 vssd1 vccd1 vccd1 _11482_/Y sky130_fd_sc_hd__o21ai_1
X_23468_ _23564_/CLK _23468_/D vssd1 vssd1 vccd1 vccd1 _23468_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_160_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23684_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13221_ _13225_/A _13221_/B vssd1 vssd1 vccd1 vccd1 _13221_/X sky130_fd_sc_hd__or2_1
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22419_ _23491_/CLK _22419_/D vssd1 vssd1 vccd1 vccd1 _22419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_326_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23399_ _23555_/CLK _23399_/D vssd1 vssd1 vccd1 vccd1 _23399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13152_ _11235_/A _13143_/Y _13147_/Y _13149_/Y _13151_/Y vssd1 vssd1 vccd1 vccd1
+ _13152_/X sky130_fd_sc_hd__o32a_1
XFILLER_353_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_341_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12103_ _12091_/A _12102_/X _11630_/A vssd1 vssd1 vccd1 vccd1 _12103_/X sky130_fd_sc_hd__o21a_1
XFILLER_341_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_298_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17960_ _22830_/Q _17956_/X _17959_/X input276/X _17951_/X vssd1 vssd1 vccd1 vccd1
+ _17960_/X sky130_fd_sc_hd__a221o_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _13083_/A vssd1 vssd1 vccd1 vccd1 _13561_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_312_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_300_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_300_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_297_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12034_ _22468_/Q _22628_/Q _22307_/Q _23443_/Q _12029_/X _12009_/X vssd1 vssd1 vccd1
+ vccd1 _12034_/X sky130_fd_sc_hd__mux4_1
X_16911_ _19261_/A vssd1 vssd1 vccd1 vccd1 _16911_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17891_ _17932_/A vssd1 vssd1 vccd1 vccd1 _17891_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_239_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19630_ _19163_/X _23461_/Q _19638_/S vssd1 vssd1 vccd1 vccd1 _19631_/A sky130_fd_sc_hd__mux2_1
X_16842_ _16841_/X _22529_/Q _16845_/S vssd1 vssd1 vccd1 vccd1 _16843_/A sky130_fd_sc_hd__mux2_1
XFILLER_254_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19561_ _19561_/A vssd1 vssd1 vccd1 vccd1 _23430_/D sky130_fd_sc_hd__clkbuf_1
X_16773_ _22509_/Q _16765_/X _16766_/X input24/X vssd1 vssd1 vccd1 vccd1 _16774_/B
+ sky130_fd_sc_hd__o22a_1
X_13985_ _13985_/A _13985_/B vssd1 vssd1 vccd1 vccd1 _13986_/A sky130_fd_sc_hd__and2_2
XFILLER_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18512_ _18507_/X _18511_/Y _18503_/X vssd1 vssd1 vccd1 vccd1 _22999_/D sky130_fd_sc_hd__a21oi_1
X_12936_ _22281_/Q _23097_/Q _23513_/Q _22442_/Q _12819_/S _11166_/A vssd1 vssd1 vccd1
+ vccd1 _12937_/B sky130_fd_sc_hd__mux4_1
X_15724_ _22933_/Q vssd1 vssd1 vccd1 vccd1 _15724_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_46_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19492_ _19175_/X _23400_/Q _19494_/S vssd1 vssd1 vccd1 vccd1 _19493_/A sky130_fd_sc_hd__mux2_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18443_ _19987_/A vssd1 vssd1 vccd1 vccd1 _19950_/A sky130_fd_sc_hd__buf_4
XFILLER_261_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ _22931_/Q _15299_/B _15644_/X _15654_/Y _14431_/A vssd1 vssd1 vccd1 vccd1
+ _15655_/X sky130_fd_sc_hd__a221o_1
XFILLER_206_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12867_ _13029_/A _13028_/A vssd1 vssd1 vccd1 vccd1 _13495_/A sky130_fd_sc_hd__and2_1
XFILLER_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _11818_/A vssd1 vssd1 vccd1 vccd1 _11819_/A sky130_fd_sc_hd__buf_2
X_14606_ _14606_/A vssd1 vssd1 vccd1 vccd1 _14606_/X sky130_fd_sc_hd__clkbuf_4
X_18374_ _14989_/X _18375_/C _22952_/Q vssd1 vssd1 vccd1 vccd1 _18376_/B sky130_fd_sc_hd__a21oi_1
X_15586_ _14632_/A _15540_/X _15581_/X _15585_/X vssd1 vssd1 vccd1 vccd1 _15586_/X
+ sky130_fd_sc_hd__o211a_2
X_12798_ _12784_/A _12796_/X _12797_/X vssd1 vssd1 vccd1 vccd1 _12798_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _17382_/A _17325_/B vssd1 vssd1 vccd1 vccd1 _17326_/C sky130_fd_sc_hd__nor2_1
X_14537_ _19090_/B vssd1 vssd1 vccd1 vccd1 _17471_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11749_ _23216_/Q _23184_/Q _23152_/Q _23120_/Q _11741_/X _12009_/A vssd1 vssd1 vccd1
+ vccd1 _11750_/B sky130_fd_sc_hd__mux4_1
XFILLER_147_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_308_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_348_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17256_ input95/X input60/X _17266_/S vssd1 vssd1 vccd1 vccd1 _17256_/X sky130_fd_sc_hd__mux2_8
XFILLER_175_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14468_ _14595_/B _14468_/B vssd1 vssd1 vccd1 vccd1 _15729_/S sky130_fd_sc_hd__or2_2
XFILLER_335_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16207_ _16288_/A vssd1 vssd1 vccd1 vccd1 _16307_/S sky130_fd_sc_hd__buf_6
X_13419_ _13470_/A vssd1 vssd1 vccd1 vccd1 _15080_/A sky130_fd_sc_hd__buf_8
X_17187_ _17169_/X _17186_/X _17107_/X _17127_/X vssd1 vssd1 vccd1 vccd1 _17187_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_351_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14399_ _14467_/C _14467_/B vssd1 vssd1 vccd1 vccd1 _14473_/A sky130_fd_sc_hd__or2_1
XFILLER_350_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16138_ _23747_/Q _23877_/Q _16138_/S vssd1 vssd1 vccd1 vccd1 _16138_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_343_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_288_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_304_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16069_ _14730_/A _16062_/X _16068_/Y _15150_/A vssd1 vssd1 vccd1 vccd1 _16070_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_335_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_297_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19828_ _19828_/A vssd1 vssd1 vccd1 vccd1 _19837_/S sky130_fd_sc_hd__buf_6
XFILLER_97_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19759_ _19249_/X _23519_/Q _19765_/S vssd1 vssd1 vccd1 vccd1 _19760_/A sky130_fd_sc_hd__mux2_1
XFILLER_284_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22770_ _23070_/CLK _22770_/D vssd1 vssd1 vccd1 vccd1 _22770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21721_ _21849_/A vssd1 vssd1 vccd1 vccd1 _21721_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21652_ _21652_/A _21867_/A vssd1 vssd1 vccd1 vccd1 _21653_/C sky130_fd_sc_hd__nand2_1
XFILLER_33_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20603_ _23722_/Q _20593_/X _20601_/X _20602_/X vssd1 vssd1 vccd1 vccd1 _23722_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21583_ _23822_/Q _23756_/Q vssd1 vssd1 vccd1 vccd1 _21585_/A sky130_fd_sc_hd__or2_1
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_327_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23322_ _23548_/CLK _23322_/D vssd1 vssd1 vccd1 vccd1 _23322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_327_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20534_ _13779_/A _20536_/B _20533_/Y _20549_/A vssd1 vssd1 vccd1 vccd1 _20535_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_192_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_326_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23253_ _23541_/CLK _23253_/D vssd1 vssd1 vccd1 vccd1 _23253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_308_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20465_ _23705_/Q _20468_/B vssd1 vssd1 vccd1 vccd1 _20465_/X sky130_fd_sc_hd__or2_1
XFILLER_119_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22204_ _22205_/A _22205_/B vssd1 vssd1 vccd1 vccd1 _22206_/A sky130_fd_sc_hd__nand2_1
XFILLER_106_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_322_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23184_ _23474_/CLK _23184_/D vssd1 vssd1 vccd1 vccd1 _23184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_334_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20396_ _20396_/A _20396_/B vssd1 vssd1 vccd1 vccd1 _20396_/X sky130_fd_sc_hd__or2_1
XTAP_7327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22135_ _22110_/A _22109_/A _22108_/Y vssd1 vssd1 vccd1 vccd1 _22136_/B sky130_fd_sc_hd__o21ai_1
XTAP_7349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput293 _14100_/X vssd1 vssd1 vccd1 vccd1 addr0[8] sky130_fd_sc_hd__buf_2
X_22066_ _22085_/A _22066_/B vssd1 vssd1 vccd1 vccd1 _22066_/X sky130_fd_sc_hd__xor2_1
XFILLER_121_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_0 _23709_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21017_ _20615_/A _21008_/X _21016_/X _21010_/X vssd1 vssd1 vccd1 vccd1 _23821_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_290_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_331_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13770_ _13807_/A _13770_/B vssd1 vssd1 vccd1 vccd1 _13770_/Y sky130_fd_sc_hd__nor2_1
XFILLER_261_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22968_ _22968_/CLK _22968_/D vssd1 vssd1 vccd1 vccd1 _22968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12721_ _12721_/A vssd1 vssd1 vccd1 vccd1 _12721_/X sky130_fd_sc_hd__buf_2
XFILLER_71_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21919_ _21919_/A _21919_/B vssd1 vssd1 vccd1 vccd1 _21919_/X sky130_fd_sc_hd__xor2_1
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22899_ _22899_/CLK _22899_/D vssd1 vssd1 vccd1 vccd1 _22899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15440_ _15440_/A vssd1 vssd1 vccd1 vccd1 _15440_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12652_ _23413_/Q _23029_/Q _23381_/Q _23349_/Q _12680_/A _12041_/A vssd1 vssd1 vccd1
+ vccd1 _12652_/X sky130_fd_sc_hd__mux4_2
XFILLER_90_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11603_ _11603_/A vssd1 vssd1 vccd1 vccd1 _12463_/A sky130_fd_sc_hd__clkbuf_4
X_15371_ _18808_/A vssd1 vssd1 vccd1 vccd1 _19201_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_212_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12583_ _12590_/A _12582_/X _11679_/A vssd1 vssd1 vccd1 vccd1 _12583_/X sky130_fd_sc_hd__o21a_1
XFILLER_230_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17110_ _17070_/X _17102_/X _17108_/X _17109_/X vssd1 vssd1 vccd1 vccd1 _17110_/X
+ sky130_fd_sc_hd__o211a_4
X_14322_ _14320_/X _14321_/X _14331_/S vssd1 vssd1 vccd1 vccd1 _14323_/A sky130_fd_sc_hd__mux2_1
X_18090_ _18105_/A vssd1 vssd1 vccd1 vccd1 _18090_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11534_ _13127_/A vssd1 vssd1 vccd1 vccd1 _11544_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_318_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_317_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17041_ input73/X input98/X _17084_/S vssd1 vssd1 vccd1 vccd1 _17041_/X sky130_fd_sc_hd__mux2_8
XFILLER_156_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14253_ _16054_/B vssd1 vssd1 vccd1 vccd1 _15582_/B sky130_fd_sc_hd__clkbuf_4
X_11465_ _13291_/A vssd1 vssd1 vccd1 vccd1 _15630_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13204_ _13084_/A _13203_/X _12816_/A vssd1 vssd1 vccd1 vccd1 _13204_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14184_ _23882_/Q vssd1 vssd1 vccd1 vccd1 _14196_/A sky130_fd_sc_hd__buf_6
XFILLER_325_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11396_ _13314_/A _11396_/B vssd1 vssd1 vccd1 vccd1 _13554_/A sky130_fd_sc_hd__nand2_4
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_297_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13135_ _11278_/A _13124_/X _13134_/X _13295_/A vssd1 vssd1 vccd1 vccd1 _20368_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18992_ _19003_/A vssd1 vssd1 vccd1 vccd1 _19001_/S sky130_fd_sc_hd__buf_2
XFILLER_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _22826_/Q _17932_/X _17942_/X _17930_/X vssd1 vssd1 vccd1 vccd1 _22826_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_300_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13066_ _13073_/A _13065_/X _11537_/X vssd1 vssd1 vccd1 vccd1 _13066_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12017_ _12025_/A vssd1 vssd1 vccd1 vccd1 _12734_/A sky130_fd_sc_hd__buf_6
XFILLER_66_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17874_ _22808_/Q _17645_/X _17874_/S vssd1 vssd1 vccd1 vccd1 _17875_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19613_ _23454_/Q _19245_/A _19621_/S vssd1 vssd1 vccd1 vccd1 _19614_/A sky130_fd_sc_hd__mux2_1
XFILLER_266_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_293_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16825_ _19175_/A vssd1 vssd1 vccd1 vccd1 _16825_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19544_ _19544_/A vssd1 vssd1 vccd1 vccd1 _23423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16756_ _16759_/A _16756_/B vssd1 vssd1 vccd1 vccd1 _16757_/A sky130_fd_sc_hd__or2_1
XFILLER_207_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13968_ _13968_/A vssd1 vssd1 vccd1 vccd1 _13968_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_281_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15707_ _22996_/Q _15780_/A _15781_/A input224/X vssd1 vssd1 vccd1 vccd1 _21888_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12919_ _12919_/A _12919_/B vssd1 vssd1 vccd1 vccd1 _12919_/Y sky130_fd_sc_hd__nor2_1
X_19475_ _23393_/Q _18862_/X _19477_/S vssd1 vssd1 vccd1 vccd1 _19476_/A sky130_fd_sc_hd__mux2_1
XFILLER_250_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16687_ _16679_/A _16691_/A _22519_/Q vssd1 vssd1 vccd1 vccd1 _16783_/A sky130_fd_sc_hd__a21oi_4
X_13899_ _21351_/A _14757_/A _13931_/A vssd1 vssd1 vccd1 vccd1 _14082_/A sky130_fd_sc_hd__mux2_8
XFILLER_250_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18426_ _18427_/A _18427_/C _22970_/Q vssd1 vssd1 vccd1 vccd1 _18428_/B sky130_fd_sc_hd__a21oi_1
XFILLER_222_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15638_ _13535_/Y _15196_/X _14761_/A _13536_/Y vssd1 vssd1 vccd1 vccd1 _15638_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_349_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18357_ _22946_/Q _22945_/Q _18357_/C vssd1 vssd1 vccd1 vccd1 _18359_/B sky130_fd_sc_hd__and3_1
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15569_ _18820_/A vssd1 vssd1 vccd1 vccd1 _19213_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_309_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_336_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17308_ _23491_/Q _17016_/X _17017_/X _17268_/X _17307_/Y vssd1 vssd1 vccd1 vccd1
+ _17308_/X sky130_fd_sc_hd__a32o_1
XFILLER_148_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18288_ _22921_/Q _22922_/Q _22923_/Q _18288_/D vssd1 vssd1 vccd1 vccd1 _18298_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_119_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17239_ _22576_/Q _17199_/X _17190_/X _17238_/X vssd1 vssd1 vccd1 vccd1 _22576_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_324_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_305_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_305_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20250_ _20250_/A _20250_/B vssd1 vssd1 vccd1 vccd1 _20250_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20181_ _20236_/A _20179_/X _20180_/Y _20174_/A vssd1 vssd1 vccd1 vccd1 _20181_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_170_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_320_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23940_ _23942_/CLK _23940_/D vssd1 vssd1 vccd1 vccd1 _23940_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23871_ _23871_/CLK _23871_/D vssd1 vssd1 vccd1 vccd1 _23871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22822_ _22822_/CLK _22822_/D vssd1 vssd1 vccd1 vccd1 _22822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_272_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22753_ _23367_/CLK _22753_/D vssd1 vssd1 vccd1 vccd1 _22753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21704_ _21667_/A _21669_/B _21667_/B vssd1 vssd1 vccd1 vccd1 _21705_/B sky130_fd_sc_hd__a21boi_1
XFILLER_240_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22684_ _23563_/CLK _22684_/D vssd1 vssd1 vccd1 vccd1 _22684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21635_ _21636_/A _21641_/A vssd1 vssd1 vccd1 vccd1 _21637_/A sky130_fd_sc_hd__nand2_1
XFILLER_233_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21566_ _21566_/A _21566_/B vssd1 vssd1 vccd1 vccd1 _21567_/B sky130_fd_sc_hd__xnor2_4
X_23305_ _23529_/CLK _23305_/D vssd1 vssd1 vccd1 vccd1 _23305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20517_ _23701_/Q _20517_/B _20517_/C vssd1 vssd1 vccd1 vccd1 _20520_/B sky130_fd_sc_hd__and3_1
XFILLER_153_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_354_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21497_ _22019_/A vssd1 vssd1 vccd1 vccd1 _22083_/A sky130_fd_sc_hd__buf_4
XFILLER_342_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_308_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23236_ _23556_/CLK _23236_/D vssd1 vssd1 vccd1 vccd1 _23236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11250_ _14132_/A _14172_/B vssd1 vssd1 vccd1 vccd1 _11382_/B sky130_fd_sc_hd__nor2_2
XFILLER_342_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_307_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20448_ _23698_/Q _20448_/B vssd1 vssd1 vccd1 vccd1 _20448_/X sky130_fd_sc_hd__or2_1
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_307_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23167_ _23582_/CLK _23167_/D vssd1 vssd1 vccd1 vccd1 _23167_/Q sky130_fd_sc_hd__dfxtp_1
X_11181_ _13091_/A vssd1 vssd1 vccd1 vccd1 _13158_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20379_ _20379_/A _21177_/A vssd1 vssd1 vccd1 vccd1 _20379_/Y sky130_fd_sc_hd__nand2_1
XFILLER_323_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22118_ _22118_/A _22118_/B vssd1 vssd1 vccd1 vccd1 _22118_/Y sky130_fd_sc_hd__xnor2_2
XTAP_7179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_322_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23098_ _23546_/CLK _23098_/D vssd1 vssd1 vccd1 vccd1 _23098_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22049_ _17246_/A _22044_/X _22047_/Y _22048_/X vssd1 vssd1 vccd1 vccd1 _22051_/B
+ sky130_fd_sc_hd__o22a_1
X_14940_ _14940_/A _14940_/B vssd1 vssd1 vccd1 vccd1 _14940_/Y sky130_fd_sc_hd__nand2_1
XTAP_6489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14871_ _23720_/Q _23850_/Q _15354_/S vssd1 vssd1 vccd1 vccd1 _14871_/X sky130_fd_sc_hd__mux2_2
XFILLER_36_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16610_ _22454_/Q _16200_/X _16618_/S vssd1 vssd1 vccd1 vccd1 _16611_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13822_ _13790_/X _13768_/Y _13820_/Y _13821_/Y vssd1 vssd1 vccd1 vccd1 _14052_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_75_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17590_ _17590_/A vssd1 vssd1 vccd1 vccd1 _22691_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_107 _13521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13753_ _13711_/B _13874_/A _13847_/A _13721_/B vssd1 vssd1 vccd1 vccd1 _13754_/B
+ sky130_fd_sc_hd__o22a_4
X_16541_ _16541_/A vssd1 vssd1 vccd1 vccd1 _22423_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_118 _20217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_129 _13695_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12704_ _12891_/A _12704_/B vssd1 vssd1 vccd1 vccd1 _12704_/Y sky130_fd_sc_hd__nand2_1
X_19260_ _19260_/A vssd1 vssd1 vccd1 vccd1 _23298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13684_ _15830_/A vssd1 vssd1 vccd1 vccd1 _14072_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16472_ _15044_/X _22394_/Q _16480_/S vssd1 vssd1 vccd1 vccd1 _16473_/A sky130_fd_sc_hd__mux2_1
XFILLER_349_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18211_ hold3/X _18202_/X _18210_/X _18206_/X vssd1 vssd1 vccd1 vccd1 _22896_/D sky130_fd_sc_hd__o211a_1
XPHY_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15423_ _15422_/X _22273_/Q _15524_/S vssd1 vssd1 vccd1 vccd1 _15424_/A sky130_fd_sc_hd__mux2_1
X_12635_ _23927_/Q _20296_/A _12739_/A vssd1 vssd1 vccd1 vccd1 _12636_/A sky130_fd_sc_hd__mux2_1
X_19191_ _19191_/A vssd1 vssd1 vccd1 vccd1 _19191_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_358_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18142_ _18142_/A _18167_/A vssd1 vssd1 vccd1 vccd1 _18164_/A sky130_fd_sc_hd__nor2_1
XPHY_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15354_ _23728_/Q _23858_/Q _15354_/S vssd1 vssd1 vccd1 vccd1 _15354_/X sky130_fd_sc_hd__mux2_1
X_12566_ _22265_/Q _23081_/Q _23497_/Q _22426_/Q _12245_/S _12292_/X vssd1 vssd1 vccd1
+ vccd1 _12567_/B sky130_fd_sc_hd__mux4_1
XFILLER_357_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_306_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11517_ _11517_/A vssd1 vssd1 vccd1 vccd1 _11517_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_145_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14305_ _13019_/Y _11939_/B _14326_/S vssd1 vssd1 vccd1 vccd1 _14305_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_345_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18073_ _22862_/Q _18066_/X _18072_/X _18060_/X vssd1 vssd1 vccd1 vccd1 _22862_/D
+ sky130_fd_sc_hd__o211a_1
X_15285_ _15285_/A vssd1 vssd1 vccd1 vccd1 _22270_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_333_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12497_ _14292_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _14687_/A sky130_fd_sc_hd__xnor2_4
XFILLER_333_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14236_ input149/X _13651_/B _15033_/S input114/X _14235_/X vssd1 vssd1 vccd1 vccd1
+ _14236_/X sky130_fd_sc_hd__a221o_4
X_17024_ _17262_/A _17283_/A vssd1 vssd1 vccd1 vccd1 _17024_/X sky130_fd_sc_hd__or2_2
XFILLER_172_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11448_ _13041_/A _11448_/B vssd1 vssd1 vccd1 vccd1 _11448_/X sky130_fd_sc_hd__or2_1
XFILLER_171_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14167_ _16962_/A _20140_/B vssd1 vssd1 vccd1 vccd1 _14167_/X sky130_fd_sc_hd__or2_4
X_11379_ _11379_/A vssd1 vssd1 vccd1 vccd1 _11483_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_152_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13118_ _23487_/Q _23583_/Q _22547_/Q _22351_/Q _13114_/X _13115_/X vssd1 vssd1 vccd1
+ vccd1 _13119_/B sky130_fd_sc_hd__mux4_2
XFILLER_298_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_286_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18975_ _16854_/X _23185_/Q _18979_/S vssd1 vssd1 vccd1 vccd1 _18976_/A sky130_fd_sc_hd__mux2_1
X_14098_ _22596_/Q _14081_/A _14097_/Y _14012_/X vssd1 vssd1 vccd1 vccd1 _14098_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17926_ _17926_/A _17987_/S vssd1 vssd1 vccd1 vccd1 _17926_/X sky130_fd_sc_hd__or2b_1
X_13049_ _13095_/A _13048_/X _11134_/A vssd1 vssd1 vccd1 vccd1 _13049_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_39_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17857_ _22800_/Q _17620_/X _17859_/S vssd1 vssd1 vccd1 vccd1 _17858_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_294_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16808_ _16808_/A _16808_/B _16808_/C _16808_/D vssd1 vssd1 vccd1 vccd1 _16809_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17788_ _17788_/A vssd1 vssd1 vccd1 vccd1 _22769_/D sky130_fd_sc_hd__clkbuf_1
X_19527_ _19226_/X _23416_/Q _19527_/S vssd1 vssd1 vccd1 vccd1 _19528_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16739_ _16739_/A vssd1 vssd1 vccd1 vccd1 _22499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19458_ _23385_/Q _18836_/X _19466_/S vssd1 vssd1 vccd1 vccd1 _19459_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18409_ _22963_/Q _22964_/Q _18409_/C vssd1 vssd1 vccd1 vccd1 _18412_/B sky130_fd_sc_hd__and3_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19389_ _19389_/A vssd1 vssd1 vccd1 vccd1 _23354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_349_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21420_ _15929_/X _15631_/A _21336_/X _14535_/X vssd1 vssd1 vccd1 vccd1 _21452_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_349_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21351_ _21351_/A _21351_/B vssd1 vssd1 vccd1 vccd1 _21352_/B sky130_fd_sc_hd__nor2_1
XFILLER_337_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_336_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_351_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20302_ _20320_/A vssd1 vssd1 vccd1 vccd1 _20302_/X sky130_fd_sc_hd__clkbuf_2
X_21282_ _21079_/B _21199_/B _21280_/Y _21281_/X vssd1 vssd1 vccd1 vccd1 _23909_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_352_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23021_ _23534_/CLK _23021_/D vssd1 vssd1 vccd1 vccd1 _23021_/Q sky130_fd_sc_hd__dfxtp_1
X_20233_ _23660_/Q _20165_/X _20232_/Y _20203_/X vssd1 vssd1 vccd1 vccd1 _23660_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_305_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20164_ _20146_/X _20543_/A _20163_/X _18547_/X vssd1 vssd1 vccd1 vccd1 _23653_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20095_ _23639_/Q _20098_/C _23637_/Q _20095_/D vssd1 vssd1 vccd1 vccd1 _20110_/C
+ sky130_fd_sc_hd__and4_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23923_ _23934_/CLK _23923_/D vssd1 vssd1 vccd1 vccd1 _23923_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23854_ _23856_/CLK _23854_/D vssd1 vssd1 vccd1 vccd1 _23854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_309_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22805_ _23073_/CLK _22805_/D vssd1 vssd1 vccd1 vccd1 _22805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23785_ _23862_/CLK _23785_/D vssd1 vssd1 vccd1 vccd1 _23785_/Q sky130_fd_sc_hd__dfxtp_4
X_20997_ _21023_/A vssd1 vssd1 vccd1 vccd1 _20997_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22736_ _23068_/CLK _22736_/D vssd1 vssd1 vccd1 vccd1 _22736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22667_ _23580_/CLK _22667_/D vssd1 vssd1 vccd1 vccd1 _22667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12420_ _23207_/Q _23175_/Q _23143_/Q _23111_/Q _12244_/A _12292_/A vssd1 vssd1 vccd1
+ vccd1 _12421_/B sky130_fd_sc_hd__mux4_1
XFILLER_346_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21618_ _21616_/Y _21617_/X _21598_/X vssd1 vssd1 vccd1 vccd1 _21618_/Y sky130_fd_sc_hd__a21oi_2
X_22598_ _22974_/CLK _22598_/D vssd1 vssd1 vccd1 vccd1 _22598_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_224_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_355_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_327_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12351_ _22780_/Q _22748_/Q _22649_/Q _22716_/Q _11112_/A _11702_/A vssd1 vssd1 vccd1
+ vccd1 _12351_/X sky130_fd_sc_hd__mux4_2
XFILLER_337_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_67_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23446_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21549_ _21549_/A vssd1 vssd1 vccd1 vccd1 _21550_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_126_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_343_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11302_ _12475_/A vssd1 vssd1 vccd1 vccd1 _12324_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15070_ _23755_/Q _15595_/A _15596_/A _15069_/X _14917_/A vssd1 vssd1 vccd1 vccd1
+ _15070_/X sky130_fd_sc_hd__a221o_1
XFILLER_138_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12282_ _12414_/A _12282_/B _12282_/C vssd1 vssd1 vccd1 vccd1 _20217_/A sky130_fd_sc_hd__nor3_4
XFILLER_316_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14021_ _14072_/B _14036_/B _14021_/C vssd1 vssd1 vccd1 vccd1 _14021_/X sky130_fd_sc_hd__and3_1
XFILLER_342_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11233_ _11233_/A vssd1 vssd1 vccd1 vccd1 _12816_/A sky130_fd_sc_hd__buf_2
X_23219_ _23507_/CLK _23219_/D vssd1 vssd1 vccd1 vccd1 _23219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_330_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11164_ _11953_/A vssd1 vssd1 vccd1 vccd1 _12685_/A sky130_fd_sc_hd__buf_6
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_310_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_296_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_295_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18760_ _18760_/A vssd1 vssd1 vccd1 vccd1 _23104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15972_ _22087_/B vssd1 vssd1 vccd1 vccd1 _22116_/B sky130_fd_sc_hd__clkbuf_4
X_11095_ _13775_/B _11095_/B _11095_/C _15081_/B vssd1 vssd1 vccd1 vccd1 _13459_/A
+ sky130_fd_sc_hd__or4b_2
XTAP_6286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17711_ _22735_/Q _17617_/X _17715_/S vssd1 vssd1 vccd1 vccd1 _17712_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14923_ _14923_/A vssd1 vssd1 vccd1 vccd1 _14923_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18691_ _23074_/Q _17639_/X _18691_/S vssd1 vssd1 vccd1 vccd1 _18692_/A sky130_fd_sc_hd__mux2_1
XFILLER_282_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_291_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17642_ _18868_/A vssd1 vssd1 vccd1 vccd1 _17642_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14854_ _14853_/X _14375_/Y _14854_/S vssd1 vssd1 vccd1 vccd1 _14855_/B sky130_fd_sc_hd__mux2_1
XFILLER_75_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_291_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13805_ _13821_/A _14015_/C vssd1 vssd1 vccd1 vccd1 _13851_/A sky130_fd_sc_hd__nor2_1
XFILLER_251_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17573_ _22686_/Q _17572_/X _17576_/S vssd1 vssd1 vccd1 vccd1 _17574_/A sky130_fd_sc_hd__mux2_1
X_11997_ _12909_/A _11997_/B vssd1 vssd1 vccd1 vccd1 _11997_/X sky130_fd_sc_hd__or2_1
X_14785_ _14354_/A _14341_/X _14840_/S vssd1 vssd1 vccd1 vccd1 _14785_/X sky130_fd_sc_hd__mux2_1
X_19312_ _19312_/A vssd1 vssd1 vccd1 vccd1 _23320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16524_ _16124_/X _22418_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _16525_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13736_ _13890_/B _13736_/B vssd1 vssd1 vccd1 vccd1 _13737_/A sky130_fd_sc_hd__nor2_2
XFILLER_177_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19243_ _19242_/X _23293_/Q _19243_/S vssd1 vssd1 vccd1 vccd1 _19244_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16455_ _16197_/X _22388_/Q _16455_/S vssd1 vssd1 vccd1 vccd1 _16456_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13667_ _13993_/A _14069_/B vssd1 vssd1 vccd1 vccd1 _14001_/A sky130_fd_sc_hd__nor2_2
XFILLER_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15406_ _22926_/Q _14588_/A _15395_/X _15405_/Y _15558_/A vssd1 vssd1 vccd1 vccd1
+ _15406_/X sky130_fd_sc_hd__a221o_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12618_ _12852_/A _12617_/X _11681_/X vssd1 vssd1 vccd1 vccd1 _12618_/Y sky130_fd_sc_hd__o21ai_1
X_19174_ _19174_/A vssd1 vssd1 vccd1 vccd1 _23271_/D sky130_fd_sc_hd__clkbuf_1
X_16386_ _16442_/A vssd1 vssd1 vccd1 vccd1 _16455_/S sky130_fd_sc_hd__buf_6
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13598_ _13532_/D _13629_/B _15678_/A vssd1 vssd1 vccd1 vccd1 _13599_/B sky130_fd_sc_hd__a21oi_2
XFILLER_129_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18125_ _18116_/Y _18123_/X _18124_/X _18121_/X vssd1 vssd1 vccd1 vccd1 _22879_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_318_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15337_ _15089_/S _14951_/Y _14860_/X vssd1 vssd1 vccd1 vccd1 _15338_/B sky130_fd_sc_hd__a21o_1
X_12549_ _13903_/A _13364_/A _14294_/A vssd1 vssd1 vccd1 vccd1 _12549_/X sky130_fd_sc_hd__or3_1
XFILLER_346_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18056_ hold4/A _18051_/X _18055_/X _18045_/X vssd1 vssd1 vccd1 vccd1 _22856_/D sky130_fd_sc_hd__o211a_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15268_ _14592_/X _15260_/X _15267_/X _14498_/X vssd1 vssd1 vccd1 vccd1 _15268_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_334_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17007_ _21351_/A _17174_/B vssd1 vssd1 vccd1 vccd1 _17007_/Y sky130_fd_sc_hd__nand2_1
X_14219_ _14219_/A vssd1 vssd1 vccd1 vccd1 _14219_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15199_ _13935_/A _14942_/X _15195_/X _14384_/X _15198_/X vssd1 vssd1 vccd1 vccd1
+ _15199_/X sky130_fd_sc_hd__o221a_1
XFILLER_113_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_302_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18958_ _18958_/A vssd1 vssd1 vccd1 vccd1 _23177_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_286_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17909_ _22815_/Q _17908_/X _17903_/X input256/X _17899_/X vssd1 vssd1 vccd1 vccd1
+ _17909_/X sky130_fd_sc_hd__a221o_1
X_18889_ _18889_/A vssd1 vssd1 vccd1 vccd1 _23146_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20920_ _20948_/A vssd1 vssd1 vccd1 vccd1 _20920_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20851_ _20705_/B _20846_/X _20847_/X _23769_/Q vssd1 vssd1 vccd1 vccd1 _20852_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23570_ _23570_/CLK _23570_/D vssd1 vssd1 vccd1 vccd1 _23570_/Q sky130_fd_sc_hd__dfxtp_1
X_20782_ _20781_/Y _20536_/B _20577_/B _20888_/C vssd1 vssd1 vccd1 vccd1 _20782_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_168_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_460 _18012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_471 _11483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22521_ _23896_/CLK _22521_/D vssd1 vssd1 vccd1 vccd1 _22521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_288_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_482 _13981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_493 _14757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22452_ _23491_/CLK _22452_/D vssd1 vssd1 vccd1 vccd1 _22452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_337_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_309_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21403_ _21403_/A _21403_/B vssd1 vssd1 vccd1 vccd1 _21404_/B sky130_fd_sc_hd__or2_1
X_22383_ _23583_/CLK _22383_/D vssd1 vssd1 vccd1 vccd1 _22383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21334_ _20500_/A _20500_/B _21333_/X vssd1 vssd1 vccd1 vccd1 _21344_/A sky130_fd_sc_hd__a21o_1
XFILLER_336_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_307_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21265_ _15674_/X _15865_/Y _21243_/A _20058_/X vssd1 vssd1 vccd1 vccd1 _21265_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_278_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23004_ _23005_/CLK _23004_/D vssd1 vssd1 vccd1 vccd1 _23004_/Q sky130_fd_sc_hd__dfxtp_4
X_20216_ _20216_/A vssd1 vssd1 vccd1 vccd1 _20279_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_235_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_320_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21196_ _21283_/B vssd1 vssd1 vccd1 vccd1 _21196_/X sky130_fd_sc_hd__buf_2
XFILLER_104_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_293_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20147_ _22712_/Q vssd1 vssd1 vccd1 vccd1 _20147_/X sky130_fd_sc_hd__buf_4
XFILLER_77_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_185_wb_clk_i _23931_/CLK vssd1 vssd1 vccd1 vccd1 _23916_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_293_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_253_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20078_ _23634_/Q _23633_/Q vssd1 vssd1 vccd1 vccd1 _20085_/D sky130_fd_sc_hd__and2_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_114_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23009_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_264_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23906_ _23907_/CLK _23906_/D vssd1 vssd1 vccd1 vccd1 _23906_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ _11920_/A vssd1 vssd1 vccd1 vccd1 _11920_/X sky130_fd_sc_hd__buf_6
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11851_ _11834_/A _11850_/X _11780_/X vssd1 vssd1 vccd1 vccd1 _11851_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23837_ _23876_/CLK _23837_/D vssd1 vssd1 vccd1 vccd1 _23837_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _15676_/A vssd1 vssd1 vccd1 vccd1 _14570_/X sky130_fd_sc_hd__buf_2
XFILLER_199_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11782_ _11890_/A _11776_/Y _11778_/Y _11781_/Y vssd1 vssd1 vccd1 vccd1 _11782_/X
+ sky130_fd_sc_hd__a31o_1
X_23768_ _23768_/CLK _23768_/D vssd1 vssd1 vccd1 vccd1 _23768_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_341_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13521_ _13521_/A _13521_/B vssd1 vssd1 vccd1 vccd1 _13528_/A sky130_fd_sc_hd__nor2_1
XFILLER_347_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22719_ _23369_/CLK _22719_/D vssd1 vssd1 vccd1 vccd1 _22719_/Q sky130_fd_sc_hd__dfxtp_1
X_23699_ _23706_/CLK _23699_/D vssd1 vssd1 vccd1 vccd1 _23699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_348_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16240_ _16307_/S vssd1 vssd1 vccd1 vccd1 _16253_/S sky130_fd_sc_hd__buf_4
X_13452_ _20533_/C vssd1 vssd1 vccd1 vccd1 _21285_/A sky130_fd_sc_hd__buf_2
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_356_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12403_ _12406_/A _12402_/X _11347_/A vssd1 vssd1 vccd1 vccd1 _12403_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16171_ _23748_/Q _23878_/Q _16171_/S vssd1 vssd1 vccd1 vccd1 _16171_/X sky130_fd_sc_hd__mux2_1
X_13383_ _13392_/B _13383_/B vssd1 vssd1 vccd1 vccd1 _13383_/X sky130_fd_sc_hd__or2_1
XFILLER_127_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_328_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12334_ _12334_/A _12334_/B vssd1 vssd1 vccd1 vccd1 _12334_/X sky130_fd_sc_hd__or2_1
X_15122_ _15122_/A _15122_/B vssd1 vssd1 vccd1 vccd1 _15122_/X sky130_fd_sc_hd__and2_1
XFILLER_316_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_316_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19930_ _19934_/B _19934_/C _18423_/X vssd1 vssd1 vccd1 vccd1 _19930_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_315_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15053_ _22493_/Q _13692_/A _14247_/X _15052_/X _14072_/A vssd1 vssd1 vccd1 vccd1
+ _15053_/X sky130_fd_sc_hd__o221a_1
XFILLER_181_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12265_ _23403_/Q _23019_/Q _23371_/Q _23339_/Q _11920_/X _11652_/A vssd1 vssd1 vccd1
+ vccd1 _12265_/X sky130_fd_sc_hd__mux4_2
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14004_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14004_/X sky130_fd_sc_hd__buf_2
XFILLER_296_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11216_ _11216_/A vssd1 vssd1 vccd1 vccd1 _11217_/A sky130_fd_sc_hd__buf_4
X_19861_ _16230_/X _23564_/Q _19865_/S vssd1 vssd1 vccd1 vccd1 _19862_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12196_ _12196_/A vssd1 vssd1 vccd1 vccd1 _12196_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_150_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18812_ _23121_/Q _18811_/X _18818_/S vssd1 vssd1 vccd1 vccd1 _18813_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11147_ _11699_/A vssd1 vssd1 vccd1 vccd1 _11148_/A sky130_fd_sc_hd__buf_6
XFILLER_123_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19792_ _19792_/A vssd1 vssd1 vccd1 vccd1 _23533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_311_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18743_ _18754_/A vssd1 vssd1 vccd1 vccd1 _18752_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_237_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15955_ _23742_/Q _23872_/Q _16103_/S vssd1 vssd1 vccd1 vccd1 _15955_/X sky130_fd_sc_hd__mux2_1
X_11078_ _13440_/C _13440_/B _13440_/A vssd1 vssd1 vccd1 vccd1 _14187_/A sky130_fd_sc_hd__and3b_2
XTAP_5371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput160 dout1[58] vssd1 vssd1 vccd1 vccd1 input160/X sky130_fd_sc_hd__buf_2
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput171 irq[0] vssd1 vssd1 vccd1 vccd1 _20517_/C sky130_fd_sc_hd__clkbuf_4
XTAP_5393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput182 irq[5] vssd1 vssd1 vccd1 vccd1 _20516_/C sky130_fd_sc_hd__clkbuf_4
X_14906_ _14906_/A vssd1 vssd1 vccd1 vccd1 _14907_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput193 localMemory_wb_adr_i[12] vssd1 vssd1 vccd1 vccd1 input193/X sky130_fd_sc_hd__clkbuf_1
X_18674_ _23066_/Q _17614_/X _18680_/S vssd1 vssd1 vccd1 vccd1 _18675_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15886_ _22937_/Q _15299_/B _15875_/X _15885_/Y _14431_/A vssd1 vssd1 vccd1 vccd1
+ _15886_/X sky130_fd_sc_hd__a221o_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17625_ _17625_/A vssd1 vssd1 vccd1 vccd1 _22702_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14837_ _15769_/A vssd1 vssd1 vccd1 vccd1 _14837_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17556_ _18782_/A vssd1 vssd1 vccd1 vccd1 _17556_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14768_ _15490_/S _14766_/X _14767_/X vssd1 vssd1 vccd1 vccd1 _14768_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_189_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16507_ _15823_/X _22410_/Q _16513_/S vssd1 vssd1 vccd1 vccd1 _16508_/A sky130_fd_sc_hd__mux2_1
X_13719_ _14015_/A _13728_/B _13810_/B vssd1 vssd1 vccd1 vccd1 _13720_/A sky130_fd_sc_hd__and3_4
XFILLER_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17487_ _17487_/A vssd1 vssd1 vccd1 vccd1 _22651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14699_ _14804_/A _14567_/Y _14695_/Y _14698_/X vssd1 vssd1 vccd1 vccd1 _14699_/X
+ sky130_fd_sc_hd__a211o_1
X_19226_ _19226_/A vssd1 vssd1 vccd1 vccd1 _19226_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_258_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16438_ _15898_/X _22380_/Q _16440_/S vssd1 vssd1 vccd1 vccd1 _16439_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_319_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19157_ _23266_/Q _18865_/X _19157_/S vssd1 vssd1 vccd1 vccd1 _19158_/A sky130_fd_sc_hd__mux2_1
X_16369_ _15975_/X _22350_/Q _16377_/S vssd1 vssd1 vccd1 vccd1 _16370_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_307_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18108_ _22874_/Q _18096_/X _18107_/X _18105_/X vssd1 vssd1 vccd1 vccd1 _22874_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_318_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19088_ _16914_/X _23236_/Q _19088_/S vssd1 vssd1 vccd1 vccd1 _19089_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_333_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18039_ _22850_/Q _18036_/X _18037_/X _22983_/Q _18038_/X vssd1 vssd1 vccd1 vccd1
+ _18039_/X sky130_fd_sc_hd__a221o_1
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_334_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21050_ _20708_/A _21047_/X _21048_/X _21049_/X vssd1 vssd1 vccd1 vccd1 _23834_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_302_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20001_ _23613_/Q _19998_/B _20000_/Y vssd1 vssd1 vccd1 vccd1 _23613_/D sky130_fd_sc_hd__o21a_1
XFILLER_286_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_302_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_290_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_286_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21952_ _21919_/A _21918_/B _21918_/A vssd1 vssd1 vccd1 vccd1 _21953_/B sky130_fd_sc_hd__a21bo_1
XFILLER_228_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20903_ _23783_/Q _20893_/X _20902_/X _20788_/X vssd1 vssd1 vccd1 vccd1 _23783_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_54_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21883_ _23831_/Q _23765_/Q vssd1 vssd1 vccd1 vccd1 _21883_/Y sky130_fd_sc_hd__nand2_1
XFILLER_270_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23622_ _23624_/CLK _23622_/D vssd1 vssd1 vccd1 vccd1 _23622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20834_ _20843_/A _20834_/B vssd1 vssd1 vccd1 vccd1 _20835_/A sky130_fd_sc_hd__and2_1
XFILLER_70_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23553_ _23553_/CLK _23553_/D vssd1 vssd1 vccd1 vccd1 _23553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20765_ _20765_/A _21301_/C vssd1 vssd1 vccd1 vccd1 _20888_/B sky130_fd_sc_hd__and2_1
XINSDIODE2_290 _18852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22504_ _23684_/CLK _22504_/D vssd1 vssd1 vccd1 vccd1 _22504_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_196_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23484_ _23546_/CLK _23484_/D vssd1 vssd1 vccd1 vccd1 _23484_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_210_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20696_ _23736_/Q _20667_/X _20695_/X _20673_/X vssd1 vssd1 vccd1 vccd1 _23736_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_338_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22435_ _23538_/CLK _22435_/D vssd1 vssd1 vccd1 vccd1 _22435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_313_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_318_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_353_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22366_ _23566_/CLK _22366_/D vssd1 vssd1 vccd1 vccd1 _22366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_272_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21317_ _21317_/A _21348_/B vssd1 vssd1 vccd1 vccd1 _21318_/B sky130_fd_sc_hd__or2_1
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22297_ _22618_/CLK _22297_/D vssd1 vssd1 vccd1 vccd1 _22297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_352_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12050_ _12700_/A _12040_/Y _12045_/Y _12047_/Y _12049_/Y vssd1 vssd1 vccd1 vccd1
+ _12050_/X sky130_fd_sc_hd__o32a_1
XFILLER_117_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21248_ _21248_/A vssd1 vssd1 vccd1 vccd1 _23895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_352_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_305_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_320_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21179_ _23874_/Q _21168_/A _21177_/Y _21178_/X _21175_/X vssd1 vssd1 vccd1 vccd1
+ _23874_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_291_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_292_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_350_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15740_ _15698_/A _15739_/X _15673_/A vssd1 vssd1 vccd1 vccd1 _15740_/X sky130_fd_sc_hd__a21o_1
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _22281_/Q _23097_/Q _23513_/Q _22442_/Q _12716_/X _12717_/X vssd1 vssd1 vccd1
+ vccd1 _12953_/B sky130_fd_sc_hd__mux4_1
XFILLER_280_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11903_ _11890_/A _11902_/X _11713_/X vssd1 vssd1 vccd1 vccd1 _11903_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _15671_/A vssd1 vssd1 vccd1 vccd1 _15671_/X sky130_fd_sc_hd__clkbuf_8
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _23418_/Q _23034_/Q _23386_/Q _23354_/Q _12922_/S _12746_/X vssd1 vssd1 vccd1
+ vccd1 _12883_/X sky130_fd_sc_hd__mux4_2
XFILLER_34_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17410_ _22618_/Q _16220_/X _17410_/S vssd1 vssd1 vccd1 vccd1 _17411_/A sky130_fd_sc_hd__mux2_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _15338_/A vssd1 vssd1 vccd1 vccd1 _14632_/A sky130_fd_sc_hd__buf_2
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _15351_/A _18392_/C _18389_/Y vssd1 vssd1 vccd1 vccd1 _22957_/D sky130_fd_sc_hd__o21a_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _11834_/A _11834_/B vssd1 vssd1 vccd1 vccd1 _11834_/Y sky130_fd_sc_hd__nor2_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _22592_/Q input209/X _17347_/S vssd1 vssd1 vccd1 vccd1 _17342_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14553_ _14553_/A _16935_/B _14553_/C vssd1 vssd1 vccd1 vccd1 _16953_/B sky130_fd_sc_hd__or3_2
X_11765_ _13521_/A _11944_/A vssd1 vssd1 vccd1 vccd1 _13337_/A sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_82_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23515_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13504_ _14791_/A _14294_/A vssd1 vssd1 vccd1 vccd1 _14794_/A sky130_fd_sc_hd__or2_4
X_17272_ _22114_/A _17271_/X _17292_/S vssd1 vssd1 vccd1 vccd1 _17272_/X sky130_fd_sc_hd__mux2_1
XFILLER_348_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14484_ _14918_/A vssd1 vssd1 vccd1 vccd1 _15067_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_11_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23534_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11696_ _12350_/A vssd1 vssd1 vccd1 vccd1 _11696_/X sky130_fd_sc_hd__buf_4
X_19011_ _19011_/A vssd1 vssd1 vccd1 vccd1 _23201_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16223_ _18788_/A vssd1 vssd1 vccd1 vccd1 _16223_/X sky130_fd_sc_hd__clkbuf_2
X_13435_ _21077_/D vssd1 vssd1 vccd1 vccd1 _13454_/A sky130_fd_sc_hd__buf_6
XFILLER_127_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16154_ _16154_/A _16154_/B vssd1 vssd1 vccd1 vccd1 _16154_/Y sky130_fd_sc_hd__nor2_1
X_13366_ _13903_/A _13366_/B vssd1 vssd1 vccd1 vccd1 _13367_/D sky130_fd_sc_hd__xnor2_1
XFILLER_343_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_315_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15105_ _15104_/X _22267_/Q _15284_/S vssd1 vssd1 vccd1 vccd1 _15106_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12317_ _23210_/Q _23178_/Q _23146_/Q _23114_/Q _12314_/X _11815_/X vssd1 vssd1 vccd1
+ vccd1 _12318_/B sky130_fd_sc_hd__mux4_1
XFILLER_138_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16085_ _16085_/A vssd1 vssd1 vccd1 vccd1 _16085_/X sky130_fd_sc_hd__buf_2
X_13297_ _11398_/A _20381_/A _13296_/X vssd1 vssd1 vccd1 vccd1 _13319_/B sky130_fd_sc_hd__o21ai_2
XFILLER_330_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19913_ _16306_/X _23588_/Q _19913_/S vssd1 vssd1 vccd1 vccd1 _19914_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12248_ _11138_/A _12247_/X _11780_/A vssd1 vssd1 vccd1 vccd1 _12248_/Y sky130_fd_sc_hd__o21ai_1
X_15036_ _14882_/A _15005_/X _15025_/Y _14822_/X _15035_/X vssd1 vssd1 vccd1 vccd1
+ _15036_/X sky130_fd_sc_hd__a32o_2
XFILLER_330_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19844_ _19900_/A vssd1 vssd1 vccd1 vccd1 _19913_/S sky130_fd_sc_hd__buf_6
XFILLER_69_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12179_ _12424_/S vssd1 vssd1 vccd1 vccd1 _12349_/S sky130_fd_sc_hd__buf_2
XFILLER_312_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_311_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19775_ _19775_/A vssd1 vssd1 vccd1 vccd1 _23525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16987_ _17230_/A vssd1 vssd1 vccd1 vccd1 _16987_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18726_ _16854_/X _23089_/Q _18730_/S vssd1 vssd1 vccd1 vccd1 _18727_/A sky130_fd_sc_hd__mux2_1
X_15938_ _15938_/A vssd1 vssd1 vccd1 vccd1 _22285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_260_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18657_ _18657_/A vssd1 vssd1 vccd1 vccd1 _23058_/D sky130_fd_sc_hd__clkbuf_1
X_15869_ _14835_/A _13592_/A _15868_/X vssd1 vssd1 vccd1 vccd1 _15871_/A sky130_fd_sc_hd__a21oi_2
XFILLER_58_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17608_ _22697_/Q _17607_/X _17608_/S vssd1 vssd1 vccd1 vccd1 _17609_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18588_ _18610_/A vssd1 vssd1 vccd1 vccd1 _18597_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_212_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17539_ _17539_/A vssd1 vssd1 vccd1 vccd1 _22675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_338_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20550_ _20724_/A vssd1 vssd1 vccd1 vccd1 _20642_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_177_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19209_ _19209_/A vssd1 vssd1 vccd1 vccd1 _23282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_326_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_295_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20481_ _23711_/Q _20416_/B _20480_/Y _20472_/X vssd1 vssd1 vccd1 vccd1 _23711_/D
+ sky130_fd_sc_hd__o211a_1
X_22220_ _22219_/X _22195_/C _22195_/B vssd1 vssd1 vccd1 vccd1 _22222_/B sky130_fd_sc_hd__a21oi_1
XFILLER_306_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22151_ _22151_/A _23774_/Q vssd1 vssd1 vccd1 vccd1 _22151_/X sky130_fd_sc_hd__or2_1
XFILLER_350_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput420 _22573_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[20] sky130_fd_sc_hd__buf_2
XFILLER_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput431 _22583_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[30] sky130_fd_sc_hd__buf_2
XFILLER_350_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21102_ _21108_/A _21102_/B vssd1 vssd1 vccd1 vccd1 _23848_/D sky130_fd_sc_hd__nor2_1
XFILLER_133_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput442 output442/A vssd1 vssd1 vccd1 vccd1 probe_env[1] sky130_fd_sc_hd__buf_2
XTAP_6808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22082_ _22082_/A _22082_/B vssd1 vssd1 vccd1 vccd1 _22083_/B sky130_fd_sc_hd__xnor2_1
Xoutput453 _22889_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[4] sky130_fd_sc_hd__buf_2
XTAP_6819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput464 _23923_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[12] sky130_fd_sc_hd__buf_2
XFILLER_259_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput475 _23933_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[22] sky130_fd_sc_hd__buf_2
XFILLER_120_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput486 _23914_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[3] sky130_fd_sc_hd__buf_2
X_21033_ _21033_/A _21043_/B vssd1 vssd1 vccd1 vccd1 _21033_/Y sky130_fd_sc_hd__nand2_1
Xoutput497 _14073_/X vssd1 vssd1 vccd1 vccd1 wmask0[0] sky130_fd_sc_hd__buf_2
XFILLER_287_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22984_ _23424_/CLK _22984_/D vssd1 vssd1 vccd1 vccd1 _22984_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21935_ _22039_/A vssd1 vssd1 vccd1 vccd1 _21935_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21866_ _15671_/A _21865_/X _21849_/X vssd1 vssd1 vccd1 vccd1 _21936_/A sky130_fd_sc_hd__o21a_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23605_ _23637_/CLK _23605_/D vssd1 vssd1 vccd1 vccd1 _23605_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20817_ _20817_/A vssd1 vssd1 vccd1 vccd1 _23759_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21797_ _21791_/A _21612_/X _21796_/Y _21581_/X vssd1 vssd1 vccd1 vccd1 _23926_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_179_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11550_ _13064_/A _11549_/X _11537_/X vssd1 vssd1 vccd1 vccd1 _11550_/X sky130_fd_sc_hd__o21a_1
XFILLER_169_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23536_ _23951_/A _23536_/D vssd1 vssd1 vccd1 vccd1 _23536_/Q sky130_fd_sc_hd__dfxtp_1
X_20748_ _23744_/Q _20729_/X _20747_/X _20737_/X vssd1 vssd1 vccd1 vccd1 _23744_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_329_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11481_ _22484_/Q _22644_/Q _22323_/Q _23459_/Q _11461_/X _11462_/X vssd1 vssd1 vccd1
+ vccd1 _11481_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23467_ _23467_/CLK _23467_/D vssd1 vssd1 vccd1 vccd1 _23467_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_326_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20679_ _23733_/Q _20667_/X _20678_/X _20673_/X vssd1 vssd1 vccd1 vccd1 _23733_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13220_ _22478_/Q _22638_/Q _22317_/Q _23453_/Q _13114_/A _13127_/A vssd1 vssd1 vccd1
+ vccd1 _13221_/B sky130_fd_sc_hd__mux4_1
XFILLER_183_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22418_ _23554_/CLK _22418_/D vssd1 vssd1 vccd1 vccd1 _22418_/Q sky130_fd_sc_hd__dfxtp_1
X_23398_ _23526_/CLK _23398_/D vssd1 vssd1 vccd1 vccd1 _23398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13151_ _13158_/A _13150_/X _11235_/A vssd1 vssd1 vccd1 vccd1 _13151_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_192_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22349_ _23515_/CLK _22349_/D vssd1 vssd1 vccd1 vccd1 _22349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_341_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12102_ _22370_/Q _22402_/Q _22691_/Q _23058_/Q _12094_/X _11457_/B vssd1 vssd1 vccd1
+ vccd1 _12102_/X sky130_fd_sc_hd__mux4_1
XFILLER_340_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13082_ _13082_/A _13082_/B vssd1 vssd1 vccd1 vccd1 _13083_/A sky130_fd_sc_hd__nor2_1
XFILLER_297_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12033_ _12998_/A _12033_/B vssd1 vssd1 vccd1 vccd1 _12033_/Y sky130_fd_sc_hd__nor2_1
X_16910_ _16910_/A vssd1 vssd1 vccd1 vccd1 _22550_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17890_ _17981_/A vssd1 vssd1 vccd1 vccd1 _17932_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16841_ _19191_/A vssd1 vssd1 vccd1 vccd1 _16841_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_293_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_293_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19560_ _23430_/Q _19169_/A _19566_/S vssd1 vssd1 vccd1 vccd1 _19561_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16772_ _16772_/A vssd1 vssd1 vccd1 vccd1 _22508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13984_ _13984_/A vssd1 vssd1 vccd1 vccd1 _13984_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18511_ _22999_/Q _18518_/B vssd1 vssd1 vccd1 vccd1 _18511_/Y sky130_fd_sc_hd__nand2_1
XFILLER_280_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15723_ _15723_/A _15723_/B vssd1 vssd1 vccd1 vccd1 _15723_/Y sky130_fd_sc_hd__nand2_4
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ _12919_/A _12934_/X _12687_/X vssd1 vssd1 vccd1 vccd1 _12935_/Y sky130_fd_sc_hd__o21ai_1
X_19491_ _19491_/A vssd1 vssd1 vccd1 vccd1 _23399_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ _22975_/Q _18438_/B _18441_/Y vssd1 vssd1 vccd1 vccd1 _22975_/D sky130_fd_sc_hd__o21a_1
XFILLER_234_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _15885_/A _15654_/B vssd1 vssd1 vccd1 vccd1 _15654_/Y sky130_fd_sc_hd__nand2_1
XFILLER_179_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12866_ _13029_/A _13028_/A vssd1 vssd1 vccd1 vccd1 _12868_/A sky130_fd_sc_hd__nor2_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_310_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _15219_/A vssd1 vssd1 vccd1 vccd1 _14605_/X sky130_fd_sc_hd__buf_2
X_18373_ _14989_/X _18375_/C _18372_/Y vssd1 vssd1 vccd1 vccd1 _22951_/D sky130_fd_sc_hd__o21a_1
XFILLER_221_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11817_ _12316_/A _11817_/B vssd1 vssd1 vccd1 vccd1 _11817_/X sky130_fd_sc_hd__or2_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _14264_/X _15542_/X _15584_/X _12665_/A vssd1 vssd1 vccd1 vccd1 _15585_/X
+ sky130_fd_sc_hd__o22a_1
X_12797_ _12797_/A vssd1 vssd1 vccd1 vccd1 _12797_/X sky130_fd_sc_hd__buf_2
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17324_ _17324_/A vssd1 vssd1 vccd1 vccd1 _17324_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14536_ _14535_/X _16942_/A _14539_/S vssd1 vssd1 vccd1 vccd1 _19090_/B sky130_fd_sc_hd__mux2_2
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11748_ _11736_/Y _11739_/Y _11744_/Y _11747_/Y _11275_/A vssd1 vssd1 vccd1 vccd1
+ _11761_/B sky130_fd_sc_hd__o221a_1
XFILLER_187_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_335_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17255_ _17255_/A vssd1 vssd1 vccd1 vccd1 _17255_/X sky130_fd_sc_hd__clkbuf_2
X_14467_ _14446_/B _14467_/B _14467_/C vssd1 vssd1 vccd1 vccd1 _14468_/B sky130_fd_sc_hd__nand3b_4
XFILLER_146_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_329_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11679_ _11679_/A vssd1 vssd1 vccd1 vccd1 _11680_/A sky130_fd_sc_hd__clkbuf_4
X_16206_ _19555_/A _19091_/A vssd1 vssd1 vccd1 vccd1 _16288_/A sky130_fd_sc_hd__nor2_4
XFILLER_317_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13418_ _13427_/A _13427_/B _15090_/A vssd1 vssd1 vccd1 vccd1 _13428_/A sky130_fd_sc_hd__o21a_1
X_17186_ _17180_/X _17184_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17186_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_344_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14398_ _21077_/D _21320_/A _20191_/A vssd1 vssd1 vccd1 vccd1 _14467_/B sky130_fd_sc_hd__mux2_2
XFILLER_289_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_350_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16137_ _23683_/Q _16137_/B vssd1 vssd1 vccd1 vccd1 _16137_/X sky130_fd_sc_hd__or2_1
XFILLER_127_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_344_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13349_ _13349_/A _13349_/B _13611_/A vssd1 vssd1 vccd1 vccd1 _13350_/B sky130_fd_sc_hd__and3_1
XFILLER_288_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_303_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16068_ _23713_/Q _15592_/X _16067_/X vssd1 vssd1 vccd1 vccd1 _16068_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15019_ _15456_/B _15018_/X _15538_/A vssd1 vssd1 vccd1 vccd1 _15019_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19827_ _19827_/A vssd1 vssd1 vccd1 vccd1 _23549_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_256_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19758_ _19758_/A vssd1 vssd1 vccd1 vccd1 _23518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18709_ _18709_/A vssd1 vssd1 vccd1 vccd1 _23081_/D sky130_fd_sc_hd__clkbuf_1
X_19689_ _19252_/X _23488_/Q _19693_/S vssd1 vssd1 vccd1 vccd1 _19690_/A sky130_fd_sc_hd__mux2_1
XFILLER_253_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21720_ _21720_/A _21865_/A vssd1 vssd1 vccd1 vccd1 _21720_/X sky130_fd_sc_hd__or2_1
XFILLER_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_342_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21651_ _21649_/Y _21650_/X _21840_/A vssd1 vssd1 vccd1 vccd1 _21653_/B sky130_fd_sc_hd__a21o_1
XFILLER_224_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20602_ _20602_/A vssd1 vssd1 vccd1 vccd1 _20602_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21582_ _13939_/B _21305_/X _21580_/X _21581_/X vssd1 vssd1 vccd1 vccd1 _23919_/D
+ sky130_fd_sc_hd__o211a_1
X_23321_ _23419_/CLK _23321_/D vssd1 vssd1 vccd1 vccd1 _23321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20533_ _20533_/A _20533_/B _20533_/C _21080_/A vssd1 vssd1 vccd1 vccd1 _20533_/Y
+ sky130_fd_sc_hd__nor4_4
XFILLER_177_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23252_ _23573_/CLK _23252_/D vssd1 vssd1 vccd1 vccd1 _23252_/Q sky130_fd_sc_hd__dfxtp_1
X_20464_ _23704_/Q _20416_/B _20463_/Y _20459_/X vssd1 vssd1 vccd1 vccd1 _23704_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_181_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_323_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22203_ _22216_/A _21867_/X _22202_/X _21865_/X vssd1 vssd1 vccd1 vccd1 _22205_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_192_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23183_ _23535_/CLK _23183_/D vssd1 vssd1 vccd1 vccd1 _23183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20395_ _17307_/A _20261_/X _20396_/B vssd1 vssd1 vccd1 vccd1 _20395_/Y sky130_fd_sc_hd__o21ai_1
XTAP_7306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_334_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22134_ _22134_/A _22134_/B vssd1 vssd1 vccd1 vccd1 _22136_/A sky130_fd_sc_hd__nor2_1
XTAP_7339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_315_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22065_ _22065_/A _22085_/B vssd1 vssd1 vccd1 vccd1 _22066_/B sky130_fd_sc_hd__nand2_1
XTAP_6649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput294 _13988_/Y vssd1 vssd1 vccd1 vccd1 addr1[0] sky130_fd_sc_hd__buf_2
XTAP_5915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_288_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_1 _22139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21016_ _23821_/Q _21028_/B vssd1 vssd1 vccd1 vccd1 _21016_/X sky130_fd_sc_hd__or2_1
XFILLER_310_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_290_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22967_ _22968_/CLK _22967_/D vssd1 vssd1 vccd1 vccd1 _22967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12720_ _12958_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _12720_/X sky130_fd_sc_hd__or2_1
XFILLER_16_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21918_ _21918_/A _21918_/B vssd1 vssd1 vccd1 vccd1 _21919_/B sky130_fd_sc_hd__nand2_1
XFILLER_215_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22898_ _23426_/CLK _22898_/D vssd1 vssd1 vccd1 vccd1 _22898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12651_ _12759_/A _12651_/B vssd1 vssd1 vccd1 vccd1 _12651_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21849_ _21849_/A vssd1 vssd1 vccd1 vccd1 _21849_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11602_ _11965_/A vssd1 vssd1 vccd1 vccd1 _12700_/A sky130_fd_sc_hd__buf_2
XFILLER_168_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12582_ _23401_/Q _23017_/Q _23369_/Q _23337_/Q _12314_/X _11815_/X vssd1 vssd1 vccd1
+ vccd1 _12582_/X sky130_fd_sc_hd__mux4_1
X_15370_ _11763_/Y _15048_/A _15368_/X _21676_/A _15321_/X vssd1 vssd1 vccd1 vccd1
+ _18808_/A sky130_fd_sc_hd__a32o_4
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14321_ _13521_/B _13022_/B _14330_/S vssd1 vssd1 vccd1 vccd1 _14321_/X sky130_fd_sc_hd__mux2_1
X_23519_ _23551_/CLK _23519_/D vssd1 vssd1 vccd1 vccd1 _23519_/Q sky130_fd_sc_hd__dfxtp_1
X_11533_ _11533_/A vssd1 vssd1 vccd1 vccd1 _13127_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_196_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17040_ _17276_/A vssd1 vssd1 vccd1 vccd1 _17084_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_317_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11464_ _21848_/A _11464_/B vssd1 vssd1 vccd1 vccd1 _11464_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14252_ _15460_/B vssd1 vssd1 vccd1 vccd1 _16054_/B sky130_fd_sc_hd__buf_2
XFILLER_333_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_319_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13203_ _23485_/Q _23581_/Q _22545_/Q _22349_/Q _13191_/S _13195_/X vssd1 vssd1 vccd1
+ vccd1 _13203_/X sky130_fd_sc_hd__mux4_1
X_11395_ _13427_/A vssd1 vssd1 vccd1 vccd1 _11396_/B sky130_fd_sc_hd__inv_2
XFILLER_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14183_ _14385_/A _14385_/B vssd1 vssd1 vccd1 vccd1 _14800_/A sky130_fd_sc_hd__nor2_2
XFILLER_325_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_2_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_13134_ _13126_/Y _13129_/Y _13131_/Y _13133_/Y _11379_/A vssd1 vssd1 vccd1 vccd1
+ _13134_/X sky130_fd_sc_hd__o221a_1
X_18991_ _18991_/A vssd1 vssd1 vccd1 vccd1 _23192_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_298_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17942_ _22825_/Q _17938_/X _17939_/X input271/X _17933_/X vssd1 vssd1 vccd1 vccd1
+ _17942_/X sky130_fd_sc_hd__a221o_1
X_13065_ _23424_/Q _23040_/Q _23392_/Q _23360_/Q _11517_/X _11519_/X vssd1 vssd1 vccd1
+ vccd1 _13065_/X sky130_fd_sc_hd__mux4_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12016_ _12852_/A _12015_/X _11285_/A vssd1 vssd1 vccd1 vccd1 _12016_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_294_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17873_ _17873_/A vssd1 vssd1 vccd1 vccd1 _22807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19612_ _19612_/A vssd1 vssd1 vccd1 vccd1 _19621_/S sky130_fd_sc_hd__buf_6
X_16824_ _16824_/A vssd1 vssd1 vccd1 vccd1 _22523_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_293_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19543_ _19249_/X _23423_/Q _19549_/S vssd1 vssd1 vccd1 vccd1 _19544_/A sky130_fd_sc_hd__mux2_1
XFILLER_253_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16755_ _22504_/Q _16747_/X _16748_/X input18/X vssd1 vssd1 vccd1 vccd1 _16756_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13967_ _13967_/A _13967_/B vssd1 vssd1 vccd1 vccd1 _13968_/A sky130_fd_sc_hd__and2_1
XFILLER_207_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15706_ _15671_/X _15672_/X _15704_/X _15705_/X vssd1 vssd1 vccd1 vccd1 _15706_/X
+ sky130_fd_sc_hd__o22a_2
X_19474_ _19474_/A vssd1 vssd1 vccd1 vccd1 _23392_/D sky130_fd_sc_hd__clkbuf_1
X_12918_ _22797_/Q _22765_/Q _22666_/Q _22733_/Q _12825_/X _12685_/X vssd1 vssd1 vccd1
+ vccd1 _12919_/B sky130_fd_sc_hd__mux4_2
XFILLER_0_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16686_ input9/X vssd1 vssd1 vccd1 vccd1 _16691_/A sky130_fd_sc_hd__inv_2
XFILLER_206_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13898_ _21293_/A vssd1 vssd1 vccd1 vccd1 _13931_/A sky130_fd_sc_hd__buf_2
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18425_ _18427_/A _18427_/C _18424_/Y vssd1 vssd1 vccd1 vccd1 _22969_/D sky130_fd_sc_hd__o21a_1
X_15637_ _13608_/Y _16031_/S _15635_/Y _15636_/X vssd1 vssd1 vccd1 vccd1 _15637_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _12897_/A _12849_/B vssd1 vssd1 vccd1 vccd1 _12849_/X sky130_fd_sc_hd__or2_1
XFILLER_181_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18356_ _16168_/A _18357_/C _22946_/Q vssd1 vssd1 vccd1 vccd1 _18358_/B sky130_fd_sc_hd__a21oi_1
XFILLER_222_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ _14210_/X _21791_/B _15567_/X vssd1 vssd1 vccd1 vccd1 _18820_/A sky130_fd_sc_hd__o21a_4
XFILLER_203_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_348_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17307_ _17307_/A vssd1 vssd1 vccd1 vccd1 _17307_/Y sky130_fd_sc_hd__inv_2
X_14519_ _14431_/X _14442_/X _14505_/X _14514_/X _14518_/X vssd1 vssd1 vccd1 vccd1
+ _14520_/B sky130_fd_sc_hd__o32a_4
XFILLER_336_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18287_ _18315_/A _18287_/B _18287_/C vssd1 vssd1 vccd1 vccd1 _22922_/D sky130_fd_sc_hd__nor3_1
X_15499_ _22960_/Q vssd1 vssd1 vccd1 vccd1 _15501_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_175_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17238_ _17167_/A _17228_/X _17236_/X _17237_/X vssd1 vssd1 vccd1 vccd1 _17238_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_190_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_305_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17169_ _17169_/A vssd1 vssd1 vccd1 vccd1 _17169_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_305_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_288_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_289_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20180_ _14756_/X _20154_/X _20179_/X vssd1 vssd1 vccd1 vccd1 _20180_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_331_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_304_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23870_ _23918_/CLK _23870_/D vssd1 vssd1 vccd1 vccd1 _23870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22821_ _23551_/CLK _22821_/D vssd1 vssd1 vccd1 vccd1 _22821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22752_ _23048_/CLK _22752_/D vssd1 vssd1 vccd1 vccd1 _22752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21703_ _21703_/A _21703_/B vssd1 vssd1 vccd1 vccd1 _21705_/A sky130_fd_sc_hd__nor2_1
X_22683_ _23564_/CLK _22683_/D vssd1 vssd1 vccd1 vccd1 _22683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_358_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21634_ _21634_/A vssd1 vssd1 vccd1 vccd1 _22215_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_339_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_139_wb_clk_i _22712_/CLK vssd1 vssd1 vccd1 vccd1 _23696_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21565_ _21533_/A _21535_/B _21533_/B vssd1 vssd1 vccd1 vccd1 _21566_/B sky130_fd_sc_hd__a21boi_4
XFILLER_197_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23304_ _23496_/CLK _23304_/D vssd1 vssd1 vccd1 vccd1 _23304_/Q sky130_fd_sc_hd__dfxtp_1
X_20516_ _23706_/Q _20517_/B _20516_/C vssd1 vssd1 vccd1 vccd1 _20520_/A sky130_fd_sc_hd__and3_1
XFILLER_315_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21496_ _21496_/A _21496_/B vssd1 vssd1 vccd1 vccd1 _21496_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_193_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23235_ _23459_/CLK _23235_/D vssd1 vssd1 vccd1 vccd1 _23235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20447_ _20467_/A vssd1 vssd1 vccd1 vccd1 _20447_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_326_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23166_ _23550_/CLK _23166_/D vssd1 vssd1 vccd1 vccd1 _23166_/Q sky130_fd_sc_hd__dfxtp_1
X_11180_ _12983_/A vssd1 vssd1 vccd1 vccd1 _13091_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_180_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20378_ _20174_/X _20375_/X _20376_/Y _22140_/B _20147_/X vssd1 vssd1 vccd1 vccd1
+ _21177_/A sky130_fd_sc_hd__o32a_4
XTAP_7136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22117_ _22065_/A _22085_/Y _22116_/Y _22087_/Y vssd1 vssd1 vccd1 vccd1 _22118_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_7169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23097_ _23100_/CLK _23097_/D vssd1 vssd1 vccd1 vccd1 _23097_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22048_ _22048_/A vssd1 vssd1 vccd1 vccd1 _22048_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14870_ _23656_/Q _15353_/B vssd1 vssd1 vccd1 vccd1 _14870_/X sky130_fd_sc_hd__or2_1
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_290_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13821_ _13821_/A _14019_/C vssd1 vssd1 vccd1 vccd1 _13821_/Y sky130_fd_sc_hd__nor2_1
XFILLER_291_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16540_ _14706_/X _22423_/Q _16546_/S vssd1 vssd1 vccd1 vccd1 _16541_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13752_ _13752_/A _14089_/A _13777_/B vssd1 vssd1 vccd1 vccd1 _13847_/A sky130_fd_sc_hd__or3_4
XINSDIODE2_108 _13521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_119 _20217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12703_ _11218_/A _12689_/X _12702_/X _11124_/A vssd1 vssd1 vccd1 vccd1 _12704_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_243_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_349_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16471_ _16528_/S vssd1 vssd1 vccd1 vccd1 _16480_/S sky130_fd_sc_hd__buf_6
X_13683_ _14833_/A vssd1 vssd1 vccd1 vccd1 _15830_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18210_ _22896_/Q _18214_/B vssd1 vssd1 vccd1 vccd1 _18210_/X sky130_fd_sc_hd__or2_1
XFILLER_204_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15422_ _19204_/A vssd1 vssd1 vccd1 vccd1 _15422_/X sky130_fd_sc_hd__clkbuf_2
XPHY_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12634_ _12634_/A _12634_/B _12634_/C vssd1 vssd1 vccd1 vccd1 _12634_/Y sky130_fd_sc_hd__nor3_4
XFILLER_203_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19190_ _19190_/A vssd1 vssd1 vccd1 vccd1 _23276_/D sky130_fd_sc_hd__clkbuf_1
XPHY_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18141_ _22893_/Q _18163_/A vssd1 vssd1 vccd1 vccd1 _18167_/A sky130_fd_sc_hd__nand2_1
XFILLER_15_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15353_ _23664_/Q _15353_/B vssd1 vssd1 vccd1 vccd1 _15353_/X sky130_fd_sc_hd__or2_1
XPHY_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12565_ _12565_/A _12565_/B vssd1 vssd1 vccd1 vccd1 _12565_/X sky130_fd_sc_hd__or2_1
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_357_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14304_ _13521_/B _13022_/B _14348_/A vssd1 vssd1 vccd1 vccd1 _14304_/X sky130_fd_sc_hd__mux2_1
XFILLER_346_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18072_ _22861_/Q _18067_/X _18068_/X _22994_/Q _18069_/X vssd1 vssd1 vccd1 vccd1
+ _18072_/X sky130_fd_sc_hd__a221o_1
X_11516_ _13216_/A vssd1 vssd1 vccd1 vccd1 _13064_/A sky130_fd_sc_hd__buf_2
X_15284_ _15283_/X _22270_/Q _15284_/S vssd1 vssd1 vccd1 vccd1 _15285_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12496_ _13506_/B vssd1 vssd1 vccd1 vccd1 _14672_/B sky130_fd_sc_hd__buf_4
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17023_ _17047_/A vssd1 vssd1 vccd1 vccd1 _17283_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_144_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14235_ _14235_/A vssd1 vssd1 vccd1 vccd1 _14235_/X sky130_fd_sc_hd__buf_2
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11447_ _23235_/Q _23203_/Q _23171_/Q _23139_/Q _13032_/S _11169_/A vssd1 vssd1 vccd1
+ vccd1 _11448_/B sky130_fd_sc_hd__mux4_1
XFILLER_236_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_298_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_298_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11378_ _11378_/A vssd1 vssd1 vccd1 vccd1 _11379_/A sky130_fd_sc_hd__clkbuf_4
X_14166_ _14553_/A _14552_/A vssd1 vssd1 vccd1 vccd1 _20140_/B sky130_fd_sc_hd__nand2_2
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13117_ _13117_/A _13117_/B vssd1 vssd1 vccd1 vccd1 _13117_/Y sky130_fd_sc_hd__nor2_1
X_18974_ _18974_/A vssd1 vssd1 vccd1 vccd1 _23184_/D sky130_fd_sc_hd__clkbuf_1
X_14097_ _14097_/A vssd1 vssd1 vccd1 vccd1 _14097_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_301_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17925_ _17991_/A vssd1 vssd1 vccd1 vccd1 _17987_/S sky130_fd_sc_hd__clkbuf_2
X_13048_ _23424_/Q _23040_/Q _23392_/Q _23360_/Q _13088_/S _13037_/X vssd1 vssd1 vccd1
+ vccd1 _13048_/X sky130_fd_sc_hd__mux4_1
XFILLER_267_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_310_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17856_ _17856_/A vssd1 vssd1 vccd1 vccd1 _22799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16807_ _13777_/A _13934_/A _13457_/A vssd1 vssd1 vccd1 vccd1 _16808_/D sky130_fd_sc_hd__o21ai_1
XFILLER_226_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17787_ _22769_/Q _17623_/X _17787_/S vssd1 vssd1 vccd1 vccd1 _17788_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14999_ _14989_/X _14998_/X _15885_/A vssd1 vssd1 vccd1 vccd1 _14999_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19526_ _19526_/A vssd1 vssd1 vccd1 vccd1 _23415_/D sky130_fd_sc_hd__clkbuf_1
X_16738_ _16741_/A _16738_/B vssd1 vssd1 vccd1 vccd1 _16739_/A sky130_fd_sc_hd__or2_1
XFILLER_223_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19457_ _19468_/A vssd1 vssd1 vccd1 vccd1 _19466_/S sky130_fd_sc_hd__buf_2
X_16669_ _22481_/Q _16294_/X _16673_/S vssd1 vssd1 vccd1 vccd1 _16670_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18408_ _15644_/A _18409_/C _22964_/Q vssd1 vssd1 vccd1 vccd1 _18410_/B sky130_fd_sc_hd__a21oi_1
X_19388_ _23354_/Q _18840_/X _19394_/S vssd1 vssd1 vccd1 vccd1 _19389_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18339_ _15950_/X _18341_/C _18338_/Y vssd1 vssd1 vccd1 vccd1 _22939_/D sky130_fd_sc_hd__o21a_1
XFILLER_300_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21350_ _21351_/A _21350_/B vssd1 vssd1 vccd1 vccd1 _21403_/A sky130_fd_sc_hd__and2_1
XFILLER_337_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_336_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20301_ _20272_/X _20675_/A _20300_/X _20285_/X vssd1 vssd1 vccd1 vccd1 _23669_/D
+ sky130_fd_sc_hd__o211a_1
X_21281_ _21281_/A vssd1 vssd1 vccd1 vccd1 _21281_/X sky130_fd_sc_hd__buf_4
XFILLER_135_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23020_ _23950_/A _23020_/D vssd1 vssd1 vccd1 vccd1 _23020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_351_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20232_ _20323_/A _21013_/A vssd1 vssd1 vccd1 vccd1 _20232_/Y sky130_fd_sc_hd__nand2_1
XFILLER_293_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_289_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_320_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20163_ _23653_/Q _20379_/A vssd1 vssd1 vccd1 vccd1 _20163_/X sky130_fd_sc_hd__or2_1
XFILLER_226_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_304_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20094_ _20098_/C _20098_/D _23639_/Q vssd1 vssd1 vccd1 vccd1 _20096_/B sky130_fd_sc_hd__a21oi_1
XFILLER_69_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23922_ _23935_/CLK _23922_/D vssd1 vssd1 vccd1 vccd1 _23922_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_285_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23853_ _23856_/CLK _23853_/D vssd1 vssd1 vccd1 vccd1 _23853_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22804_ _23391_/CLK _22804_/D vssd1 vssd1 vccd1 vccd1 _22804_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_309_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20996_ _20996_/A _20996_/B vssd1 vssd1 vccd1 vccd1 _20996_/Y sky130_fd_sc_hd__nand2_1
X_23784_ _23911_/CLK _23784_/D vssd1 vssd1 vccd1 vccd1 _23784_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22735_ _22801_/CLK _22735_/D vssd1 vssd1 vccd1 vccd1 _22735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_347_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22666_ _22666_/CLK _22666_/D vssd1 vssd1 vccd1 vccd1 _22666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21617_ _14195_/X _21518_/X _21868_/A _15318_/B vssd1 vssd1 vccd1 vccd1 _21617_/X
+ sky130_fd_sc_hd__a211o_1
X_22597_ _22974_/CLK _22597_/D vssd1 vssd1 vccd1 vccd1 _22597_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_21_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ _12350_/A _12350_/B vssd1 vssd1 vccd1 vccd1 _12350_/Y sky130_fd_sc_hd__nand2_1
XFILLER_354_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21548_ _21548_/A _21548_/B vssd1 vssd1 vccd1 vccd1 _21559_/A sky130_fd_sc_hd__nor2_2
XFILLER_127_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11301_ _23894_/Q vssd1 vssd1 vccd1 vccd1 _12475_/A sky130_fd_sc_hd__buf_4
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12281_ _12274_/Y _12276_/Y _12278_/Y _12280_/Y _11826_/A vssd1 vssd1 vccd1 vccd1
+ _12282_/C sky130_fd_sc_hd__o221a_1
XFILLER_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21479_ _21479_/A vssd1 vssd1 vccd1 vccd1 _21479_/X sky130_fd_sc_hd__clkbuf_4
X_11232_ _11232_/A vssd1 vssd1 vccd1 vccd1 _11233_/A sky130_fd_sc_hd__buf_2
X_14020_ input243/X _14004_/X _14019_/X vssd1 vssd1 vccd1 vccd1 _14020_/X sky130_fd_sc_hd__a21o_4
X_23218_ _23538_/CLK _23218_/D vssd1 vssd1 vccd1 vccd1 _23218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_323_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_323_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_296_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11163_ _11163_/A vssd1 vssd1 vccd1 vccd1 _11953_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_310_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23149_ _23407_/CLK _23149_/D vssd1 vssd1 vccd1 vccd1 _23149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_36_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23448_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_350_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_311_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15971_ _23003_/Q _16084_/A _16085_/A input232/X vssd1 vssd1 vccd1 vccd1 _22087_/B
+ sky130_fd_sc_hd__a22o_4
X_11094_ _23893_/Q _23892_/Q vssd1 vssd1 vccd1 vccd1 _15081_/B sky130_fd_sc_hd__nand2_2
XTAP_6265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17710_ _17710_/A vssd1 vssd1 vccd1 vccd1 _22734_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14922_ _14922_/A vssd1 vssd1 vccd1 vccd1 _14923_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18690_ _18690_/A vssd1 vssd1 vccd1 vccd1 _23073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17641_ _17641_/A vssd1 vssd1 vccd1 vccd1 _22707_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14853_ _14644_/X _14646_/X _14853_/S vssd1 vssd1 vccd1 vccd1 _14853_/X sky130_fd_sc_hd__mux2_1
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_291_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _12704_/B _13798_/B _13781_/A vssd1 vssd1 vccd1 vccd1 _13804_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17572_ _18798_/A vssd1 vssd1 vccd1 vccd1 _17572_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_302_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14784_ _14784_/A vssd1 vssd1 vccd1 vccd1 _14784_/Y sky130_fd_sc_hd__inv_2
X_11996_ _22792_/Q _22760_/Q _22661_/Q _22728_/Q _12716_/A _11669_/X vssd1 vssd1 vccd1
+ vccd1 _11997_/B sky130_fd_sc_hd__mux4_1
XFILLER_205_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19311_ _19226_/X _23320_/Q _19311_/S vssd1 vssd1 vccd1 vccd1 _19312_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16523_ _16523_/A vssd1 vssd1 vccd1 vccd1 _22417_/D sky130_fd_sc_hd__clkbuf_1
X_13735_ _14216_/B vssd1 vssd1 vccd1 vccd1 _13736_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_232_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19242_ _19242_/A vssd1 vssd1 vccd1 vccd1 _19242_/X sky130_fd_sc_hd__clkbuf_2
X_16454_ _16454_/A vssd1 vssd1 vccd1 vccd1 _22387_/D sky130_fd_sc_hd__clkbuf_1
X_13666_ _13993_/A _14069_/B _14002_/A vssd1 vssd1 vccd1 vccd1 _13666_/X sky130_fd_sc_hd__o21a_4
XFILLER_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15405_ _15735_/A _15405_/B vssd1 vssd1 vccd1 vccd1 _15405_/Y sky130_fd_sc_hd__nand2_1
X_12617_ _23413_/Q _23029_/Q _23381_/Q _23349_/Q _12013_/X _12710_/A vssd1 vssd1 vccd1
+ vccd1 _12617_/X sky130_fd_sc_hd__mux4_2
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19173_ _19172_/X _23271_/Q _19179_/S vssd1 vssd1 vccd1 vccd1 _19174_/A sky130_fd_sc_hd__mux2_1
X_16385_ _19267_/A _18625_/B vssd1 vssd1 vccd1 vccd1 _16442_/A sky130_fd_sc_hd__or2_4
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ _13532_/A _13612_/A _13538_/B vssd1 vssd1 vccd1 vccd1 _13629_/B sky130_fd_sc_hd__a21o_2
XFILLER_157_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18124_ _18116_/A _14107_/X _22879_/Q vssd1 vssd1 vccd1 vccd1 _18124_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15336_ _13393_/Y _14940_/B _15335_/Y _15010_/A vssd1 vssd1 vccd1 vccd1 _15336_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_247_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12548_ _14687_/A _14687_/B _12547_/X vssd1 vssd1 vccd1 vccd1 _13358_/B sky130_fd_sc_hd__a21oi_2
XFILLER_8_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_346_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_318_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18055_ _22855_/Q _18052_/X _18053_/X _22988_/Q _18054_/X vssd1 vssd1 vccd1 vccd1
+ _18055_/X sky130_fd_sc_hd__a221o_1
X_15267_ _23694_/Q _15210_/X _15266_/X vssd1 vssd1 vccd1 vccd1 _15267_/X sky130_fd_sc_hd__o21a_2
XFILLER_172_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12479_ _23302_/Q _23270_/Q _23238_/Q _23526_/Q _12475_/X _12476_/X vssd1 vssd1 vccd1
+ vccd1 _12480_/B sky130_fd_sc_hd__mux4_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17006_ _13455_/Y _16932_/A _17022_/A vssd1 vssd1 vccd1 vccd1 _17006_/X sky130_fd_sc_hd__a21o_1
X_14218_ _14725_/A vssd1 vssd1 vccd1 vccd1 _14218_/X sky130_fd_sc_hd__clkbuf_2
X_15198_ _15198_/A _15198_/B vssd1 vssd1 vccd1 vccd1 _15198_/X sky130_fd_sc_hd__or2_1
XFILLER_302_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_342_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14149_ _16971_/B _16966_/A vssd1 vssd1 vccd1 vccd1 _16917_/A sky130_fd_sc_hd__or2_1
XFILLER_301_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18957_ _16828_/X _23177_/Q _18957_/S vssd1 vssd1 vccd1 vccd1 _18958_/A sky130_fd_sc_hd__mux2_1
XFILLER_343_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17908_ _17908_/A _18097_/A vssd1 vssd1 vccd1 vccd1 _17908_/X sky130_fd_sc_hd__or2_1
XFILLER_267_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_295_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18888_ _23146_/Q _18788_/X _18896_/S vssd1 vssd1 vccd1 vccd1 _18889_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17839_ _17861_/A vssd1 vssd1 vccd1 vccd1 _17848_/S sky130_fd_sc_hd__buf_4
XFILLER_255_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20850_ _20850_/A vssd1 vssd1 vccd1 vccd1 _23768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19509_ _19509_/A vssd1 vssd1 vccd1 vccd1 _23407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20781_ _20781_/A vssd1 vssd1 vccd1 vccd1 _20781_/Y sky130_fd_sc_hd__inv_2
XFILLER_288_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_450 _21871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_461 _20708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_472 _13803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22520_ _22520_/CLK _22520_/D vssd1 vssd1 vccd1 vccd1 _22520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_483 _13979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_288_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_494 _14097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_298_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22451_ _23522_/CLK _22451_/D vssd1 vssd1 vccd1 vccd1 _22451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21402_ _13895_/A _21350_/B _21319_/A _21348_/Y _21318_/A vssd1 vssd1 vccd1 vccd1
+ _21403_/B sky130_fd_sc_hd__o221a_1
X_22382_ _23583_/CLK _22382_/D vssd1 vssd1 vccd1 vccd1 _22382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_309_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21333_ _21333_/A _21333_/B vssd1 vssd1 vccd1 vccd1 _21333_/X sky130_fd_sc_hd__and2_1
XFILLER_108_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_351_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21264_ _21077_/B _21196_/X _21263_/X vssd1 vssd1 vccd1 vccd1 _23901_/D sky130_fd_sc_hd__o21ba_2
XFILLER_2_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_351_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_305_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_333_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23003_ _23005_/CLK _23003_/D vssd1 vssd1 vccd1 vccd1 _23003_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_278_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20215_ _20254_/A vssd1 vssd1 vccd1 vccd1 _20215_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_278_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21195_ _21214_/S vssd1 vssd1 vccd1 vccd1 _21283_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20146_ _20213_/A vssd1 vssd1 vccd1 vccd1 _20146_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20077_ _23633_/Q _20085_/C _23634_/Q vssd1 vssd1 vccd1 vccd1 _20080_/B sky130_fd_sc_hd__a21oi_1
XFILLER_286_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23905_ _23907_/CLK _23905_/D vssd1 vssd1 vccd1 vccd1 _23905_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23836_ _23876_/CLK _23836_/D vssd1 vssd1 vccd1 vccd1 _23836_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _23406_/Q _23022_/Q _23374_/Q _23342_/Q _11719_/A _12246_/A vssd1 vssd1 vccd1
+ vccd1 _11850_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_154_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23755_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11781_ _11582_/A _11779_/X _11780_/X vssd1 vssd1 vccd1 vccd1 _11781_/Y sky130_fd_sc_hd__o21ai_1
X_23767_ _23768_/CLK _23767_/D vssd1 vssd1 vccd1 vccd1 _23767_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20979_ _23809_/Q _20969_/X _20977_/X _20978_/X vssd1 vssd1 vccd1 vccd1 _23809_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_260_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13520_ _13935_/B _13935_/C _13518_/Y _13935_/A _13646_/A vssd1 vssd1 vccd1 vccd1
+ _13621_/B sky130_fd_sc_hd__a2111o_1
XFILLER_201_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22718_ _23048_/CLK _22718_/D vssd1 vssd1 vccd1 vccd1 _22718_/Q sky130_fd_sc_hd__dfxtp_1
X_23698_ _23704_/CLK _23698_/D vssd1 vssd1 vccd1 vccd1 _23698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_347_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_348_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13451_ _13451_/A vssd1 vssd1 vccd1 vccd1 _20533_/C sky130_fd_sc_hd__clkbuf_4
X_22649_ _23048_/CLK _22649_/D vssd1 vssd1 vccd1 vccd1 _22649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12402_ _23399_/Q _23015_/Q _23367_/Q _23335_/Q _11920_/X _11652_/A vssd1 vssd1 vccd1
+ vccd1 _12402_/X sky130_fd_sc_hd__mux4_2
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16170_ _23684_/Q _16170_/B vssd1 vssd1 vccd1 vccd1 _16170_/X sky130_fd_sc_hd__or2_1
XFILLER_356_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_316_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13382_ _13948_/A _13382_/B _13382_/C vssd1 vssd1 vccd1 vccd1 _13383_/B sky130_fd_sc_hd__and3_1
XFILLER_154_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15121_ _14724_/A _15176_/C _15113_/Y _15120_/X vssd1 vssd1 vccd1 vccd1 _15121_/X
+ sky130_fd_sc_hd__a211o_4
X_12333_ _23402_/Q _23018_/Q _23370_/Q _23338_/Q _11920_/A _12329_/A vssd1 vssd1 vccd1
+ vccd1 _12334_/B sky130_fd_sc_hd__mux4_1
XFILLER_182_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15052_ input138/X input167/X _15052_/S vssd1 vssd1 vccd1 vccd1 _15052_/X sky130_fd_sc_hd__mux2_8
XFILLER_142_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12264_ _12401_/A _12264_/B vssd1 vssd1 vccd1 vccd1 _12264_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14003_ _14041_/A vssd1 vssd1 vccd1 vccd1 _14058_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11215_ _11215_/A vssd1 vssd1 vccd1 vccd1 _11216_/A sky130_fd_sc_hd__buf_6
X_12195_ _12565_/A _12194_/X _11844_/X vssd1 vssd1 vccd1 vccd1 _12195_/Y sky130_fd_sc_hd__o21ai_1
X_19860_ _19860_/A vssd1 vssd1 vccd1 vccd1 _23563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_268_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_323_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18811_ _18811_/A vssd1 vssd1 vccd1 vccd1 _18811_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_6040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11146_ _11146_/A vssd1 vssd1 vccd1 vccd1 _11699_/A sky130_fd_sc_hd__buf_4
XTAP_6051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19791_ _23533_/Q _19191_/A _19793_/S vssd1 vssd1 vccd1 vccd1 _19792_/A sky130_fd_sc_hd__mux2_1
XTAP_6062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18742_ _18742_/A vssd1 vssd1 vccd1 vccd1 _23096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_295_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15954_ _23678_/Q _16102_/B vssd1 vssd1 vccd1 vccd1 _15954_/X sky130_fd_sc_hd__or2_1
X_11077_ _14132_/A vssd1 vssd1 vccd1 vccd1 _13440_/A sky130_fd_sc_hd__buf_4
XTAP_6095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput150 dout1[49] vssd1 vssd1 vccd1 vccd1 input150/X sky130_fd_sc_hd__buf_2
XFILLER_295_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput161 dout1[59] vssd1 vssd1 vccd1 vccd1 input161/X sky130_fd_sc_hd__buf_2
XFILLER_283_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput172 irq[10] vssd1 vssd1 vccd1 vccd1 _20506_/C sky130_fd_sc_hd__buf_2
X_14905_ _14905_/A vssd1 vssd1 vccd1 vccd1 _14905_/X sky130_fd_sc_hd__buf_6
XFILLER_264_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18673_ _18673_/A vssd1 vssd1 vccd1 vccd1 _23065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15885_ _15885_/A _15885_/B vssd1 vssd1 vccd1 vccd1 _15885_/Y sky130_fd_sc_hd__nand2_1
XFILLER_236_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput183 irq[6] vssd1 vssd1 vccd1 vccd1 _20519_/C sky130_fd_sc_hd__buf_2
Xinput194 localMemory_wb_adr_i[13] vssd1 vssd1 vccd1 vccd1 input194/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_236_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17624_ _22702_/Q _17623_/X _17624_/S vssd1 vssd1 vccd1 vccd1 _17625_/A sky130_fd_sc_hd__mux2_1
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14836_ _14836_/A vssd1 vssd1 vccd1 vccd1 _15769_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _17555_/A vssd1 vssd1 vccd1 vccd1 _22680_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14767_ _14767_/A vssd1 vssd1 vccd1 vccd1 _14767_/X sky130_fd_sc_hd__clkbuf_2
X_11979_ _11217_/A _11967_/X _11978_/X _12660_/A vssd1 vssd1 vccd1 vccd1 _13875_/A
+ sky130_fd_sc_hd__a211oi_4
X_16506_ _16506_/A vssd1 vssd1 vccd1 vccd1 _22409_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13718_ _13718_/A _13718_/B _13718_/C _13718_/D vssd1 vssd1 vccd1 vccd1 _13810_/B
+ sky130_fd_sc_hd__and4_4
XFILLER_177_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17486_ _22651_/Q _16223_/X _17494_/S vssd1 vssd1 vccd1 vccd1 _17487_/A sky130_fd_sc_hd__mux2_1
XFILLER_338_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14698_ _15162_/A vssd1 vssd1 vccd1 vccd1 _14698_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19225_ _19225_/A vssd1 vssd1 vccd1 vccd1 _23287_/D sky130_fd_sc_hd__clkbuf_1
X_16437_ _16437_/A vssd1 vssd1 vccd1 vccd1 _22379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13649_ _13652_/A vssd1 vssd1 vccd1 vccd1 _13650_/A sky130_fd_sc_hd__buf_2
XFILLER_31_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_347_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19156_ _19156_/A vssd1 vssd1 vccd1 vccd1 _23265_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_353_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_319_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_318_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16368_ _16368_/A vssd1 vssd1 vccd1 vccd1 _16377_/S sky130_fd_sc_hd__buf_8
XFILLER_157_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18107_ _22873_/Q _18097_/X _18098_/X _23006_/Q _18099_/X vssd1 vssd1 vccd1 vccd1
+ _18107_/X sky130_fd_sc_hd__a221o_1
XFILLER_258_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15319_ _15161_/A _15314_/X _15318_/Y _15162_/X vssd1 vssd1 vccd1 vccd1 _15319_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_306_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19087_ _19087_/A vssd1 vssd1 vccd1 vccd1 _23235_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16299_ _16299_/A vssd1 vssd1 vccd1 vccd1 _22321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18038_ _18054_/A vssd1 vssd1 vccd1 vccd1 _18038_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20000_ _23613_/Q _19998_/B _19962_/X vssd1 vssd1 vccd1 vccd1 _20000_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_87_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19989_ _20027_/A _19994_/C vssd1 vssd1 vccd1 vccd1 _19989_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_287_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_286_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21951_ _21951_/A _21951_/B vssd1 vssd1 vccd1 vccd1 _21953_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20902_ _14713_/A _20894_/X _20577_/B _20897_/X vssd1 vssd1 vccd1 vccd1 _20902_/X
+ sky130_fd_sc_hd__a211o_1
X_21882_ _23831_/Q _23765_/Q vssd1 vssd1 vccd1 vccd1 _21884_/A sky130_fd_sc_hd__nor2_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23621_ _23624_/CLK _23621_/D vssd1 vssd1 vccd1 vccd1 _23621_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20833_ _20672_/B _20828_/X _20829_/X _23764_/Q vssd1 vssd1 vccd1 vccd1 _20834_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23552_ _23552_/CLK _23552_/D vssd1 vssd1 vccd1 vccd1 _23552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20764_ _23747_/Q _20628_/A _20762_/X _20763_/X vssd1 vssd1 vccd1 vccd1 _23747_/D
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_280 _15842_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_291 _18852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22503_ _23704_/CLK _22503_/D vssd1 vssd1 vccd1 vccd1 _22503_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_329_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23483_ _23515_/CLK _23483_/D vssd1 vssd1 vccd1 vccd1 _23483_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_168_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20695_ _20695_/A _20695_/B _20695_/C vssd1 vssd1 vccd1 vccd1 _20695_/X sky130_fd_sc_hd__or3_1
Xclkbuf_4_13_0_wb_clk_i clkbuf_3_6_1_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _22712_/CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_196_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22434_ _23505_/CLK _22434_/D vssd1 vssd1 vccd1 vccd1 _22434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_353_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22365_ _23565_/CLK _22365_/D vssd1 vssd1 vccd1 vccd1 _22365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_309_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_353_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_340_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21316_ _23912_/Q _21348_/B vssd1 vssd1 vccd1 vccd1 _21318_/A sky130_fd_sc_hd__nand2_1
X_22296_ _23368_/CLK _22296_/D vssd1 vssd1 vccd1 vccd1 _22296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_306_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_352_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21247_ _21258_/A _21247_/B vssd1 vssd1 vccd1 vccd1 _21248_/A sky130_fd_sc_hd__and2_1
XFILLER_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_334_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_313_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21178_ _21083_/A _20525_/A _21150_/X vssd1 vssd1 vccd1 vccd1 _21178_/X sky130_fd_sc_hd__a21o_1
XFILLER_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20129_ _23649_/Q _20127_/C _20128_/Y vssd1 vssd1 vccd1 vccd1 _23649_/D sky130_fd_sc_hd__a21oi_1
XFILLER_120_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _12745_/A _12944_/X _12946_/X _12950_/X vssd1 vssd1 vccd1 vccd1 _12951_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_274_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _23405_/Q _23021_/Q _23373_/Q _23341_/Q _11574_/A _11696_/X vssd1 vssd1 vccd1
+ vccd1 _11902_/X sky130_fd_sc_hd__mux4_2
X_15670_ _15670_/A vssd1 vssd1 vccd1 vccd1 _22278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _12886_/A _12882_/B vssd1 vssd1 vccd1 vccd1 _12882_/Y sky130_fd_sc_hd__nor2_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14621_ _14621_/A vssd1 vssd1 vccd1 vccd1 _15338_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23819_ _23824_/CLK _23819_/D vssd1 vssd1 vccd1 vccd1 _23819_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _23214_/Q _23182_/Q _23150_/Q _23118_/Q _11770_/A _11621_/A vssd1 vssd1 vccd1
+ vccd1 _11834_/B sky130_fd_sc_hd__mux4_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _17340_/A vssd1 vssd1 vccd1 vccd1 _22591_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14552_/A _14552_/B _14552_/C vssd1 vssd1 vccd1 vccd1 _14553_/C sky130_fd_sc_hd__or3_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _11763_/B _21648_/A _11763_/Y vssd1 vssd1 vccd1 vccd1 _11944_/A sky130_fd_sc_hd__o21a_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _14313_/A _13508_/B vssd1 vssd1 vccd1 vccd1 _13503_/Y sky130_fd_sc_hd__nand2_1
X_17271_ _21078_/A _17270_/X _17291_/S vssd1 vssd1 vccd1 vccd1 _17271_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14483_ _14483_/A _14595_/B vssd1 vssd1 vccd1 vccd1 _14918_/A sky130_fd_sc_hd__nor2_4
XFILLER_202_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11695_ _12241_/A vssd1 vssd1 vccd1 vccd1 _11698_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_329_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19010_ _16905_/X _23201_/Q _19012_/S vssd1 vssd1 vccd1 vccd1 _19011_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16222_ _16222_/A vssd1 vssd1 vccd1 vccd1 _22297_/D sky130_fd_sc_hd__clkbuf_1
X_13434_ _13434_/A vssd1 vssd1 vccd1 vccd1 _21077_/D sky130_fd_sc_hd__buf_8
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_328_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16153_ _16165_/B _16153_/B vssd1 vssd1 vccd1 vccd1 _16154_/B sky130_fd_sc_hd__nor2_2
X_13365_ _13897_/A _13358_/B _13364_/X vssd1 vssd1 vccd1 vccd1 _13366_/B sky130_fd_sc_hd__o21ai_1
XFILLER_316_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_51_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23505_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_315_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15104_ _19185_/A vssd1 vssd1 vccd1 vccd1 _15104_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_308_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ _12316_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _12316_/X sky130_fd_sc_hd__or2_1
XFILLER_343_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16084_ _16084_/A vssd1 vssd1 vccd1 vccd1 _16944_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_315_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13296_ _23939_/Q _13296_/B vssd1 vssd1 vccd1 vccd1 _13296_/X sky130_fd_sc_hd__or2_1
XFILLER_138_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_308_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15035_ _15032_/Y _15034_/X _15865_/A vssd1 vssd1 vccd1 vccd1 _15035_/X sky130_fd_sc_hd__mux2_4
X_19912_ _19912_/A vssd1 vssd1 vccd1 vccd1 _23587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12247_ _22783_/Q _22751_/Q _22652_/Q _22719_/Q _11413_/A _12425_/A vssd1 vssd1 vccd1
+ vccd1 _12247_/X sky130_fd_sc_hd__mux4_1
XFILLER_268_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_312_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19843_ _19843_/A _19843_/B vssd1 vssd1 vccd1 vccd1 _19900_/A sky130_fd_sc_hd__or2_4
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12178_ _12537_/S vssd1 vssd1 vccd1 vccd1 _12424_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_268_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11129_ _11713_/A vssd1 vssd1 vccd1 vccd1 _12371_/A sky130_fd_sc_hd__buf_6
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19774_ _23525_/Q _19163_/A _19782_/S vssd1 vssd1 vccd1 vccd1 _19775_/A sky130_fd_sc_hd__mux2_1
XFILLER_288_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16986_ _17033_/B vssd1 vssd1 vccd1 vccd1 _17174_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18725_ _18725_/A vssd1 vssd1 vccd1 vccd1 _23088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_329_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15937_ _15936_/X _22285_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15938_/A sky130_fd_sc_hd__mux2_1
XTAP_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18656_ _23058_/Q _17588_/X _18658_/S vssd1 vssd1 vccd1 vccd1 _18657_/A sky130_fd_sc_hd__mux2_1
X_15868_ _12868_/A _15996_/B _14259_/X _13495_/Y _15769_/A vssd1 vssd1 vccd1 vccd1
+ _15868_/X sky130_fd_sc_hd__a221o_1
XFILLER_97_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17607_ _18833_/A vssd1 vssd1 vccd1 vccd1 _17607_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14819_ _15318_/A vssd1 vssd1 vccd1 vccd1 _14819_/X sky130_fd_sc_hd__clkbuf_2
X_18587_ _18587_/A vssd1 vssd1 vccd1 vccd1 _23027_/D sky130_fd_sc_hd__clkbuf_1
X_15799_ _12916_/B _15582_/B _14259_/X _13493_/Y _15798_/Y vssd1 vssd1 vccd1 vccd1
+ _15799_/X sky130_fd_sc_hd__a221o_1
XFILLER_18_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17538_ _22675_/Q _16300_/X _17538_/S vssd1 vssd1 vccd1 vccd1 _17539_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17469_ _22645_/Q _16306_/X _17469_/S vssd1 vssd1 vccd1 vccd1 _17470_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_349_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19208_ _19207_/X _23282_/Q _19211_/S vssd1 vssd1 vccd1 vccd1 _19209_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20480_ _21173_/A _20482_/B vssd1 vssd1 vccd1 vccd1 _20480_/Y sky130_fd_sc_hd__nand2_1
XFILLER_121_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_335_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19139_ _19139_/A vssd1 vssd1 vccd1 vccd1 _23257_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22150_ _22148_/Y _22150_/B vssd1 vssd1 vccd1 vccd1 _22153_/A sky130_fd_sc_hd__and2b_1
XFILLER_336_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_307_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput410 _22564_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[11] sky130_fd_sc_hd__buf_2
Xoutput421 _22574_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[21] sky130_fd_sc_hd__buf_2
XFILLER_321_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_306_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21101_ _23848_/Q _21096_/X _21098_/X _20996_/A vssd1 vssd1 vccd1 vccd1 _21102_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xoutput432 _22584_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[31] sky130_fd_sc_hd__buf_2
X_22081_ _22081_/A _22081_/B vssd1 vssd1 vccd1 vccd1 _22082_/B sky130_fd_sc_hd__nor2_1
Xoutput443 _23943_/Q vssd1 vssd1 vccd1 vccd1 probe_errorCode[0] sky130_fd_sc_hd__buf_2
XTAP_6809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput454 _23879_/Q vssd1 vssd1 vccd1 vccd1 probe_opcode[0] sky130_fd_sc_hd__buf_2
Xoutput465 _23924_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[13] sky130_fd_sc_hd__buf_2
XFILLER_299_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput476 _23934_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[23] sky130_fd_sc_hd__buf_2
X_21032_ _20660_/A _21027_/X _21031_/X _21023_/X vssd1 vssd1 vccd1 vccd1 _23827_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_321_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput487 _23915_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[4] sky130_fd_sc_hd__buf_2
Xoutput498 _14075_/X vssd1 vssd1 vccd1 vccd1 wmask0[1] sky130_fd_sc_hd__buf_2
XFILLER_302_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_330_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_302_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_287_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22983_ _23424_/CLK _22983_/D vssd1 vssd1 vccd1 vccd1 _22983_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21934_ _21934_/A _21934_/B _21934_/C vssd1 vssd1 vccd1 vccd1 _22039_/A sky130_fd_sc_hd__and3_1
XFILLER_271_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_1_wb_clk_i clkbuf_2_3_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21865_ _21865_/A vssd1 vssd1 vccd1 vccd1 _21865_/X sky130_fd_sc_hd__buf_2
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23604_ _23652_/CLK _23604_/D vssd1 vssd1 vccd1 vccd1 _23604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20816_ _20825_/A _20816_/B vssd1 vssd1 vccd1 vccd1 _20817_/A sky130_fd_sc_hd__and2_1
XFILLER_249_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21796_ _22234_/A _21782_/X _21795_/X _21329_/X vssd1 vssd1 vccd1 vccd1 _21796_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_51_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_329_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23535_ _23535_/CLK _23535_/D vssd1 vssd1 vccd1 vccd1 _23535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20747_ _20757_/A _20747_/B _20747_/C vssd1 vssd1 vccd1 vccd1 _20747_/X sky130_fd_sc_hd__or3_1
XFILLER_169_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_345_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11480_ _15630_/A _11480_/B vssd1 vssd1 vccd1 vccd1 _11480_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23466_ _23466_/CLK _23466_/D vssd1 vssd1 vccd1 vccd1 _23466_/Q sky130_fd_sc_hd__dfxtp_4
X_20678_ _20695_/A _20678_/B _20678_/C vssd1 vssd1 vccd1 vccd1 _20678_/X sky130_fd_sc_hd__or3_1
XFILLER_338_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22417_ _23073_/CLK _22417_/D vssd1 vssd1 vccd1 vccd1 _22417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23397_ _23397_/CLK _23397_/D vssd1 vssd1 vccd1 vccd1 _23397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_325_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13150_ _22382_/Q _22414_/Q _22703_/Q _23070_/Q _13034_/S _13096_/X vssd1 vssd1 vccd1
+ vccd1 _13150_/X sky130_fd_sc_hd__mux4_2
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22348_ _23576_/CLK _22348_/D vssd1 vssd1 vccd1 vccd1 _22348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_313_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_312_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_297_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12101_ _12105_/A _12101_/B vssd1 vssd1 vccd1 vccd1 _12101_/X sky130_fd_sc_hd__or2_1
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13081_ _13249_/A _14276_/B vssd1 vssd1 vccd1 vccd1 _13082_/B sky130_fd_sc_hd__nor2_1
X_22279_ _23420_/CLK _22279_/D vssd1 vssd1 vccd1 vccd1 _22279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_340_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_340_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12032_ _22791_/Q _22759_/Q _22660_/Q _22727_/Q _12024_/X _12025_/X vssd1 vssd1 vccd1
+ vccd1 _12033_/B sky130_fd_sc_hd__mux4_1
XFILLER_137_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16840_ _16840_/A vssd1 vssd1 vccd1 vccd1 _22528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16771_ _16777_/A _16771_/B vssd1 vssd1 vccd1 vccd1 _16772_/A sky130_fd_sc_hd__or2_1
XFILLER_120_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13983_ _13983_/A _13985_/B vssd1 vssd1 vccd1 vccd1 _13984_/A sky130_fd_sc_hd__and2_2
XFILLER_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18510_ _18507_/X _18509_/Y _18503_/X vssd1 vssd1 vccd1 vccd1 _22998_/D sky130_fd_sc_hd__a21oi_1
XFILLER_281_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15722_ _15798_/A _15384_/X _15387_/X _14621_/A _15721_/Y vssd1 vssd1 vccd1 vccd1
+ _15723_/B sky130_fd_sc_hd__o221a_1
X_12934_ _23481_/Q _23577_/Q _22541_/Q _22345_/Q _12977_/S _12685_/X vssd1 vssd1 vccd1
+ vccd1 _12934_/X sky130_fd_sc_hd__mux4_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ _19172_/X _23399_/Q _19494_/S vssd1 vssd1 vccd1 vccd1 _19491_/A sky130_fd_sc_hd__mux2_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18441_ _18441_/A _18444_/B vssd1 vssd1 vccd1 vccd1 _18441_/Y sky130_fd_sc_hd__nor2_1
X_15653_ _14516_/A _15645_/X _15651_/Y _15652_/X vssd1 vssd1 vccd1 vccd1 _15654_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_206_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12865_ _12841_/Y _20347_/A _13500_/A vssd1 vssd1 vccd1 vccd1 _13028_/A sky130_fd_sc_hd__mux2_4
XFILLER_61_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _14916_/A vssd1 vssd1 vccd1 vccd1 _15219_/A sky130_fd_sc_hd__clkbuf_2
X_18372_ _14989_/X _18375_/C _18337_/X vssd1 vssd1 vccd1 vccd1 _18372_/Y sky130_fd_sc_hd__a21oi_1
X_11816_ _22271_/Q _23087_/Q _23503_/Q _22432_/Q _11814_/X _11815_/X vssd1 vssd1 vccd1
+ vccd1 _11817_/B sky130_fd_sc_hd__mux4_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15584_ _15582_/A _14942_/A _15582_/Y _15583_/X vssd1 vssd1 vccd1 vccd1 _15584_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _22472_/Q _22632_/Q _22311_/Q _23447_/Q _11308_/A _11320_/A vssd1 vssd1 vccd1
+ vccd1 _12796_/X sky130_fd_sc_hd__mux4_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _17322_/Y _16927_/B _16973_/X vssd1 vssd1 vccd1 vccd1 _22585_/D sky130_fd_sc_hd__a21oi_1
XFILLER_202_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _23890_/Q vssd1 vssd1 vccd1 vccd1 _14535_/X sky130_fd_sc_hd__buf_4
XFILLER_42_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _12139_/A _11746_/X _11284_/A vssd1 vssd1 vccd1 vccd1 _11747_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17254_ _22577_/Q _17199_/X _17240_/X _17253_/X vssd1 vssd1 vccd1 vccd1 _22577_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_169_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14466_ _14609_/A _14601_/A vssd1 vssd1 vccd1 vccd1 _14595_/B sky130_fd_sc_hd__or2_4
XFILLER_105_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_348_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11678_ _11678_/A vssd1 vssd1 vccd1 vccd1 _11679_/A sky130_fd_sc_hd__buf_4
XFILLER_335_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_317_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16205_ _19699_/B vssd1 vssd1 vccd1 vccd1 _19091_/A sky130_fd_sc_hd__buf_6
X_13417_ _20205_/A _20214_/A vssd1 vssd1 vccd1 vccd1 _15090_/A sky130_fd_sc_hd__nor2_2
X_17185_ _17250_/A vssd1 vssd1 vccd1 vccd1 _17235_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_190_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14397_ _22896_/Q _14394_/X _14164_/X _22589_/Q vssd1 vssd1 vccd1 vccd1 _21320_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_317_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16136_ _20034_/B _14901_/A _14902_/A _23651_/Q vssd1 vssd1 vccd1 vccd1 _16136_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_183_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ _13615_/A _13348_/B vssd1 vssd1 vccd1 vccd1 _13387_/B sky130_fd_sc_hd__xnor2_1
XFILLER_289_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_289_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16067_ _23841_/Q _15593_/X _16063_/X _16066_/X _14738_/X vssd1 vssd1 vccd1 vccd1
+ _16067_/X sky130_fd_sc_hd__a221o_1
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_332_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13279_ _23425_/Q _23041_/Q _23393_/Q _23361_/Q _11364_/A _11365_/A vssd1 vssd1 vccd1
+ vccd1 _13279_/X sky130_fd_sc_hd__mux4_1
XFILLER_170_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15018_ _15017_/Y _14655_/X _15018_/S vssd1 vssd1 vccd1 vccd1 _15018_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_303_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_312_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_312_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_296_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19826_ _23549_/Q _19242_/A _19826_/S vssd1 vssd1 vccd1 vccd1 _19827_/A sky130_fd_sc_hd__mux2_1
XFILLER_284_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_311_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_300_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19757_ _19245_/X _23518_/Q _19765_/S vssd1 vssd1 vccd1 vccd1 _19758_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16969_ _16939_/X _16948_/X _16951_/X _16965_/X _16968_/X vssd1 vssd1 vccd1 vccd1
+ _16969_/X sky130_fd_sc_hd__a221o_1
XFILLER_37_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18708_ _16828_/X _23081_/Q _18708_/S vssd1 vssd1 vccd1 vccd1 _18709_/A sky130_fd_sc_hd__mux2_1
XFILLER_351_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19688_ _19688_/A vssd1 vssd1 vccd1 vccd1 _23487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18639_ _23050_/Q _17562_/X _18647_/S vssd1 vssd1 vccd1 vccd1 _18640_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21650_ _14195_/X _21518_/X _21868_/A _15330_/Y vssd1 vssd1 vccd1 vccd1 _21650_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_342_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20601_ _20626_/A _20601_/B _20601_/C vssd1 vssd1 vccd1 vccd1 _20601_/X sky130_fd_sc_hd__or3_1
XFILLER_33_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21581_ _22122_/A vssd1 vssd1 vccd1 vccd1 _21581_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23320_ _23354_/CLK _23320_/D vssd1 vssd1 vccd1 vccd1 _23320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20532_ _20532_/A _20532_/B _20532_/C _20532_/D vssd1 vssd1 vccd1 vccd1 _21080_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_327_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_326_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23251_ _23510_/CLK _23251_/D vssd1 vssd1 vccd1 vccd1 _23251_/Q sky130_fd_sc_hd__dfxtp_1
X_20463_ _21153_/A _20463_/B vssd1 vssd1 vccd1 vccd1 _20463_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22202_ _20394_/A _22045_/X _16154_/B _22046_/X vssd1 vssd1 vccd1 vccd1 _22202_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_323_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23182_ _23502_/CLK _23182_/D vssd1 vssd1 vccd1 vccd1 _23182_/Q sky130_fd_sc_hd__dfxtp_1
X_20394_ _20394_/A _20394_/B vssd1 vssd1 vccd1 vccd1 _20396_/B sky130_fd_sc_hd__nand2_1
XTAP_7307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22133_ _22151_/A _23774_/Q vssd1 vssd1 vccd1 vccd1 _22134_/B sky130_fd_sc_hd__and2_1
XFILLER_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22064_ _22064_/A _22067_/A vssd1 vssd1 vccd1 vccd1 _22085_/B sky130_fd_sc_hd__or2_1
XFILLER_121_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput295 _13989_/Y vssd1 vssd1 vccd1 vccd1 addr1[1] sky130_fd_sc_hd__buf_2
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_287_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_2 _22139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21015_ _21051_/A vssd1 vssd1 vccd1 vccd1 _21028_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_287_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_290_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22966_ _22968_/CLK _22966_/D vssd1 vssd1 vccd1 vccd1 _22966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_255_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21917_ _23930_/Q _21920_/A vssd1 vssd1 vccd1 vccd1 _21918_/B sky130_fd_sc_hd__or2_1
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22897_ _23426_/CLK _22897_/D vssd1 vssd1 vccd1 vccd1 _22897_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_349_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12650_ _23317_/Q _23285_/Q _23253_/Q _23541_/Q _12751_/S _12671_/A vssd1 vssd1 vccd1
+ vccd1 _12651_/B sky130_fd_sc_hd__mux4_2
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21848_ _21848_/A _22048_/A vssd1 vssd1 vccd1 vccd1 _21848_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11601_ _11570_/Y _11577_/Y _11600_/X vssd1 vssd1 vccd1 vccd1 _11601_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_90_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12581_ _12586_/A _12581_/B vssd1 vssd1 vccd1 vccd1 _12581_/X sky130_fd_sc_hd__or2_1
X_21779_ _21779_/A _21779_/B vssd1 vssd1 vccd1 vccd1 _21799_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14320_ _13019_/Y _11939_/B _14329_/S vssd1 vssd1 vccd1 vccd1 _14320_/X sky130_fd_sc_hd__mux2_1
X_23518_ _23582_/CLK _23518_/D vssd1 vssd1 vccd1 vccd1 _23518_/Q sky130_fd_sc_hd__dfxtp_1
X_11532_ _11532_/A vssd1 vssd1 vccd1 vccd1 _11532_/X sky130_fd_sc_hd__buf_4
XFILLER_184_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_356_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14251_ _14251_/A vssd1 vssd1 vccd1 vccd1 _15460_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_345_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23449_ _23449_/CLK _23449_/D vssd1 vssd1 vccd1 vccd1 _23449_/Q sky130_fd_sc_hd__dfxtp_1
X_11463_ _22291_/Q _23107_/Q _23523_/Q _22452_/Q _11461_/X _11462_/X vssd1 vssd1 vccd1
+ vccd1 _11464_/B sky130_fd_sc_hd__mux4_1
XFILLER_137_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13202_ _13206_/A _13202_/B vssd1 vssd1 vccd1 vccd1 _13202_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_326_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14182_ _21335_/A _14524_/B _14370_/C vssd1 vssd1 vccd1 vccd1 _14385_/B sky130_fd_sc_hd__and3_2
XFILLER_319_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11394_ _11394_/A _14356_/B vssd1 vssd1 vccd1 vccd1 _13427_/A sky130_fd_sc_hd__and2_2
X_13133_ _13117_/A _13132_/X _11352_/A vssd1 vssd1 vccd1 vccd1 _13133_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18990_ _16876_/X _23192_/Q _18990_/S vssd1 vssd1 vccd1 vccd1 _18991_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_314_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_340_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17941_ _22825_/Q _17932_/X _17940_/X _17930_/X vssd1 vssd1 vccd1 vccd1 _22825_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_301_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13064_ _13064_/A _13064_/B vssd1 vssd1 vccd1 vccd1 _13064_/Y sky130_fd_sc_hd__nor2_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_305_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12015_ _23475_/Q _23571_/Q _22535_/Q _22339_/Q _12013_/X _12710_/A vssd1 vssd1 vccd1
+ vccd1 _12015_/X sky130_fd_sc_hd__mux4_1
X_17872_ _22807_/Q _17642_/X _17874_/S vssd1 vssd1 vccd1 vccd1 _17873_/A sky130_fd_sc_hd__mux2_1
XFILLER_266_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_294_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19611_ _19611_/A vssd1 vssd1 vccd1 vccd1 _23453_/D sky130_fd_sc_hd__clkbuf_1
X_16823_ _16822_/X _22523_/Q _16829_/S vssd1 vssd1 vccd1 vccd1 _16824_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19542_ _19542_/A vssd1 vssd1 vccd1 vccd1 _23422_/D sky130_fd_sc_hd__clkbuf_1
X_13966_ _13966_/A _13974_/B vssd1 vssd1 vccd1 vccd1 _13966_/Y sky130_fd_sc_hd__nor2_1
X_16754_ _16754_/A vssd1 vssd1 vccd1 vccd1 _22503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_321_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12917_ _13492_/B vssd1 vssd1 vccd1 vccd1 _13605_/A sky130_fd_sc_hd__clkinv_2
X_15705_ _15479_/A _13629_/Y _14529_/A vssd1 vssd1 vccd1 vccd1 _15705_/X sky130_fd_sc_hd__a21o_1
XFILLER_326_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19473_ _23392_/Q _18859_/X _19477_/S vssd1 vssd1 vccd1 vccd1 _19474_/A sky130_fd_sc_hd__mux2_1
X_16685_ _16779_/A vssd1 vssd1 vccd1 vccd1 _16704_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_321_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13897_ _13897_/A _13897_/B vssd1 vssd1 vccd1 vccd1 _14757_/A sky130_fd_sc_hd__xnor2_4
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_321_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18424_ _18427_/A _18427_/C _18423_/X vssd1 vssd1 vccd1 vccd1 _18424_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_221_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12848_ _23484_/Q _23580_/Q _22544_/Q _22348_/Q _12843_/X _12844_/X vssd1 vssd1 vccd1
+ vccd1 _12849_/B sky130_fd_sc_hd__mux4_1
XFILLER_221_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15636_ _15636_/A vssd1 vssd1 vccd1 vccd1 _15636_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18355_ _16168_/A _18357_/C _18354_/Y vssd1 vssd1 vccd1 vccd1 _22945_/D sky130_fd_sc_hd__o21a_1
X_15567_ _17149_/A _15375_/X _15564_/Y _15566_/X _15746_/A vssd1 vssd1 vccd1 vccd1
+ _15567_/X sky130_fd_sc_hd__a221o_1
X_12779_ _12784_/A _12779_/B vssd1 vssd1 vccd1 vccd1 _12779_/Y sky130_fd_sc_hd__nor2_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ _14518_/A vssd1 vssd1 vccd1 vccd1 _14518_/X sky130_fd_sc_hd__clkbuf_4
X_17306_ _22216_/A vssd1 vssd1 vccd1 vccd1 _22217_/A sky130_fd_sc_hd__buf_8
XFILLER_230_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18286_ _18286_/A _22922_/Q _18286_/C vssd1 vssd1 vccd1 vccd1 _18287_/C sky130_fd_sc_hd__and3_1
X_15498_ _16057_/A _15489_/X _15494_/Y _15497_/Y vssd1 vssd1 vccd1 vccd1 _15498_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_308_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14449_ _15589_/A vssd1 vssd1 vccd1 vccd1 _14450_/A sky130_fd_sc_hd__buf_2
X_17237_ _17237_/A vssd1 vssd1 vccd1 vccd1 _17237_/X sky130_fd_sc_hd__buf_2
XFILLER_175_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17168_ input86/X input51/X _17200_/S vssd1 vssd1 vccd1 vccd1 _17168_/X sky130_fd_sc_hd__mux2_8
XFILLER_174_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_344_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16119_ _21076_/A _15617_/X _15618_/X vssd1 vssd1 vccd1 vccd1 _16119_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_289_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17099_ _17073_/X _17098_/X _16968_/X _17078_/X vssd1 vssd1 vccd1 vccd1 _17099_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_305_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_288_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_332_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_331_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_331_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_296_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19809_ _23541_/Q _19217_/A _19815_/S vssd1 vssd1 vccd1 vccd1 _19810_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22820_ _23551_/CLK _22820_/D vssd1 vssd1 vccd1 vccd1 _22820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22751_ _23369_/CLK _22751_/D vssd1 vssd1 vccd1 vccd1 _22751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21702_ _23825_/Q _23759_/Q vssd1 vssd1 vccd1 vccd1 _21703_/B sky130_fd_sc_hd__nor2_1
XFILLER_225_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22682_ _23561_/CLK _22682_/D vssd1 vssd1 vccd1 vccd1 _22682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_358_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21633_ _23823_/Q _21632_/Y _21973_/S vssd1 vssd1 vccd1 vccd1 _21633_/X sky130_fd_sc_hd__mux2_4
XFILLER_240_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21564_ _21564_/A _21563_/Y vssd1 vssd1 vccd1 vccd1 _21566_/A sky130_fd_sc_hd__or2b_2
XFILLER_138_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_355_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_354_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23303_ _23527_/CLK _23303_/D vssd1 vssd1 vccd1 vccd1 _23303_/Q sky130_fd_sc_hd__dfxtp_1
X_20515_ _20515_/A _20515_/B _20515_/C _20515_/D vssd1 vssd1 vccd1 vccd1 _20526_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_138_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_327_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21495_ _21460_/A _21462_/B _21459_/Y vssd1 vssd1 vccd1 vccd1 _21496_/B sky130_fd_sc_hd__o21ai_1
XFILLER_193_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_179_wb_clk_i _23931_/CLK vssd1 vssd1 vccd1 vccd1 _23935_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_308_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23234_ _23554_/CLK _23234_/D vssd1 vssd1 vccd1 vccd1 _23234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20446_ _23697_/Q _20413_/X _20444_/Y _20445_/X vssd1 vssd1 vccd1 vccd1 _23697_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_108_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23551_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_326_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_307_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23165_ _23549_/CLK _23165_/D vssd1 vssd1 vccd1 vccd1 _23165_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_7115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20377_ _22139_/B vssd1 vssd1 vccd1 vccd1 _22140_/B sky130_fd_sc_hd__inv_2
XFILLER_106_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_7137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_7148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22116_ _22116_/A _22116_/B vssd1 vssd1 vccd1 vccd1 _22116_/Y sky130_fd_sc_hd__nand2_1
XTAP_7159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23096_ _23420_/CLK _23096_/D vssd1 vssd1 vccd1 vccd1 _23096_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_6425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22047_ _20353_/A _22045_/X _15926_/X _22046_/X vssd1 vssd1 vccd1 vccd1 _22047_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_6469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_342_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13820_ _12989_/B _13808_/A _13781_/A vssd1 vssd1 vccd1 vccd1 _13820_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_291_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_291_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13751_ _15113_/A vssd1 vssd1 vccd1 vccd1 _13874_/A sky130_fd_sc_hd__clkbuf_2
X_22949_ _23602_/CLK _22949_/D vssd1 vssd1 vccd1 vccd1 _22949_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_109 _13521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12702_ _12691_/Y _12694_/Y _12697_/Y _12701_/Y _11559_/X vssd1 vssd1 vccd1 vccd1
+ _12702_/X sky130_fd_sc_hd__o221a_1
XFILLER_204_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16470_ _16470_/A vssd1 vssd1 vccd1 vccd1 _22393_/D sky130_fd_sc_hd__clkbuf_1
X_13682_ _15901_/A vssd1 vssd1 vccd1 vccd1 _14833_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_325_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15421_ _18811_/A vssd1 vssd1 vccd1 vccd1 _19204_/A sky130_fd_sc_hd__clkbuf_2
X_12633_ _12626_/Y _12628_/Y _12630_/Y _12632_/Y _11657_/X vssd1 vssd1 vccd1 vccd1
+ _12634_/C sky130_fd_sc_hd__o221a_2
XPHY_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_346_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18140_ _22892_/Q vssd1 vssd1 vccd1 vccd1 _18163_/A sky130_fd_sc_hd__clkbuf_2
X_15352_ _23600_/Q _14901_/X _14902_/X _23632_/Q vssd1 vssd1 vccd1 vccd1 _15352_/X
+ sky130_fd_sc_hd__o22a_2
XPHY_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12564_ _23465_/Q _23561_/Q _22525_/Q _22329_/Q _12245_/S _12292_/X vssd1 vssd1 vccd1
+ vccd1 _12565_/B sky130_fd_sc_hd__mux4_1
XFILLER_357_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14303_ _14299_/X _14302_/X _14639_/A vssd1 vssd1 vccd1 vccd1 _14303_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11515_ _11515_/A vssd1 vssd1 vccd1 vccd1 _13216_/A sky130_fd_sc_hd__clkbuf_2
X_18071_ _22861_/Q _18066_/X _18070_/X _18060_/X vssd1 vssd1 vccd1 vccd1 _22861_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15283_ _19194_/A vssd1 vssd1 vccd1 vccd1 _15283_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12495_ _12596_/B _12493_/X _12494_/X vssd1 vssd1 vccd1 vccd1 _13506_/B sky130_fd_sc_hd__o21a_2
X_17022_ _17022_/A _17022_/B vssd1 vssd1 vccd1 vccd1 _17047_/A sky130_fd_sc_hd__and2_1
XFILLER_138_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14234_ _14234_/A _15119_/A vssd1 vssd1 vccd1 vccd1 _14235_/A sky130_fd_sc_hd__or2b_4
XFILLER_144_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_345_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11446_ _11502_/A _11446_/B vssd1 vssd1 vccd1 vccd1 _11446_/X sky130_fd_sc_hd__or2_1
XFILLER_138_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_291_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14165_ _22909_/Q _14394_/A _14164_/X _22602_/Q vssd1 vssd1 vccd1 vccd1 _14552_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_314_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_298_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11377_ _11657_/A vssd1 vssd1 vccd1 vccd1 _11378_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_4_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_291_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13116_ _22287_/Q _23103_/Q _23519_/Q _22448_/Q _13114_/X _13115_/X vssd1 vssd1 vccd1
+ vccd1 _13117_/B sky130_fd_sc_hd__mux4_2
XFILLER_316_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18973_ _16851_/X _23184_/Q _18979_/S vssd1 vssd1 vccd1 vccd1 _18974_/A sky130_fd_sc_hd__mux2_1
X_14096_ _22595_/Q _14081_/A _14095_/Y _14012_/X vssd1 vssd1 vccd1 vccd1 _14096_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_301_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_316_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17924_ _22820_/Q _17914_/X _17923_/X _17912_/X vssd1 vssd1 vccd1 vccd1 _22820_/D
+ sky130_fd_sc_hd__o211a_1
X_13047_ _13191_/S vssd1 vssd1 vccd1 vccd1 _13088_/S sky130_fd_sc_hd__buf_4
XFILLER_79_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17855_ _22799_/Q _17617_/X _17859_/S vssd1 vssd1 vccd1 vccd1 _17856_/A sky130_fd_sc_hd__mux2_1
XFILLER_266_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16806_ input9/X _16806_/B vssd1 vssd1 vccd1 vccd1 _16808_/C sky130_fd_sc_hd__or2_1
XFILLER_293_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17786_ _17786_/A vssd1 vssd1 vccd1 vccd1 _22768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_282_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14998_ _15346_/A _14991_/X _14997_/X _14748_/X vssd1 vssd1 vccd1 vccd1 _14998_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_226_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19525_ _19223_/X _23415_/Q _19527_/S vssd1 vssd1 vccd1 vccd1 _19526_/A sky130_fd_sc_hd__mux2_1
X_16737_ _22499_/Q _16729_/X _16730_/X input13/X vssd1 vssd1 vccd1 vccd1 _16738_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_241_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13949_ _23921_/Q vssd1 vssd1 vccd1 vccd1 _21636_/A sky130_fd_sc_hd__buf_2
XFILLER_46_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19456_ _19456_/A vssd1 vssd1 vccd1 vccd1 _23384_/D sky130_fd_sc_hd__clkbuf_1
X_16668_ _16668_/A vssd1 vssd1 vccd1 vccd1 _22480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18407_ _19932_/A vssd1 vssd1 vccd1 vccd1 _19923_/A sky130_fd_sc_hd__buf_6
XFILLER_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15619_ _17159_/A _15617_/X _15618_/X vssd1 vssd1 vccd1 vccd1 _15619_/Y sky130_fd_sc_hd__o21ai_2
X_19387_ _19387_/A vssd1 vssd1 vccd1 vccd1 _23353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_349_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16599_ _16089_/X _22450_/Q _16601_/S vssd1 vssd1 vccd1 vccd1 _16600_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18338_ _15950_/X _18341_/C _18337_/X vssd1 vssd1 vccd1 vccd1 _18338_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_188_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_6_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23369_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_337_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18269_ _22917_/Q _18264_/C _18268_/Y vssd1 vssd1 vccd1 vccd1 _22917_/D sky130_fd_sc_hd__o21a_1
XFILLER_175_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20300_ _23669_/Q _20338_/B vssd1 vssd1 vccd1 vccd1 _20300_/X sky130_fd_sc_hd__or2_1
XFILLER_357_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21280_ _21280_/A _21283_/B vssd1 vssd1 vccd1 vccd1 _21280_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_201_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23048_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20231_ _20226_/X _21515_/A _20230_/X vssd1 vssd1 vccd1 vccd1 _21013_/A sky130_fd_sc_hd__a21oi_4
XFILLER_289_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_304_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20162_ _20344_/A vssd1 vssd1 vccd1 vccd1 _20379_/A sky130_fd_sc_hd__buf_2
XFILLER_320_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_320_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20093_ _20121_/A vssd1 vssd1 vccd1 vccd1 _20120_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23921_ _23926_/CLK _23921_/D vssd1 vssd1 vccd1 vccd1 _23921_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23852_ _23856_/CLK _23852_/D vssd1 vssd1 vccd1 vccd1 _23852_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22803_ _23583_/CLK _22803_/D vssd1 vssd1 vccd1 vccd1 _22803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_309_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23783_ _23911_/CLK _23783_/D vssd1 vssd1 vccd1 vccd1 _23783_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20995_ _21072_/B vssd1 vssd1 vccd1 vccd1 _20996_/B sky130_fd_sc_hd__buf_4
XFILLER_25_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22734_ _23068_/CLK _22734_/D vssd1 vssd1 vccd1 vccd1 _22734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22665_ _23571_/CLK _22665_/D vssd1 vssd1 vccd1 vccd1 _22665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_336_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_328_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21616_ _21616_/A _21870_/A vssd1 vssd1 vccd1 vccd1 _21616_/Y sky130_fd_sc_hd__nand2_1
XFILLER_139_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22596_ _22974_/CLK _22596_/D vssd1 vssd1 vccd1 vccd1 _22596_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_138_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21547_ _21428_/B _21542_/X _21543_/X _21545_/X _21546_/X vssd1 vssd1 vccd1 vccd1
+ _21548_/B sky130_fd_sc_hd__a311o_4
XFILLER_194_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11300_ _11343_/A vssd1 vssd1 vccd1 vccd1 _13278_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_342_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12280_ _12401_/A _12279_/X _11680_/A vssd1 vssd1 vccd1 vccd1 _12280_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_107_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21478_ _13910_/X _21305_/X _21477_/X _21281_/X vssd1 vssd1 vccd1 vccd1 _23916_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11231_ _11965_/A vssd1 vssd1 vccd1 vccd1 _11232_/A sky130_fd_sc_hd__buf_2
X_23217_ _23507_/CLK _23217_/D vssd1 vssd1 vccd1 vccd1 _23217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20429_ _23691_/Q _20429_/B vssd1 vssd1 vccd1 vccd1 _20429_/X sky130_fd_sc_hd__or2_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_311_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23148_ _23950_/A _23148_/D vssd1 vssd1 vccd1 vccd1 _23148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11162_ _12246_/A vssd1 vssd1 vccd1 vccd1 _11163_/A sky130_fd_sc_hd__buf_4
XFILLER_323_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_296_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_296_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15970_ _21078_/B _15617_/X _15618_/X vssd1 vssd1 vccd1 vccd1 _15970_/Y sky130_fd_sc_hd__o21ai_1
X_11093_ _23885_/Q _23884_/Q _23883_/Q vssd1 vssd1 vccd1 vccd1 _11095_/C sky130_fd_sc_hd__or3_1
X_23079_ _23555_/CLK _23079_/D vssd1 vssd1 vccd1 vccd1 _23079_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14921_ _23753_/Q _14911_/X _14913_/X _14915_/X _14920_/X vssd1 vssd1 vccd1 vccd1
+ _14921_/X sky130_fd_sc_hd__a221o_1
XTAP_6299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_76_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23549_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17640_ _22707_/Q _17639_/X _17640_/S vssd1 vssd1 vccd1 vccd1 _17641_/A sky130_fd_sc_hd__mux2_1
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14852_ _14850_/X _14851_/X _14852_/S vssd1 vssd1 vccd1 vccd1 _14852_/X sky130_fd_sc_hd__mux2_2
XFILLER_91_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13803_ _13803_/A _13875_/B vssd1 vssd1 vccd1 vccd1 _13852_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17571_ _17571_/A vssd1 vssd1 vccd1 vccd1 _22685_/D sky130_fd_sc_hd__clkbuf_1
X_14783_ _14781_/X _14782_/X _14852_/S vssd1 vssd1 vccd1 vccd1 _14784_/A sky130_fd_sc_hd__mux2_2
X_11995_ _12900_/A _11994_/X _11631_/A vssd1 vssd1 vccd1 vccd1 _11995_/X sky130_fd_sc_hd__o21a_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19310_ _19310_/A vssd1 vssd1 vccd1 vccd1 _23319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16522_ _16089_/X _22417_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _16523_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13734_ _13745_/B vssd1 vssd1 vccd1 vccd1 _13771_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_44_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_323_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19241_ _19241_/A vssd1 vssd1 vccd1 vccd1 _23292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13665_ _13665_/A _13670_/A _13670_/B _13670_/C vssd1 vssd1 vccd1 vccd1 _14002_/A
+ sky130_fd_sc_hd__or4_4
X_16453_ _16161_/X _22387_/Q _16455_/S vssd1 vssd1 vccd1 vccd1 _16454_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12616_ _12708_/A _12616_/B vssd1 vssd1 vccd1 vccd1 _12616_/Y sky130_fd_sc_hd__nor2_1
X_15404_ _14745_/A _15397_/X _15403_/Y _15652_/A vssd1 vssd1 vccd1 vccd1 _15405_/B
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16384_ _18770_/A _19090_/A _19090_/B vssd1 vssd1 vccd1 vccd1 _18625_/B sky130_fd_sc_hd__or3b_4
X_19172_ _19172_/A vssd1 vssd1 vccd1 vccd1 _19172_/X sky130_fd_sc_hd__clkbuf_2
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13596_ _13619_/A _13531_/X _12005_/Y _13611_/A vssd1 vssd1 vccd1 vccd1 _13612_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_346_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18123_ _22886_/Q _22878_/Q _18126_/S vssd1 vssd1 vccd1 vccd1 _18123_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15335_ _15335_/A _15335_/B vssd1 vssd1 vccd1 vccd1 _15335_/Y sky130_fd_sc_hd__nor2_1
X_12547_ _14292_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _12547_/X sky130_fd_sc_hd__and2b_1
XFILLER_145_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_346_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18054_ _18054_/A vssd1 vssd1 vccd1 vccd1 _18054_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15266_ _21630_/A _15211_/X _15262_/X _15265_/X _14612_/X vssd1 vssd1 vccd1 vccd1
+ _15266_/X sky130_fd_sc_hd__a221o_2
X_12478_ _12489_/A _12477_/X _11818_/A vssd1 vssd1 vccd1 vccd1 _12478_/X sky130_fd_sc_hd__o21a_1
XFILLER_333_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_327_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17005_ _20508_/B _16978_/Y _16932_/A _16947_/X vssd1 vssd1 vccd1 vccd1 _17005_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_172_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14217_ _15109_/A vssd1 vssd1 vccd1 vccd1 _14725_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11429_ _13095_/A vssd1 vssd1 vccd1 vccd1 _11497_/A sky130_fd_sc_hd__buf_4
XFILLER_160_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15197_ _13942_/A _15196_/X _14761_/A vssd1 vssd1 vccd1 vccd1 _15198_/B sky130_fd_sc_hd__a21oi_1
XFILLER_302_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_299_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14148_ _14148_/A _14148_/B _14148_/C _13662_/B vssd1 vssd1 vccd1 vccd1 _16966_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_141_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_342_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14079_ _14083_/A _14724_/A _14009_/X _22812_/Q vssd1 vssd1 vccd1 vccd1 _14079_/X
+ sky130_fd_sc_hd__a22o_4
X_18956_ _18956_/A vssd1 vssd1 vccd1 vccd1 _23176_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17907_ _22815_/Q _17891_/X _17906_/X _17657_/X vssd1 vssd1 vccd1 vccd1 _22815_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_301_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18887_ _18944_/S vssd1 vssd1 vccd1 vccd1 _18896_/S sky130_fd_sc_hd__buf_4
XFILLER_239_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17838_ _17838_/A vssd1 vssd1 vccd1 vccd1 _22791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17769_ _17769_/A vssd1 vssd1 vccd1 vccd1 _22760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_270_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19508_ _19197_/X _23407_/Q _19516_/S vssd1 vssd1 vccd1 vccd1 _19509_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20780_ _23750_/Q _20786_/B _20779_/X _20763_/X vssd1 vssd1 vccd1 vccd1 _23750_/D
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_440 _23916_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_451 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19439_ _19439_/A vssd1 vssd1 vccd1 vccd1 _23376_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_462 _20723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_473 _21616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_484 _14224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_495 _14099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22450_ _23489_/CLK _22450_/D vssd1 vssd1 vccd1 vccd1 _22450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21401_ _21401_/A _21400_/Y vssd1 vssd1 vccd1 vccd1 _21404_/A sky130_fd_sc_hd__or2b_1
X_22381_ _23451_/CLK _22381_/D vssd1 vssd1 vccd1 vccd1 _22381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_325_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_324_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21332_ _21663_/A vssd1 vssd1 vccd1 vccd1 _21942_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_325_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_336_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21263_ _15674_/X _15830_/Y _21242_/A _20058_/X vssd1 vssd1 vccd1 vccd1 _21263_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23002_ _23592_/CLK _23002_/D vssd1 vssd1 vccd1 vccd1 _23002_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_305_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20214_ _20214_/A _20214_/B vssd1 vssd1 vccd1 vccd1 _20254_/A sky130_fd_sc_hd__nor2_1
XFILLER_351_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_333_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21194_ _21260_/S vssd1 vssd1 vccd1 vccd1 _21214_/S sky130_fd_sc_hd__buf_2
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_320_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20145_ _20333_/A vssd1 vssd1 vccd1 vccd1 _20213_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_277_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ _23632_/Q _20079_/B _20076_/C _20076_/D vssd1 vssd1 vccd1 vccd1 _20085_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_286_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23904_ _23910_/CLK _23904_/D vssd1 vssd1 vccd1 vccd1 _23904_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23835_ _23876_/CLK _23835_/D vssd1 vssd1 vccd1 vccd1 _23835_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23766_ _23768_/CLK _23766_/D vssd1 vssd1 vccd1 vccd1 _23766_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11780_ _11780_/A vssd1 vssd1 vccd1 vccd1 _11780_/X sky130_fd_sc_hd__buf_4
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20978_ _21023_/A vssd1 vssd1 vccd1 vccd1 _20978_/X sky130_fd_sc_hd__buf_4
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22717_ _23054_/CLK _22717_/D vssd1 vssd1 vccd1 vccd1 _22717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23697_ _23704_/CLK _23697_/D vssd1 vssd1 vccd1 vccd1 _23697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_194_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23526_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_41_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13450_ _13473_/B vssd1 vssd1 vccd1 vccd1 _13451_/A sky130_fd_sc_hd__buf_2
XFILLER_347_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22648_ _23054_/CLK _22648_/D vssd1 vssd1 vccd1 vccd1 _22648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_327_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_123_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23643_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_278_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12401_ _12401_/A _12401_/B vssd1 vssd1 vccd1 vccd1 _12401_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13381_ _13382_/B _13382_/C _13948_/A vssd1 vssd1 vccd1 vccd1 _13392_/B sky130_fd_sc_hd__a21oi_1
X_22579_ _23643_/CLK _22579_/D vssd1 vssd1 vccd1 vccd1 _22579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15120_ _13879_/A _15116_/Y _15532_/A _13834_/A vssd1 vssd1 vccd1 vccd1 _15120_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_154_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12332_ _23306_/Q _23274_/Q _23242_/Q _23530_/Q _12314_/X _12325_/X vssd1 vssd1 vccd1
+ vccd1 _12332_/X sky130_fd_sc_hd__mux4_2
XFILLER_194_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15051_ _15159_/B _15051_/B vssd1 vssd1 vccd1 vccd1 _15051_/Y sky130_fd_sc_hd__nor2_1
X_12263_ _23307_/Q _23275_/Q _23243_/Q _23531_/Q _11455_/A _11733_/A vssd1 vssd1 vccd1
+ vccd1 _12264_/B sky130_fd_sc_hd__mux4_1
XFILLER_107_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_324_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14002_ _14002_/A _14072_/C vssd1 vssd1 vccd1 vccd1 _14041_/A sky130_fd_sc_hd__nor2_2
XFILLER_324_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11214_ _11214_/A vssd1 vssd1 vccd1 vccd1 _11215_/A sky130_fd_sc_hd__buf_6
XFILLER_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12194_ _23404_/Q _23020_/Q _23372_/Q _23340_/Q _12242_/S _11611_/A vssd1 vssd1 vccd1
+ vccd1 _12194_/X sky130_fd_sc_hd__mux4_2
XFILLER_269_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18810_ _18810_/A vssd1 vssd1 vccd1 vccd1 _23120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11145_ _13041_/A vssd1 vssd1 vccd1 vccd1 _13259_/A sky130_fd_sc_hd__buf_2
XFILLER_123_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_311_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19790_ _19790_/A vssd1 vssd1 vccd1 vccd1 _23532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18741_ _16876_/X _23096_/Q _18741_/S vssd1 vssd1 vccd1 vccd1 _18742_/A sky130_fd_sc_hd__mux2_1
XTAP_6074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15953_ _23614_/Q _15589_/X _15590_/X _23646_/Q vssd1 vssd1 vccd1 vccd1 _15953_/X
+ sky130_fd_sc_hd__o22a_2
XTAP_6085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11076_ _23885_/Q vssd1 vssd1 vccd1 vccd1 _14132_/A sky130_fd_sc_hd__clkbuf_2
XTAP_6096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput140 dout1[3] vssd1 vssd1 vccd1 vccd1 input140/X sky130_fd_sc_hd__clkbuf_1
XFILLER_209_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_313_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput151 dout1[4] vssd1 vssd1 vccd1 vccd1 input151/X sky130_fd_sc_hd__clkbuf_1
Xinput162 dout1[5] vssd1 vssd1 vccd1 vccd1 input162/X sky130_fd_sc_hd__clkbuf_1
XTAP_5373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14904_ _15592_/A vssd1 vssd1 vccd1 vccd1 _14905_/A sky130_fd_sc_hd__buf_2
XTAP_5384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18672_ _23065_/Q _17610_/X _18680_/S vssd1 vssd1 vccd1 vccd1 _18673_/A sky130_fd_sc_hd__mux2_1
Xinput173 irq[11] vssd1 vssd1 vccd1 vccd1 _20521_/C sky130_fd_sc_hd__buf_2
X_15884_ _14730_/X _15877_/X _15883_/Y _15150_/X vssd1 vssd1 vccd1 vccd1 _15885_/B
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_5395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput184 irq[7] vssd1 vssd1 vccd1 vccd1 _20514_/C sky130_fd_sc_hd__buf_2
XFILLER_49_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput195 localMemory_wb_adr_i[14] vssd1 vssd1 vccd1 vccd1 input195/X sky130_fd_sc_hd__clkbuf_1
XFILLER_264_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17623_ _18849_/A vssd1 vssd1 vccd1 vccd1 _17623_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_236_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ _14835_/A vssd1 vssd1 vccd1 vccd1 _20186_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_252_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _22680_/Q _17553_/X _17560_/S vssd1 vssd1 vccd1 vccd1 _17555_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11978_ _11969_/Y _11971_/Y _11975_/Y _11977_/Y _11244_/A vssd1 vssd1 vccd1 vccd1
+ _11978_/X sky130_fd_sc_hd__o221a_1
XFILLER_205_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14766_ _14854_/S _14648_/X _14376_/X vssd1 vssd1 vccd1 vccd1 _14766_/X sky130_fd_sc_hd__o21a_1
XFILLER_45_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16505_ _15785_/X _22409_/Q _16513_/S vssd1 vssd1 vccd1 vccd1 _16506_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13717_ _14072_/B vssd1 vssd1 vccd1 vccd1 _14015_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_260_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14697_ _16191_/A vssd1 vssd1 vccd1 vccd1 _15162_/A sky130_fd_sc_hd__clkbuf_2
X_17485_ _17542_/S vssd1 vssd1 vccd1 vccd1 _17494_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_177_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19224_ _19223_/X _23287_/Q _19227_/S vssd1 vssd1 vccd1 vccd1 _19225_/A sky130_fd_sc_hd__mux2_1
XFILLER_338_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16436_ _15861_/X _22379_/Q _16440_/S vssd1 vssd1 vccd1 vccd1 _16437_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13648_ _21293_/A _21673_/A _13490_/X _13647_/Y vssd1 vssd1 vccd1 vccd1 _13652_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_319_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _23265_/Q _18862_/X _19157_/S vssd1 vssd1 vccd1 vccd1 _19156_/A sky130_fd_sc_hd__mux2_1
X_16367_ _16367_/A vssd1 vssd1 vccd1 vccd1 _22349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13579_ _13579_/A _13579_/B vssd1 vssd1 vccd1 vccd1 _13580_/B sky130_fd_sc_hd__or2_1
XFILLER_158_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_347_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_318_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18106_ _22873_/Q _18096_/X _18104_/X _18105_/X vssd1 vssd1 vccd1 vccd1 _22873_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_346_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15318_ _15318_/A _15318_/B vssd1 vssd1 vccd1 vccd1 _15318_/Y sky130_fd_sc_hd__nor2_1
XFILLER_318_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16298_ _22321_/Q _16297_/X _16301_/S vssd1 vssd1 vccd1 vccd1 _16299_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19086_ _16911_/X _23235_/Q _19088_/S vssd1 vssd1 vccd1 vccd1 _19087_/A sky130_fd_sc_hd__mux2_1
XFILLER_338_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_318_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_334_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_5_1_wb_clk_i clkbuf_3_5_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_1_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_274_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18037_ _18053_/A vssd1 vssd1 vccd1 vccd1 _18037_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_219_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15249_ _14659_/X _14642_/X _15249_/S vssd1 vssd1 vccd1 vccd1 _15250_/A sky130_fd_sc_hd__mux2_1
XFILLER_321_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_299_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_302_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_342_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19988_ _23609_/Q _23608_/Q _19988_/C vssd1 vssd1 vccd1 vccd1 _19994_/C sky130_fd_sc_hd__and3_1
XFILLER_287_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_302_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_286_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18939_ _18939_/A vssd1 vssd1 vccd1 vccd1 _23169_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_268_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21950_ _21950_/A _21954_/A vssd1 vssd1 vccd1 vccd1 _21951_/B sky130_fd_sc_hd__or2_1
XFILLER_55_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20901_ _23782_/Q _20893_/X _20900_/X _20788_/X vssd1 vssd1 vccd1 vccd1 _23782_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21881_ _21837_/A _21837_/B _21836_/A vssd1 vssd1 vccd1 vccd1 _21885_/A sky130_fd_sc_hd__a21oi_1
XFILLER_254_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23620_ _23624_/CLK _23620_/D vssd1 vssd1 vccd1 vccd1 _23620_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_270_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20832_ _20832_/A vssd1 vssd1 vccd1 vccd1 _23763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_299_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23551_ _23551_/CLK _23551_/D vssd1 vssd1 vccd1 vccd1 _23551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20763_ _20763_/A vssd1 vssd1 vccd1 vccd1 _20763_/X sky130_fd_sc_hd__buf_2
XFILLER_251_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_270 _18827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_357_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_281 _15883_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22502_ _23684_/CLK _22502_/D vssd1 vssd1 vccd1 vccd1 _22502_/Q sky130_fd_sc_hd__dfxtp_4
XINSDIODE2_292 _18852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23482_ _23546_/CLK _23482_/D vssd1 vssd1 vccd1 vccd1 _23482_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_210_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20694_ _21899_/A _20648_/X _20693_/Y vssd1 vssd1 vccd1 vccd1 _20695_/C sky130_fd_sc_hd__a21oi_2
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22433_ _23504_/CLK _22433_/D vssd1 vssd1 vccd1 vccd1 _22433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_309_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_353_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22364_ _23500_/CLK _22364_/D vssd1 vssd1 vccd1 vccd1 _22364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21315_ _17655_/A _23911_/Q vssd1 vssd1 vccd1 vccd1 _21319_/A sky130_fd_sc_hd__nand2b_1
X_22295_ _22779_/CLK _22295_/D vssd1 vssd1 vccd1 vccd1 _22295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_312_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_306_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21246_ _17159_/A _15579_/X _21257_/S vssd1 vssd1 vccd1 vccd1 _21247_/B sky130_fd_sc_hd__mux2_1
XFILLER_305_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_334_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_321_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21177_ _21177_/A _21177_/B vssd1 vssd1 vccd1 vccd1 _21177_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20128_ _23649_/Q _20127_/C _20101_/X vssd1 vssd1 vccd1 vccd1 _20128_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_277_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12950_ _13006_/A _12947_/X _12949_/X _12721_/X vssd1 vssd1 vccd1 vccd1 _12950_/X
+ sky130_fd_sc_hd__o211a_1
X_20059_ _23629_/Q _20066_/A _20066_/B _20066_/C _20058_/X vssd1 vssd1 vccd1 vccd1
+ _20059_/X sky130_fd_sc_hd__a41o_1
XFILLER_18_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11901_ _11905_/A _11901_/B vssd1 vssd1 vccd1 vccd1 _11901_/Y sky130_fd_sc_hd__nor2_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _23322_/Q _23290_/Q _23258_/Q _23546_/Q _12755_/X _11594_/A vssd1 vssd1 vccd1
+ vccd1 _12882_/B sky130_fd_sc_hd__mux4_1
XFILLER_218_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14620_ _14762_/A vssd1 vssd1 vccd1 vccd1 _14621_/A sky130_fd_sc_hd__clkbuf_2
X_11832_ _11853_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11832_/Y sky130_fd_sc_hd__nor2_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23818_ _23818_/CLK _23818_/D vssd1 vssd1 vccd1 vccd1 _23818_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14551_ _14551_/A _14551_/B _14551_/C vssd1 vssd1 vccd1 vccd1 _16935_/B sky130_fd_sc_hd__or3_1
XFILLER_214_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23749_ _23911_/CLK _23749_/D vssd1 vssd1 vccd1 vccd1 _23749_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _21652_/A _11763_/B vssd1 vssd1 vccd1 vccd1 _11763_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _13502_/A vssd1 vssd1 vccd1 vccd1 _13508_/B sky130_fd_sc_hd__inv_2
X_17270_ _23487_/Q _17230_/X _17231_/X _17268_/X _17269_/Y vssd1 vssd1 vccd1 vccd1
+ _17270_/X sky130_fd_sc_hd__a32o_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _15215_/A vssd1 vssd1 vccd1 vccd1 _14482_/X sky130_fd_sc_hd__buf_2
XFILLER_13_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11694_ _12196_/A vssd1 vssd1 vccd1 vccd1 _12241_/A sky130_fd_sc_hd__buf_4
XFILLER_201_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13433_ _13433_/A vssd1 vssd1 vccd1 vccd1 _13433_/X sky130_fd_sc_hd__clkbuf_1
X_16221_ _22297_/Q _16220_/X _16221_/S vssd1 vssd1 vccd1 vccd1 _16222_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_328_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_329_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16152_ _22219_/A _16151_/C _22216_/A vssd1 vssd1 vccd1 vccd1 _16153_/B sky130_fd_sc_hd__a21oi_1
XFILLER_356_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13364_ _13364_/A _14294_/A vssd1 vssd1 vccd1 vccd1 _13364_/X sky130_fd_sc_hd__or2_1
XFILLER_177_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_355_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_343_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12315_ _22362_/Q _22394_/Q _22683_/Q _23050_/Q _12314_/X _11815_/X vssd1 vssd1 vccd1
+ vccd1 _12316_/B sky130_fd_sc_hd__mux4_2
XFILLER_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15103_ _18792_/A vssd1 vssd1 vccd1 vccd1 _19185_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_315_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16083_ _16080_/X _16081_/X _21605_/A _15375_/X vssd1 vssd1 vccd1 vccd1 _16083_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_304_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13295_ _13295_/A _13295_/B _13295_/C vssd1 vssd1 vccd1 vccd1 _20381_/A sky130_fd_sc_hd__nor3_4
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_308_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_315_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ _22492_/Q _14232_/X _14247_/X _15033_/X _14071_/A vssd1 vssd1 vccd1 vccd1
+ _15034_/X sky130_fd_sc_hd__o221a_1
X_19911_ _16303_/X _23587_/Q _19913_/S vssd1 vssd1 vccd1 vccd1 _19912_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12246_ _12246_/A _12246_/B vssd1 vssd1 vccd1 vccd1 _12246_/Y sky130_fd_sc_hd__nand2_1
XFILLER_308_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_91_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23880_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_296_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_296_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19842_ _19842_/A vssd1 vssd1 vccd1 vccd1 _23556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12177_ _23899_/Q vssd1 vssd1 vccd1 vccd1 _12537_/S sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_20_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _22779_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_311_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_324_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ _11780_/A vssd1 vssd1 vccd1 vccd1 _11713_/A sky130_fd_sc_hd__buf_4
XFILLER_288_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19773_ _19841_/S vssd1 vssd1 vccd1 vccd1 _19782_/S sky130_fd_sc_hd__clkbuf_8
X_16985_ _17224_/B vssd1 vssd1 vccd1 vccd1 _17033_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_324_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18724_ _16851_/X _23088_/Q _18730_/S vssd1 vssd1 vccd1 vccd1 _18725_/A sky130_fd_sc_hd__mux2_1
X_15936_ _19242_/A vssd1 vssd1 vccd1 vccd1 _15936_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_265_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18655_ _18655_/A vssd1 vssd1 vccd1 vccd1 _23057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15867_ _13400_/C _13592_/Y _15867_/S vssd1 vssd1 vccd1 vccd1 _15867_/X sky130_fd_sc_hd__mux2_1
XFILLER_329_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17606_ _17606_/A vssd1 vssd1 vccd1 vccd1 _22696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_252_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14818_ _16079_/A vssd1 vssd1 vccd1 vccd1 _15318_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_340_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18586_ _16860_/X _23027_/Q _18586_/S vssd1 vssd1 vccd1 vccd1 _18587_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15798_ _15798_/A _15798_/B vssd1 vssd1 vccd1 vccd1 _15798_/Y sky130_fd_sc_hd__nor2_2
X_17537_ _17537_/A vssd1 vssd1 vccd1 vccd1 _22674_/D sky130_fd_sc_hd__clkbuf_1
X_14749_ _14730_/X _14735_/X _14747_/X _14748_/X vssd1 vssd1 vccd1 vccd1 _14749_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_339_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17468_ _17468_/A vssd1 vssd1 vccd1 vccd1 _22644_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19207_ _19207_/A vssd1 vssd1 vccd1 vccd1 _19207_/X sky130_fd_sc_hd__clkbuf_2
X_16419_ _16419_/A vssd1 vssd1 vccd1 vccd1 _22371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_349_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17399_ _19555_/A _19164_/A vssd1 vssd1 vccd1 vccd1 _17456_/A sky130_fd_sc_hd__nor2_4
XFILLER_193_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19138_ _23257_/Q _18836_/X _19146_/S vssd1 vssd1 vccd1 vccd1 _19139_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_334_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19069_ _16886_/X _23227_/Q _19073_/S vssd1 vssd1 vccd1 vccd1 _19070_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput400 _14017_/X vssd1 vssd1 vccd1 vccd1 din0[4] sky130_fd_sc_hd__buf_2
XFILLER_322_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput411 _22565_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[12] sky130_fd_sc_hd__buf_2
X_21100_ _21108_/A _21100_/B vssd1 vssd1 vccd1 vccd1 _23847_/D sky130_fd_sc_hd__nor2_1
XFILLER_173_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput422 _22575_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[22] sky130_fd_sc_hd__buf_2
XFILLER_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_306_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput433 _22556_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[3] sky130_fd_sc_hd__buf_2
X_22080_ _23838_/Q _23772_/Q vssd1 vssd1 vccd1 vccd1 _22081_/B sky130_fd_sc_hd__nor2_1
XFILLER_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput444 _23944_/Q vssd1 vssd1 vccd1 vccd1 probe_errorCode[1] sky130_fd_sc_hd__buf_2
Xoutput455 _23880_/Q vssd1 vssd1 vccd1 vccd1 probe_opcode[1] sky130_fd_sc_hd__buf_2
XFILLER_271_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput466 _23925_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[14] sky130_fd_sc_hd__buf_2
X_21031_ _23827_/Q _21048_/B vssd1 vssd1 vccd1 vccd1 _21031_/X sky130_fd_sc_hd__or2_1
Xoutput477 _23935_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[24] sky130_fd_sc_hd__buf_2
Xoutput488 _23916_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[5] sky130_fd_sc_hd__buf_2
Xoutput499 _14076_/X vssd1 vssd1 vccd1 vccd1 wmask0[2] sky130_fd_sc_hd__buf_2
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_287_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22982_ _23424_/CLK _22982_/D vssd1 vssd1 vccd1 vccd1 _22982_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21933_ _21933_/A _21933_/B vssd1 vssd1 vccd1 vccd1 _21934_/C sky130_fd_sc_hd__nor2_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21864_ _21856_/A _21714_/A _21839_/X _21863_/Y _21681_/X vssd1 vssd1 vccd1 vccd1
+ _23928_/D sky130_fd_sc_hd__o221a_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23603_ _23651_/CLK _23603_/D vssd1 vssd1 vccd1 vccd1 _23603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20815_ _20635_/B _20810_/X _20811_/X _23759_/Q vssd1 vssd1 vccd1 vccd1 _20816_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21795_ _22061_/A _21788_/X _21794_/X _21408_/X vssd1 vssd1 vccd1 vccd1 _21795_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_24_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23534_ _23534_/CLK _23534_/D vssd1 vssd1 vccd1 vccd1 _23534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20746_ _22140_/A _20732_/X _20745_/Y vssd1 vssd1 vccd1 vccd1 _20747_/C sky130_fd_sc_hd__a21oi_4
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23465_ _23555_/CLK _23465_/D vssd1 vssd1 vccd1 vccd1 _23465_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_326_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20677_ _17163_/A _20632_/X _20676_/X vssd1 vssd1 vccd1 vccd1 _20678_/C sky130_fd_sc_hd__o21a_2
XFILLER_137_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22416_ _23584_/CLK _22416_/D vssd1 vssd1 vccd1 vccd1 _22416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_338_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23396_ _23578_/CLK _23396_/D vssd1 vssd1 vccd1 vccd1 _23396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_337_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22347_ _23515_/CLK _22347_/D vssd1 vssd1 vccd1 vccd1 _22347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12100_ _23218_/Q _23186_/Q _23154_/Q _23122_/Q _12094_/X _11755_/A vssd1 vssd1 vccd1
+ vccd1 _12101_/B sky130_fd_sc_hd__mux4_1
XFILLER_151_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_352_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13080_ _13080_/A vssd1 vssd1 vccd1 vccd1 _13082_/A sky130_fd_sc_hd__inv_2
X_22278_ _23510_/CLK _22278_/D vssd1 vssd1 vccd1 vccd1 _22278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12031_ _12708_/A _12030_/X _11631_/X vssd1 vssd1 vccd1 vccd1 _12031_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21229_ _21242_/A vssd1 vssd1 vccd1 vccd1 _21229_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_239_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_321_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_320_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_293_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16770_ _22508_/Q _16765_/X _16766_/X input23/X vssd1 vssd1 vccd1 vccd1 _16771_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_65_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13982_ _13982_/A vssd1 vssd1 vccd1 vccd1 _13982_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15721_ _13599_/A _14674_/A _15720_/X vssd1 vssd1 vccd1 vccd1 _15721_/Y sky130_fd_sc_hd__a21oi_2
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _12919_/A _12932_/X _11133_/A vssd1 vssd1 vccd1 vccd1 _12933_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_274_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18440_ _22974_/Q _22975_/Q _18440_/C vssd1 vssd1 vccd1 vccd1 _18444_/B sky130_fd_sc_hd__and3_1
XFILLER_234_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _15652_/A vssd1 vssd1 vccd1 vccd1 _15652_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12864_ _12864_/A _12864_/B _12864_/C vssd1 vssd1 vccd1 vccd1 _20347_/A sky130_fd_sc_hd__nand3_4
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _14603_/A vssd1 vssd1 vccd1 vccd1 _14916_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18371_ _22950_/Q _18369_/B _18370_/Y vssd1 vssd1 vccd1 vccd1 _22950_/D sky130_fd_sc_hd__o21a_1
XFILLER_221_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11815_ _11815_/A vssd1 vssd1 vccd1 vccd1 _11815_/X sky130_fd_sc_hd__buf_8
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _12906_/A _12795_/B vssd1 vssd1 vccd1 vccd1 _12795_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _15583_/A vssd1 vssd1 vccd1 vccd1 _15583_/X sky130_fd_sc_hd__buf_2
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_310_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _22585_/Q vssd1 vssd1 vccd1 vccd1 _17322_/Y sky130_fd_sc_hd__inv_2
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _22272_/Q _23088_/Q _23504_/Q _22433_/Q _11745_/X _12014_/A vssd1 vssd1 vccd1
+ vccd1 _11746_/X sky130_fd_sc_hd__mux4_1
X_14534_ _19163_/A vssd1 vssd1 vccd1 vccd1 _14534_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_348_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17253_ _17242_/X _17243_/X _17252_/X _17237_/X vssd1 vssd1 vccd1 vccd1 _17253_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11677_ _22471_/Q _22631_/Q _22310_/Q _23446_/Q _12716_/A _12844_/A vssd1 vssd1 vccd1
+ vccd1 _11677_/X sky130_fd_sc_hd__mux4_1
X_14465_ _14465_/A _14465_/B _14465_/C _14451_/B vssd1 vssd1 vccd1 vccd1 _14601_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_329_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16204_ _16457_/B _16310_/A vssd1 vssd1 vccd1 vccd1 _19699_/B sky130_fd_sc_hd__or2_4
XFILLER_317_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13416_ _13436_/A vssd1 vssd1 vccd1 vccd1 _20205_/A sky130_fd_sc_hd__buf_4
X_17184_ _15671_/X _17183_/X _17234_/S vssd1 vssd1 vccd1 vccd1 _17184_/X sky130_fd_sc_hd__mux2_1
X_14396_ _14393_/X _16936_/C _14421_/S vssd1 vssd1 vccd1 vccd1 _14467_/C sky130_fd_sc_hd__mux2_2
XFILLER_174_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_316_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16135_ _23619_/Q vssd1 vssd1 vccd1 vccd1 _20034_/B sky130_fd_sc_hd__buf_2
XFILLER_317_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13347_ _13618_/A _13351_/B _12168_/Y vssd1 vssd1 vccd1 vccd1 _13348_/B sky130_fd_sc_hd__a21bo_1
XFILLER_182_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_294_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_332_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13278_ _13278_/A _13278_/B vssd1 vssd1 vccd1 vccd1 _13278_/Y sky130_fd_sc_hd__nor2_1
X_16066_ _23777_/Q _15595_/X _15596_/X _16064_/X _16065_/X vssd1 vssd1 vccd1 vccd1
+ _16066_/X sky130_fd_sc_hd__a221o_2
XFILLER_335_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_331_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_335_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12229_ _12519_/A _12229_/B _12229_/C vssd1 vssd1 vccd1 vccd1 _21517_/A sky130_fd_sc_hd__and3_4
X_15017_ _15017_/A vssd1 vssd1 vccd1 vccd1 _15017_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_300_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19825_ _19825_/A vssd1 vssd1 vccd1 vccd1 _23548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_271_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19756_ _19756_/A vssd1 vssd1 vccd1 vccd1 _19765_/S sky130_fd_sc_hd__buf_6
X_16968_ _16996_/A vssd1 vssd1 vccd1 vccd1 _16968_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18707_ _18707_/A vssd1 vssd1 vccd1 vccd1 _23080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15919_ _16057_/A _15137_/X _15918_/X _13439_/A vssd1 vssd1 vccd1 vccd1 _15920_/C
+ sky130_fd_sc_hd__o22a_1
X_19687_ _19249_/X _23487_/Q _19693_/S vssd1 vssd1 vccd1 vccd1 _19688_/A sky130_fd_sc_hd__mux2_1
XFILLER_271_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16899_ _19249_/A vssd1 vssd1 vccd1 vccd1 _16899_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18638_ _18695_/S vssd1 vssd1 vccd1 vccd1 _18647_/S sky130_fd_sc_hd__buf_6
XFILLER_37_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18569_ _16835_/X _23019_/Q _18575_/S vssd1 vssd1 vccd1 vccd1 _18570_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20600_ _13910_/X _20563_/X _20599_/X vssd1 vssd1 vccd1 vccd1 _20601_/C sky130_fd_sc_hd__o21a_1
XFILLER_33_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_339_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21580_ _13960_/X _21561_/X _21568_/X _21579_/Y vssd1 vssd1 vccd1 vccd1 _21580_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_296_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20531_ _20531_/A _20531_/B vssd1 vssd1 vccd1 vccd1 _21093_/A sky130_fd_sc_hd__nor2_4
XFILLER_221_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_308_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23250_ _23474_/CLK _23250_/D vssd1 vssd1 vccd1 vccd1 _23250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20462_ _23703_/Q _20413_/X _20461_/Y _20459_/X vssd1 vssd1 vccd1 vccd1 _23703_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_319_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_335_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22201_ _22177_/B _22183_/B _22182_/A _22177_/A vssd1 vssd1 vccd1 vccd1 _22207_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_323_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23181_ _23407_/CLK _23181_/D vssd1 vssd1 vccd1 vccd1 _23181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_334_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20393_ _20213_/A _20754_/A _20391_/X _20392_/X vssd1 vssd1 vccd1 vccd1 _23682_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_335_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_323_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_334_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22132_ _22151_/A _23774_/Q vssd1 vssd1 vccd1 vccd1 _22134_/A sky130_fd_sc_hd__nor2_1
XTAP_7319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_323_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_350_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22063_ _22064_/A _22067_/A vssd1 vssd1 vccd1 vccd1 _22065_/A sky130_fd_sc_hd__nand2_1
XTAP_6629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput285 _14084_/X vssd1 vssd1 vccd1 vccd1 addr0[0] sky130_fd_sc_hd__buf_2
XFILLER_87_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_288_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput296 _13990_/Y vssd1 vssd1 vccd1 vccd1 addr1[2] sky130_fd_sc_hd__buf_2
X_21014_ _23820_/Q _20993_/X _21013_/Y _21010_/X vssd1 vssd1 vccd1 vccd1 _23820_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_3 _22139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_287_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_302_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22965_ _23696_/CLK _22965_/D vssd1 vssd1 vccd1 vccd1 _22965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21916_ _21916_/A _21920_/A vssd1 vssd1 vccd1 vccd1 _21918_/A sky130_fd_sc_hd__nand2_1
X_22896_ _23424_/CLK _22896_/D vssd1 vssd1 vccd1 vccd1 _22896_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_244_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21847_ _21847_/A vssd1 vssd1 vccd1 vccd1 _22048_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_358_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11600_ _12698_/A _11587_/Y _11594_/Y _11599_/Y vssd1 vssd1 vccd1 vccd1 _11600_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12580_ _23305_/Q _23273_/Q _23241_/Q _23529_/Q _12324_/X _12329_/X vssd1 vssd1 vccd1
+ vccd1 _12581_/B sky130_fd_sc_hd__mux4_1
XFILLER_358_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21778_ _21799_/B _21778_/B vssd1 vssd1 vccd1 vccd1 _21801_/D sky130_fd_sc_hd__nor2_2
XFILLER_196_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11531_ _13229_/A vssd1 vssd1 vccd1 vccd1 _13180_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23517_ _23547_/CLK _23517_/D vssd1 vssd1 vccd1 vccd1 _23517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20729_ _20729_/A vssd1 vssd1 vccd1 vccd1 _20729_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_345_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14250_ _14250_/A vssd1 vssd1 vccd1 vccd1 _14835_/A sky130_fd_sc_hd__buf_4
X_23448_ _23448_/CLK _23448_/D vssd1 vssd1 vccd1 vccd1 _23448_/Q sky130_fd_sc_hd__dfxtp_1
X_11462_ _11469_/A vssd1 vssd1 vccd1 vccd1 _11462_/X sky130_fd_sc_hd__buf_2
XFILLER_109_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ _22285_/Q _23101_/Q _23517_/Q _22446_/Q _13090_/S _13195_/X vssd1 vssd1 vccd1
+ vccd1 _13202_/B sky130_fd_sc_hd__mux4_1
XFILLER_326_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14181_ _14175_/Y _14177_/Y _20533_/A vssd1 vssd1 vccd1 vccd1 _14370_/C sky130_fd_sc_hd__a21bo_1
XFILLER_341_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23379_ _23507_/CLK _23379_/D vssd1 vssd1 vccd1 vccd1 _23379_/Q sky130_fd_sc_hd__dfxtp_1
X_11393_ _11394_/A _14356_/B vssd1 vssd1 vccd1 vccd1 _13314_/A sky130_fd_sc_hd__or2_1
XFILLER_326_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_314_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13132_ _22480_/Q _22640_/Q _22319_/Q _23455_/Q _13114_/X _13115_/X vssd1 vssd1 vccd1
+ vccd1 _13132_/X sky130_fd_sc_hd__mux4_2
XFILLER_353_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_297_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17940_ _22824_/Q _17938_/X _17939_/X input264/X _17933_/X vssd1 vssd1 vccd1 vccd1
+ _17940_/X sky130_fd_sc_hd__a221o_1
XFILLER_341_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13063_ _23328_/Q _23296_/Q _23264_/Q _23552_/Q _11543_/X _13276_/A vssd1 vssd1 vccd1
+ vccd1 _13064_/B sky130_fd_sc_hd__mux4_1
XFILLER_340_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_340_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12014_ _12014_/A vssd1 vssd1 vccd1 vccd1 _12710_/A sky130_fd_sc_hd__buf_6
XFILLER_305_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17871_ _17871_/A vssd1 vssd1 vccd1 vccd1 _22806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19610_ _23453_/Q _19242_/A _19610_/S vssd1 vssd1 vccd1 vccd1 _19611_/A sky130_fd_sc_hd__mux2_1
XFILLER_266_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16822_ _19172_/A vssd1 vssd1 vccd1 vccd1 _16822_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_294_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19541_ _19245_/X _23422_/Q _19549_/S vssd1 vssd1 vccd1 vccd1 _19542_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16753_ _16759_/A _16753_/B vssd1 vssd1 vccd1 vccd1 _16754_/A sky130_fd_sc_hd__or2_1
XFILLER_19_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13965_ _13965_/A _13965_/B vssd1 vssd1 vccd1 vccd1 _13965_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_321_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15704_ _15891_/A _15677_/Y _15699_/X _15703_/Y _15818_/A vssd1 vssd1 vccd1 vccd1
+ _15704_/X sky130_fd_sc_hd__o311a_1
X_19472_ _19472_/A vssd1 vssd1 vccd1 vccd1 _23391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12916_ _12916_/A _12916_/B vssd1 vssd1 vccd1 vccd1 _13492_/B sky130_fd_sc_hd__nor2_2
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16684_ input42/X _16680_/A _17382_/A vssd1 vssd1 vccd1 vccd1 _16779_/A sky130_fd_sc_hd__a21o_4
XFILLER_46_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13896_ _13505_/X _13464_/B _13506_/X vssd1 vssd1 vccd1 vccd1 _13897_/B sky130_fd_sc_hd__a21o_1
XFILLER_326_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18423_ _18423_/A vssd1 vssd1 vccd1 vccd1 _18423_/X sky130_fd_sc_hd__buf_4
XFILLER_261_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_321_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15635_ _15635_/A _15718_/B vssd1 vssd1 vccd1 vccd1 _15635_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _12852_/A vssd1 vssd1 vccd1 vccd1 _12897_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18354_ _16168_/A _18357_/C _18337_/X vssd1 vssd1 vccd1 vccd1 _18354_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_221_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ _15818_/A _13615_/Y _15574_/A vssd1 vssd1 vccd1 vccd1 _15566_/X sky130_fd_sc_hd__o21a_1
XFILLER_348_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12778_ _22279_/Q _23095_/Q _23511_/Q _22440_/Q _12776_/X _12777_/X vssd1 vssd1 vccd1
+ vccd1 _12779_/B sky130_fd_sc_hd__mux4_2
XFILLER_221_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17305_ input101/X input66/X _17314_/S vssd1 vssd1 vccd1 vccd1 _17305_/X sky130_fd_sc_hd__mux2_8
X_14517_ _14936_/A vssd1 vssd1 vccd1 vccd1 _14518_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_203_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_348_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18285_ _18286_/A _18286_/C _22922_/Q vssd1 vssd1 vccd1 vccd1 _18287_/B sky130_fd_sc_hd__a21oi_1
X_11729_ _12157_/S _13500_/B vssd1 vssd1 vccd1 vccd1 _13521_/A sky130_fd_sc_hd__and2_1
XFILLER_30_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15497_ _13386_/A _15718_/B _15496_/Y vssd1 vssd1 vccd1 vccd1 _15497_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_147_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17236_ _17169_/A _17235_/X _17195_/X _17215_/X vssd1 vssd1 vccd1 vccd1 _17236_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14448_ _14731_/A vssd1 vssd1 vccd1 vccd1 _15589_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17167_ _17167_/A vssd1 vssd1 vccd1 vccd1 _17167_/X sky130_fd_sc_hd__buf_2
XFILLER_162_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14379_ _15385_/S _14377_/X _14767_/A vssd1 vssd1 vccd1 vccd1 _14380_/A sky130_fd_sc_hd__o21a_1
XFILLER_116_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_317_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_305_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_304_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16118_ _16118_/A vssd1 vssd1 vccd1 vccd1 _21076_/A sky130_fd_sc_hd__buf_6
XFILLER_6_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_346_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17098_ _13951_/B _17096_/X _17137_/S vssd1 vssd1 vccd1 vccd1 _17098_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_304_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_288_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16049_ _19252_/A vssd1 vssd1 vccd1 vccd1 _16049_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_276_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19808_ _19808_/A vssd1 vssd1 vccd1 vccd1 _23540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_300_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19739_ _19220_/X _23510_/Q _19743_/S vssd1 vssd1 vccd1 vccd1 _19740_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22750_ _23048_/CLK _22750_/D vssd1 vssd1 vccd1 vccd1 _22750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21701_ _23825_/Q _23759_/Q vssd1 vssd1 vccd1 vccd1 _21703_/A sky130_fd_sc_hd__and2_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22681_ _23048_/CLK _22681_/D vssd1 vssd1 vccd1 vccd1 _22681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21632_ _21632_/A _21632_/B vssd1 vssd1 vccd1 vccd1 _21632_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_197_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_327_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21563_ _23821_/Q _23755_/Q vssd1 vssd1 vccd1 vccd1 _21563_/Y sky130_fd_sc_hd__nand2_1
XFILLER_139_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23302_ _23494_/CLK _23302_/D vssd1 vssd1 vccd1 vccd1 _23302_/Q sky130_fd_sc_hd__dfxtp_1
X_20514_ _23708_/Q _20524_/B _20514_/C vssd1 vssd1 vccd1 vccd1 _20515_/D sky130_fd_sc_hd__and3_1
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21494_ _21494_/A _21494_/B vssd1 vssd1 vccd1 vccd1 _21496_/A sky130_fd_sc_hd__nand2_1
XFILLER_176_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23233_ _23451_/CLK _23233_/D vssd1 vssd1 vccd1 vccd1 _23233_/Q sky130_fd_sc_hd__dfxtp_1
X_20445_ _20445_/A vssd1 vssd1 vccd1 vccd1 _20445_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_238_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23164_ _23420_/CLK _23164_/D vssd1 vssd1 vccd1 vccd1 _23164_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_7105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20376_ _20376_/A _20376_/B vssd1 vssd1 vccd1 vccd1 _20376_/Y sky130_fd_sc_hd__nor2_1
XTAP_7116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_7138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22115_ _22115_/A _22114_/Y vssd1 vssd1 vccd1 vccd1 _22118_/A sky130_fd_sc_hd__or2b_1
XFILLER_134_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_7149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23095_ _23511_/CLK _23095_/D vssd1 vssd1 vccd1 vccd1 _23095_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_322_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22046_ _22046_/A vssd1 vssd1 vccd1 vccd1 _22046_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_310_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_290_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_290_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13750_ _15576_/A _13831_/B vssd1 vssd1 vccd1 vccd1 _15113_/A sky130_fd_sc_hd__nand2_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22948_ _23602_/CLK _22948_/D vssd1 vssd1 vccd1 vccd1 _22948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_290_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12701_ _12919_/A _12699_/X _12700_/X vssd1 vssd1 vccd1 vccd1 _12701_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_271_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13681_ _13890_/B _13831_/B vssd1 vssd1 vccd1 vccd1 _15901_/A sky130_fd_sc_hd__nor2_2
XFILLER_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22879_ _23584_/CLK _22879_/D vssd1 vssd1 vccd1 vccd1 _22879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15420_ _15415_/X _21708_/B _15708_/S vssd1 vssd1 vccd1 vccd1 _18811_/A sky130_fd_sc_hd__mux2_8
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12632_ _12708_/A _12631_/X _12721_/A vssd1 vssd1 vccd1 vccd1 _12632_/Y sky130_fd_sc_hd__o21ai_1
XPHY_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15351_ _15351_/A _16070_/A vssd1 vssd1 vccd1 vccd1 _15351_/X sky130_fd_sc_hd__or2_1
XFILLER_212_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12563_ _11780_/X _12553_/X _12558_/X _12562_/X _11243_/A vssd1 vssd1 vccd1 vccd1
+ _13718_/B sky130_fd_sc_hd__a311o_4
XPHY_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_346_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14302_ _14300_/X _14301_/X _14310_/S vssd1 vssd1 vccd1 vccd1 _14302_/X sky130_fd_sc_hd__mux2_1
X_11514_ _23940_/Q vssd1 vssd1 vccd1 vccd1 _16114_/A sky130_fd_sc_hd__clkinv_2
X_18070_ _22860_/Q _18067_/X _18068_/X _22993_/Q _18069_/X vssd1 vssd1 vccd1 vccd1
+ _18070_/X sky130_fd_sc_hd__a221o_1
XFILLER_141_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_345_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15282_ _18801_/A vssd1 vssd1 vccd1 vccd1 _19194_/A sky130_fd_sc_hd__clkbuf_2
X_12494_ _23912_/Q _12520_/S vssd1 vssd1 vccd1 vccd1 _12494_/X sky130_fd_sc_hd__or2_1
XFILLER_346_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17021_ _17033_/B _17019_/X _17020_/Y _16951_/A vssd1 vssd1 vccd1 vccd1 _17021_/X
+ sky130_fd_sc_hd__o211a_1
X_14233_ _15030_/S vssd1 vssd1 vccd1 vccd1 _15033_/S sky130_fd_sc_hd__clkbuf_4
X_11445_ _22387_/Q _22419_/Q _22708_/Q _23075_/Q _11493_/S _11169_/A vssd1 vssd1 vccd1
+ vccd1 _11446_/B sky130_fd_sc_hd__mux4_2
XFILLER_50_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14164_ _14164_/A vssd1 vssd1 vccd1 vccd1 _14164_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_299_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11376_ _11826_/A vssd1 vssd1 vccd1 vccd1 _11657_/A sky130_fd_sc_hd__buf_4
XFILLER_313_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_299_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13115_ _13127_/A vssd1 vssd1 vccd1 vccd1 _13115_/X sky130_fd_sc_hd__buf_2
XFILLER_252_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14095_ _14095_/A vssd1 vssd1 vccd1 vccd1 _14095_/Y sky130_fd_sc_hd__inv_2
X_18972_ _18972_/A vssd1 vssd1 vccd1 vccd1 _23183_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_316_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_341_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17923_ _22819_/Q _17922_/X _17918_/X input260/X _17915_/X vssd1 vssd1 vccd1 vccd1
+ _17923_/X sky130_fd_sc_hd__a221o_1
X_13046_ _13107_/A _13046_/B vssd1 vssd1 vccd1 vccd1 _13046_/Y sky130_fd_sc_hd__nor2_1
XFILLER_279_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_316_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17854_ _17854_/A vssd1 vssd1 vccd1 vccd1 _22798_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_332_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16805_ _16805_/A vssd1 vssd1 vccd1 vccd1 _22518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_281_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17785_ _22768_/Q _17620_/X _17787_/S vssd1 vssd1 vccd1 vccd1 _17786_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14997_ _23690_/Q _14905_/X _14996_/X vssd1 vssd1 vccd1 vccd1 _14997_/X sky130_fd_sc_hd__o21a_2
XFILLER_94_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19524_ _19524_/A vssd1 vssd1 vccd1 vccd1 _23414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16736_ _16736_/A vssd1 vssd1 vccd1 vccd1 _22498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13948_ _13948_/A _13948_/B vssd1 vssd1 vccd1 vccd1 _13948_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_223_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19455_ _23384_/Q _18833_/X _19455_/S vssd1 vssd1 vccd1 vccd1 _19456_/A sky130_fd_sc_hd__mux2_1
X_16667_ _22480_/Q _16291_/X _16673_/S vssd1 vssd1 vccd1 vccd1 _16668_/A sky130_fd_sc_hd__mux2_1
X_13879_ _13879_/A _13879_/B vssd1 vssd1 vccd1 vccd1 _14246_/A sky130_fd_sc_hd__or2_4
XFILLER_90_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18406_ _15644_/A _18409_/C _18405_/Y vssd1 vssd1 vccd1 vccd1 _22963_/D sky130_fd_sc_hd__o21a_1
XFILLER_179_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15618_ _15618_/A vssd1 vssd1 vccd1 vccd1 _15618_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19386_ _23353_/Q _18836_/X _19394_/S vssd1 vssd1 vccd1 vccd1 _19387_/A sky130_fd_sc_hd__mux2_1
X_16598_ _16598_/A vssd1 vssd1 vccd1 vccd1 _22449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_349_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_349_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18337_ _18423_/A vssd1 vssd1 vccd1 vccd1 _18337_/X sky130_fd_sc_hd__buf_2
XFILLER_309_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15549_ _23604_/Q _14901_/A _14902_/A _23636_/Q vssd1 vssd1 vccd1 vccd1 _15549_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_277_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18268_ _18268_/A _18275_/C vssd1 vssd1 vccd1 vccd1 _18268_/Y sky130_fd_sc_hd__nor2_1
XFILLER_348_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17219_ input92/X input57/X _17219_/S vssd1 vssd1 vccd1 vccd1 _17219_/X sky130_fd_sc_hd__mux2_8
XFILLER_129_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_357_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18199_ _23012_/Q vssd1 vssd1 vccd1 vccd1 _18549_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_144_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20230_ _20227_/X _20228_/Y _20229_/X _20196_/X vssd1 vssd1 vccd1 vccd1 _20230_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_332_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_304_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_293_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_289_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20161_ _20161_/A _21097_/B vssd1 vssd1 vccd1 vccd1 _20344_/A sky130_fd_sc_hd__nor2_2
XFILLER_226_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_320_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20092_ _20098_/C _20098_/D _20091_/Y vssd1 vssd1 vccd1 vccd1 _23638_/D sky130_fd_sc_hd__a21oi_1
XFILLER_226_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_276_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_301_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23920_ _23935_/CLK _23920_/D vssd1 vssd1 vccd1 vccd1 _23920_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_58_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_301_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23851_ _23851_/CLK _23851_/D vssd1 vssd1 vccd1 vccd1 _23851_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22802_ _23070_/CLK _22802_/D vssd1 vssd1 vccd1 vccd1 _22802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_272_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23782_ _23911_/CLK _23782_/D vssd1 vssd1 vccd1 vccd1 _23782_/Q sky130_fd_sc_hd__dfxtp_4
X_20994_ _21051_/A vssd1 vssd1 vccd1 vccd1 _21072_/B sky130_fd_sc_hd__clkbuf_4
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22733_ _23068_/CLK _22733_/D vssd1 vssd1 vccd1 vccd1 _22733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22664_ _23575_/CLK _22664_/D vssd1 vssd1 vccd1 vccd1 _22664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21615_ _21615_/A vssd1 vssd1 vccd1 vccd1 _21870_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_231_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22595_ _22600_/CLK _22595_/D vssd1 vssd1 vccd1 vccd1 _22595_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_328_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_327_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21546_ _21546_/A _21546_/B vssd1 vssd1 vccd1 vccd1 _21546_/X sky130_fd_sc_hd__and2_1
XFILLER_139_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_355_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21477_ _13960_/X _21455_/X _21464_/X _21476_/Y vssd1 vssd1 vccd1 vccd1 _21477_/X
+ sky130_fd_sc_hd__a211o_1
X_23216_ _23474_/CLK _23216_/D vssd1 vssd1 vccd1 vccd1 _23216_/Q sky130_fd_sc_hd__dfxtp_1
X_11230_ _11230_/A vssd1 vssd1 vccd1 vccd1 _11965_/A sky130_fd_sc_hd__buf_4
XFILLER_355_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20428_ _20428_/A vssd1 vssd1 vccd1 vccd1 _20428_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_355_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23147_ _23531_/CLK _23147_/D vssd1 vssd1 vccd1 vccd1 _23147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11161_ _12425_/A vssd1 vssd1 vccd1 vccd1 _12246_/A sky130_fd_sc_hd__buf_2
XFILLER_122_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20359_ _20963_/A vssd1 vssd1 vccd1 vccd1 _20445_/A sky130_fd_sc_hd__clkbuf_4
XTAP_6201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_323_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ _13472_/A vssd1 vssd1 vccd1 vccd1 _13779_/A sky130_fd_sc_hd__buf_12
X_23078_ _23494_/CLK _23078_/D vssd1 vssd1 vccd1 vccd1 _23078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_310_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22029_ _22029_/A _22032_/A vssd1 vssd1 vccd1 vccd1 _22030_/B sky130_fd_sc_hd__nor2_1
X_14920_ _23785_/Q _14917_/X _14919_/X vssd1 vssd1 vccd1 vccd1 _14920_/X sky130_fd_sc_hd__a21o_1
XTAP_6289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14851_ _14638_/X _14643_/X _14853_/S vssd1 vssd1 vccd1 vccd1 _14851_/X sky130_fd_sc_hd__mux2_1
XFILLER_275_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13802_ _13802_/A vssd1 vssd1 vccd1 vccd1 _13802_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17570_ _22685_/Q _17569_/X _17576_/S vssd1 vssd1 vccd1 vccd1 _17571_/A sky130_fd_sc_hd__mux2_1
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14782_ _14331_/X _14299_/X _14841_/S vssd1 vssd1 vccd1 vccd1 _14782_/X sky130_fd_sc_hd__mux2_1
X_11994_ _22372_/Q _22404_/Q _22693_/Q _23060_/Q _12716_/A _12844_/A vssd1 vssd1 vccd1
+ vccd1 _11994_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16521_ _16521_/A vssd1 vssd1 vccd1 vccd1 _22416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_302_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13733_ _13765_/C _13777_/B vssd1 vssd1 vccd1 vccd1 _13745_/B sky130_fd_sc_hd__nor2_1
XFILLER_16_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_290_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23474_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_43_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19240_ _19239_/X _23292_/Q _19243_/S vssd1 vssd1 vccd1 vccd1 _19241_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16452_ _16452_/A vssd1 vssd1 vccd1 vccd1 _22386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13664_ _22604_/Q _22605_/Q _22606_/Q vssd1 vssd1 vccd1 vccd1 _13670_/C sky130_fd_sc_hd__or3_4
XFILLER_204_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15403_ _23697_/Q _14491_/A _15402_/X vssd1 vssd1 vccd1 vccd1 _15403_/Y sky130_fd_sc_hd__o21ai_4
X_12615_ _23317_/Q _23285_/Q _23253_/Q _23541_/Q _12008_/X _12009_/X vssd1 vssd1 vccd1
+ vccd1 _12616_/B sky130_fd_sc_hd__mux4_2
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19171_ _19171_/A vssd1 vssd1 vccd1 vccd1 _23270_/D sky130_fd_sc_hd__clkbuf_1
X_16383_ _19627_/A vssd1 vssd1 vccd1 vccd1 _19267_/A sky130_fd_sc_hd__clkbuf_4
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ _17229_/A _13884_/A _13592_/Y _14198_/B vssd1 vssd1 vccd1 vccd1 _13977_/A
+ sky130_fd_sc_hd__a22o_4
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18122_ _18116_/Y _18117_/X _18119_/X _18121_/X vssd1 vssd1 vccd1 vccd1 _22878_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15334_ _14829_/Y _15181_/X _15183_/X _15333_/Y vssd1 vssd1 vccd1 vccd1 _21233_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_40_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12546_ _12546_/A _13362_/B _13361_/B vssd1 vssd1 vccd1 vccd1 _14687_/B sky130_fd_sc_hd__or3b_2
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18053_ _18053_/A vssd1 vssd1 vccd1 vccd1 _18053_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_185_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15265_ _23758_/Q _15215_/X _15216_/X _15263_/X _15264_/X vssd1 vssd1 vccd1 vccd1
+ _15265_/X sky130_fd_sc_hd__a221o_1
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12477_ _23462_/Q _23558_/Q _22522_/Q _22326_/Q _12475_/X _12476_/X vssd1 vssd1 vccd1
+ vccd1 _12477_/X sky130_fd_sc_hd__mux4_1
X_17004_ _20524_/B vssd1 vssd1 vccd1 vccd1 _20508_/B sky130_fd_sc_hd__buf_6
X_14216_ _14216_/A _14216_/B vssd1 vssd1 vccd1 vccd1 _15109_/A sky130_fd_sc_hd__or2_1
X_11428_ _13084_/A vssd1 vssd1 vccd1 vccd1 _13095_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_172_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15196_ _15460_/B vssd1 vssd1 vccd1 vccd1 _15196_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_99_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_342_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_299_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14147_ _14211_/A _14147_/B vssd1 vssd1 vccd1 vccd1 _16971_/B sky130_fd_sc_hd__nor2_2
X_11359_ _12519_/A vssd1 vssd1 vccd1 vccd1 _12594_/A sky130_fd_sc_hd__buf_6
XFILLER_302_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_298_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_301_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_302_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14078_ _15056_/A vssd1 vssd1 vccd1 vccd1 _14724_/A sky130_fd_sc_hd__clkbuf_4
X_18955_ _16825_/X _23176_/Q _18957_/S vssd1 vssd1 vccd1 vccd1 _18956_/A sky130_fd_sc_hd__mux2_1
XFILLER_258_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_343_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17906_ _22814_/Q _17894_/X _17903_/X input255/X _17899_/X vssd1 vssd1 vccd1 vccd1
+ _17906_/X sky130_fd_sc_hd__a221o_1
X_13029_ _13029_/A _13029_/B vssd1 vssd1 vccd1 vccd1 _13029_/Y sky130_fd_sc_hd__nand2_1
XFILLER_343_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_295_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18886_ _18886_/A vssd1 vssd1 vccd1 vccd1 _23145_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_267_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17837_ _22791_/Q _17591_/X _17837_/S vssd1 vssd1 vccd1 vccd1 _17838_/A sky130_fd_sc_hd__mux2_1
XFILLER_266_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17768_ _22760_/Q _17594_/X _17776_/S vssd1 vssd1 vccd1 vccd1 _17769_/A sky130_fd_sc_hd__mux2_1
XFILLER_270_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19507_ _19553_/S vssd1 vssd1 vccd1 vccd1 _19516_/S sky130_fd_sc_hd__buf_4
X_16719_ _22494_/Q _16711_/X _16712_/X input39/X vssd1 vssd1 vccd1 vccd1 _16720_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_35_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17699_ _17699_/A vssd1 vssd1 vccd1 vccd1 _22729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_430 _22887_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_441 _23916_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_452 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19438_ _23376_/Q _18808_/X _19444_/S vssd1 vssd1 vccd1 vccd1 _19439_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_463 _20754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_357_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_474 _20234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_485 _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_496 _14235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_356_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_298_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19369_ _19369_/A vssd1 vssd1 vccd1 vccd1 _23345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21400_ _21400_/A _21406_/A vssd1 vssd1 vccd1 vccd1 _21400_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22380_ _23449_/CLK _22380_/D vssd1 vssd1 vccd1 vccd1 _22380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_309_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21331_ _21317_/A _21305_/X _21330_/Y _21281_/X vssd1 vssd1 vccd1 vccd1 _23912_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_336_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_351_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21262_ _21262_/A vssd1 vssd1 vccd1 vccd1 _23900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_274_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_351_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23001_ _23592_/CLK _23001_/D vssd1 vssd1 vccd1 vccd1 _23001_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_144_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20213_ _20213_/A vssd1 vssd1 vccd1 vccd1 _20213_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21193_ _21193_/A _21308_/B _21193_/C vssd1 vssd1 vccd1 vccd1 _21260_/S sky130_fd_sc_hd__and3_2
XFILLER_104_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_305_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20144_ _20161_/A _20890_/B vssd1 vssd1 vccd1 vccd1 _20333_/A sky130_fd_sc_hd__or2_1
XFILLER_131_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20075_ _23633_/Q _20072_/B _20074_/Y vssd1 vssd1 vccd1 vccd1 _23633_/D sky130_fd_sc_hd__o21a_1
XFILLER_292_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_301_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23903_ _23903_/CLK _23903_/D vssd1 vssd1 vccd1 vccd1 _23903_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23834_ _23876_/CLK _23834_/D vssd1 vssd1 vccd1 vccd1 _23834_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_73_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23765_ _23768_/CLK _23765_/D vssd1 vssd1 vccd1 vccd1 _23765_/Q sky130_fd_sc_hd__dfxtp_2
X_20977_ _22166_/A _20966_/X _20752_/B _20970_/X vssd1 vssd1 vccd1 vccd1 _20977_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22716_ _23048_/CLK _22716_/D vssd1 vssd1 vccd1 vccd1 _22716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_348_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23696_ _23696_/CLK _23696_/D vssd1 vssd1 vccd1 vccd1 _23696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22647_ _23496_/CLK _22647_/D vssd1 vssd1 vccd1 vccd1 _22647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_348_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12400_ _23303_/Q _23271_/Q _23239_/Q _23527_/Q _11647_/A _12269_/X vssd1 vssd1 vccd1
+ vccd1 _12401_/B sky130_fd_sc_hd__mux4_1
XFILLER_139_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13380_ _13380_/A vssd1 vssd1 vccd1 vccd1 _13948_/A sky130_fd_sc_hd__buf_4
X_22578_ _23643_/CLK _22578_/D vssd1 vssd1 vccd1 vccd1 _22578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_316_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12331_ _12590_/A _12331_/B vssd1 vssd1 vccd1 vccd1 _12331_/X sky130_fd_sc_hd__or2_1
XFILLER_355_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21529_ _23788_/Q _21683_/A _21528_/Y _21346_/A vssd1 vssd1 vccd1 vccd1 _21529_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_108_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_309_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_163_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _23878_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_315_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12262_ _12135_/A _13724_/A _12261_/Y vssd1 vssd1 vccd1 vccd1 _12606_/A sky130_fd_sc_hd__a21oi_4
XFILLER_147_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15050_ _15037_/A _15049_/C _21500_/A vssd1 vssd1 vccd1 vccd1 _15051_/B sky130_fd_sc_hd__a21oi_1
XFILLER_107_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14001_ _14001_/A vssd1 vssd1 vccd1 vccd1 _14072_/C sky130_fd_sc_hd__clkbuf_2
X_11213_ _11240_/A vssd1 vssd1 vccd1 vccd1 _11214_/A sky130_fd_sc_hd__buf_4
XFILLER_108_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12193_ _12244_/A vssd1 vssd1 vccd1 vccd1 _12242_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_269_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_323_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11144_ _13199_/A vssd1 vssd1 vccd1 vccd1 _13041_/A sky130_fd_sc_hd__buf_4
XTAP_6020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_6031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_296_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18740_ _18740_/A vssd1 vssd1 vccd1 vccd1 _23095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_311_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15952_ _22971_/Q _16144_/S vssd1 vssd1 vccd1 vccd1 _15952_/X sky130_fd_sc_hd__or2_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11075_ _14172_/B vssd1 vssd1 vccd1 vccd1 _13440_/B sky130_fd_sc_hd__buf_4
XTAP_6075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput130 dout1[30] vssd1 vssd1 vccd1 vccd1 input130/X sky130_fd_sc_hd__clkbuf_1
XTAP_6086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput141 dout1[40] vssd1 vssd1 vccd1 vccd1 input141/X sky130_fd_sc_hd__buf_2
XTAP_6097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput152 dout1[50] vssd1 vssd1 vccd1 vccd1 input152/X sky130_fd_sc_hd__buf_2
X_14903_ _23593_/Q _14901_/X _14902_/X _23625_/Q vssd1 vssd1 vccd1 vccd1 _14903_/X
+ sky130_fd_sc_hd__o22a_2
XTAP_5363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput163 dout1[60] vssd1 vssd1 vccd1 vccd1 input163/X sky130_fd_sc_hd__buf_2
XTAP_5374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18671_ _18682_/A vssd1 vssd1 vccd1 vccd1 _18680_/S sky130_fd_sc_hd__buf_2
XTAP_5385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _23708_/Q _14905_/X _15882_/X vssd1 vssd1 vccd1 vccd1 _15883_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_248_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput174 irq[12] vssd1 vssd1 vccd1 vccd1 _20505_/C sky130_fd_sc_hd__buf_2
XFILLER_37_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput185 irq[8] vssd1 vssd1 vccd1 vccd1 _20522_/C sky130_fd_sc_hd__buf_2
XFILLER_291_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput196 localMemory_wb_adr_i[15] vssd1 vssd1 vccd1 vccd1 input196/X sky130_fd_sc_hd__clkbuf_1
X_17622_ _17622_/A vssd1 vssd1 vccd1 vccd1 _22701_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834_ _14830_/Y _14832_/X _15865_/A vssd1 vssd1 vccd1 vccd1 _14834_/X sky130_fd_sc_hd__mux2_4
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17553_ _18779_/A vssd1 vssd1 vccd1 vccd1 _17553_/X sky130_fd_sc_hd__buf_2
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _15249_/S vssd1 vssd1 vccd1 vccd1 _15490_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11977_ _12754_/A _11976_/X _11965_/A vssd1 vssd1 vccd1 vccd1 _11977_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_189_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16504_ _16515_/A vssd1 vssd1 vccd1 vccd1 _16513_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_45_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13716_ _13716_/A vssd1 vssd1 vccd1 vccd1 _13716_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_339_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17484_ _17484_/A vssd1 vssd1 vccd1 vccd1 _22650_/D sky130_fd_sc_hd__clkbuf_1
X_14696_ _16005_/A vssd1 vssd1 vccd1 vccd1 _16191_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_205_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19223_ _19223_/A vssd1 vssd1 vccd1 vccd1 _19223_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_260_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16435_ _16435_/A vssd1 vssd1 vccd1 vccd1 _22378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13647_ _13647_/A _15335_/A vssd1 vssd1 vccd1 vccd1 _13647_/Y sky130_fd_sc_hd__nand2_1
XFILLER_258_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19154_ _19154_/A vssd1 vssd1 vccd1 vccd1 _23264_/D sky130_fd_sc_hd__clkbuf_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _15936_/X _22349_/Q _16366_/S vssd1 vssd1 vccd1 vccd1 _16367_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _13492_/X _13540_/A _13632_/B _13540_/X vssd1 vssd1 vccd1 vccd1 _13579_/B
+ sky130_fd_sc_hd__o22a_1
X_18105_ _18105_/A vssd1 vssd1 vccd1 vccd1 _18105_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_307_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_297_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15317_ _15376_/C _15317_/B vssd1 vssd1 vccd1 vccd1 _15318_/B sky130_fd_sc_hd__or2_2
XFILLER_306_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19085_ _19085_/A vssd1 vssd1 vccd1 vccd1 _23234_/D sky130_fd_sc_hd__clkbuf_1
X_12529_ _12532_/A _12529_/B vssd1 vssd1 vccd1 vccd1 _12529_/Y sky130_fd_sc_hd__nor2_1
XFILLER_334_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_319_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16297_ _18862_/A vssd1 vssd1 vccd1 vccd1 _16297_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_258_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_333_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_318_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_306_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18036_ _18052_/A vssd1 vssd1 vccd1 vccd1 _18036_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_333_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15248_ _20186_/A _13943_/A _15247_/X vssd1 vssd1 vccd1 vccd1 _15248_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_334_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_322_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_321_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_314_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15179_ _15179_/A _15901_/B vssd1 vssd1 vccd1 vccd1 _15483_/B sky130_fd_sc_hd__nor2_1
XFILLER_113_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_302_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_354_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19987_ _19987_/A vssd1 vssd1 vccd1 vccd1 _20027_/A sky130_fd_sc_hd__buf_2
XFILLER_87_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_287_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18938_ _23169_/Q _18862_/X _18940_/S vssd1 vssd1 vccd1 vccd1 _18939_/A sky130_fd_sc_hd__mux2_1
.ends

