* NGSPICE file created from SPI.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

.subckt SPI clk peripheralBus_address[0] peripheralBus_address[10] peripheralBus_address[11]
+ peripheralBus_address[12] peripheralBus_address[13] peripheralBus_address[14] peripheralBus_address[15]
+ peripheralBus_address[16] peripheralBus_address[17] peripheralBus_address[18] peripheralBus_address[19]
+ peripheralBus_address[1] peripheralBus_address[20] peripheralBus_address[21] peripheralBus_address[22]
+ peripheralBus_address[23] peripheralBus_address[2] peripheralBus_address[3] peripheralBus_address[4]
+ peripheralBus_address[5] peripheralBus_address[6] peripheralBus_address[7] peripheralBus_address[8]
+ peripheralBus_address[9] peripheralBus_busy peripheralBus_data[0] peripheralBus_data[10]
+ peripheralBus_data[11] peripheralBus_data[12] peripheralBus_data[13] peripheralBus_data[14]
+ peripheralBus_data[15] peripheralBus_data[16] peripheralBus_data[17] peripheralBus_data[18]
+ peripheralBus_data[19] peripheralBus_data[1] peripheralBus_data[20] peripheralBus_data[21]
+ peripheralBus_data[22] peripheralBus_data[23] peripheralBus_data[24] peripheralBus_data[25]
+ peripheralBus_data[26] peripheralBus_data[27] peripheralBus_data[28] peripheralBus_data[29]
+ peripheralBus_data[2] peripheralBus_data[30] peripheralBus_data[31] peripheralBus_data[3]
+ peripheralBus_data[4] peripheralBus_data[5] peripheralBus_data[6] peripheralBus_data[7]
+ peripheralBus_data[8] peripheralBus_data[9] peripheralBus_oe peripheralBus_we rst
+ spi_clk[0] spi_clk[1] spi_cs[0] spi_cs[1] spi_en[0] spi_en[1] spi_miso[0] spi_miso[1]
+ spi_mosi[0] spi_mosi[1] vccd1 vssd1
XFILLER_54_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1381__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1462__94 vssd1 vssd1 vccd1 vccd1 _1462__94/HI _1584_/A sky130_fd_sc_hd__conb_1
XFILLER_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1270_ _1270_/A vssd1 vssd1 vccd1 vccd1 _1383_/D sky130_fd_sc_hd__clkbuf_1
X_0985_ _0991_/A _0991_/B _0985_/C _0985_/D vssd1 vssd1 vccd1 vccd1 _0986_/A sky130_fd_sc_hd__or4_1
X_1606_ _1606_/A _0899_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[7] sky130_fd_sc_hd__ebufn_8
X_1537_ _1537_/A _1044_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[2] sky130_fd_sc_hd__ebufn_8
X_1399_ _1404_/CLK _1399_/D vssd1 vssd1 vccd1 vccd1 _1399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0770_ _0867_/A vssd1 vssd1 vccd1 vccd1 _0789_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1253_ _1267_/A vssd1 vssd1 vccd1 vccd1 _1253_/X sky130_fd_sc_hd__buf_2
X_1322_ _1334_/A _1322_/B vssd1 vssd1 vccd1 vccd1 _1323_/A sky130_fd_sc_hd__or2_1
X_1184_ _1184_/A vssd1 vssd1 vccd1 vccd1 _1365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0968_ _0968_/A vssd1 vssd1 vccd1 vccd1 _0968_/X sky130_fd_sc_hd__clkbuf_1
X_0899_ _0899_/A vssd1 vssd1 vccd1 vccd1 _0899_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1432__64 vssd1 vssd1 vccd1 vccd1 _1432__64/HI _1546_/A sky130_fd_sc_hd__conb_1
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1336__A0 _1185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0822_ _0891_/A vssd1 vssd1 vccd1 vccd1 _0845_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0801__A _0931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1327__A0 peripheralBus_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0753_ _0753_/A _0753_/B _0753_/C _0753_/D vssd1 vssd1 vccd1 vccd1 _0756_/B sky130_fd_sc_hd__or4_1
X_1236_ _1236_/A _1379_/Q _1236_/C vssd1 vssd1 vccd1 vccd1 _1236_/X sky130_fd_sc_hd__or3_1
X_1305_ _1303_/X _1304_/X _1305_/S vssd1 vssd1 vccd1 vccd1 _1305_/X sky130_fd_sc_hd__mux2_1
X_1167_ _1177_/A _1167_/B vssd1 vssd1 vccd1 vccd1 _1168_/A sky130_fd_sc_hd__and2_1
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1098_ _1098_/A vssd1 vssd1 vccd1 vccd1 _1098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1318__A0 peripheralBus_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487__119 vssd1 vssd1 vccd1 vccd1 _1487__119/HI _1617_/A sky130_fd_sc_hd__conb_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1021_ _1021_/A _1021_/B _1029_/C _1029_/D vssd1 vssd1 vccd1 vccd1 _1022_/A sky130_fd_sc_hd__or4_1
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0805_ _0805_/A vssd1 vssd1 vccd1 vccd1 _0805_/X sky130_fd_sc_hd__clkbuf_1
X_0736_ _0752_/A input1/X _0755_/A _0753_/A vssd1 vssd1 vccd1 vccd1 _0737_/D sky130_fd_sc_hd__or4_1
XFILLER_55_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1219_ _1269_/A _1219_/B vssd1 vssd1 vccd1 vccd1 _1220_/A sky130_fd_sc_hd__and2_1
XFILLER_25_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1211__S _1225_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input18_A peripheralBus_address[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1570_ _1570_/A _0919_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[3] sky130_fd_sc_hd__ebufn_8
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1004_ _1004_/A vssd1 vssd1 vccd1 vccd1 _1004_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1357__A _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput31 _1603_/A vssd1 vssd1 vccd1 vccd1 spi_clk[0] sky130_fd_sc_hd__buf_2
XANTENNA__1267__A _1267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1622_ _1622_/A _0839_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[23] sky130_fd_sc_hd__ebufn_8
XFILLER_8_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1553_ _1553_/A _1086_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[18] sky130_fd_sc_hd__ebufn_8
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1438__70 vssd1 vssd1 vccd1 vccd1 _1438__70/HI _1552_/A sky130_fd_sc_hd__conb_1
X_0984_ _0984_/A vssd1 vssd1 vccd1 vccd1 _0984_/X sky130_fd_sc_hd__clkbuf_1
X_1536_ _1536_/A _1042_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[1] sky130_fd_sc_hd__ebufn_8
X_1605_ _1605_/A _0897_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[6] sky130_fd_sc_hd__ebufn_8
X_1398_ _1404_/CLK _1398_/D vssd1 vssd1 vccd1 vccd1 _1606_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_63_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1280__A _1295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1371__CLK _1378_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1252_ _1404_/Q vssd1 vssd1 vccd1 vccd1 _1267_/A sky130_fd_sc_hd__clkinv_2
X_1321_ peripheralBus_data[2] _1601_/A _1333_/S vssd1 vssd1 vccd1 vccd1 _1322_/B sky130_fd_sc_hd__mux2_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1183_ _1208_/A _1183_/B vssd1 vssd1 vccd1 vccd1 _1184_/A sky130_fd_sc_hd__and2_1
XFILLER_24_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0967_ _0977_/A _0977_/B _0972_/C _0969_/D vssd1 vssd1 vccd1 vccd1 _0968_/A sky130_fd_sc_hd__or4_2
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1519_ _1519_/A _0996_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[16] sky130_fd_sc_hd__ebufn_8
X_0898_ _0904_/A _0904_/B _0898_/C _0902_/D vssd1 vssd1 vccd1 vccd1 _0899_/A sky130_fd_sc_hd__or4_1
XFILLER_59_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1275__A _1295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1394__CLK _1396_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0821_ _0821_/A vssd1 vssd1 vccd1 vccd1 _0821_/X sky130_fd_sc_hd__clkbuf_1
X_1408__40 vssd1 vssd1 vccd1 vccd1 _1408__40/HI _1514_/A sky130_fd_sc_hd__conb_1
X_0752_ _0752_/A input1/X vssd1 vssd1 vccd1 vccd1 _0756_/A sky130_fd_sc_hd__or2_1
XANTENNA__1185__A peripheralBus_data[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1166_ peripheralBus_data[3] _1144_/X _1165_/X _1155_/X vssd1 vssd1 vccd1 vccd1 _1167_/B
+ sky130_fd_sc_hd__a22o_1
X_1235_ _1233_/X _1234_/Y _1537_/A _1536_/A vssd1 vssd1 vccd1 vccd1 _1236_/C sky130_fd_sc_hd__a211o_1
X_1304_ _1568_/A _1573_/A _1604_/A vssd1 vssd1 vccd1 vccd1 _1304_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1097_ _1105_/A _1105_/B _1099_/C _1099_/D vssd1 vssd1 vccd1 vccd1 _1098_/A sky130_fd_sc_hd__or4_1
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1020_ _1020_/A vssd1 vssd1 vccd1 vccd1 _1020_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0804_ _0808_/A _0808_/B _0808_/C _0813_/D vssd1 vssd1 vccd1 vccd1 _0805_/A sky130_fd_sc_hd__or4_1
XANTENNA__0812__A _0928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0735_ _0753_/B _0753_/C _0753_/D _0754_/A vssd1 vssd1 vccd1 vccd1 _0737_/C sky130_fd_sc_hd__or4_1
X_1470__102 vssd1 vssd1 vccd1 vccd1 _1470__102/HI _1592_/A sky130_fd_sc_hd__conb_1
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1218_ peripheralBus_data[4] _1539_/A _1228_/S vssd1 vssd1 vccd1 vccd1 _1219_/B sky130_fd_sc_hd__mux2_1
XFILLER_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1149_ _1297_/A vssd1 vssd1 vccd1 vccd1 _1337_/A sky130_fd_sc_hd__buf_2
XFILLER_40_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1003_ _1005_/A _1005_/B _1015_/C _1015_/D vssd1 vssd1 vccd1 vccd1 _1004_/A sky130_fd_sc_hd__or4_1
XFILLER_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1218__A0 peripheralBus_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput32 _1539_/A vssd1 vssd1 vccd1 vccd1 spi_clk[1] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1621_ _1621_/A _0761_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[22] sky130_fd_sc_hd__ebufn_8
X_1552_ _1552_/A _1084_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[17] sky130_fd_sc_hd__ebufn_8
XFILLER_12_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0983_ _0991_/A _0991_/B _0985_/C _0985_/D vssd1 vssd1 vccd1 vccd1 _0984_/A sky130_fd_sc_hd__or4_1
X_1453__85 vssd1 vssd1 vccd1 vccd1 _1453__85/HI _1575_/A sky130_fd_sc_hd__conb_1
X_1535_ _1535_/A _0837_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[0] sky130_fd_sc_hd__ebufn_8
X_1604_ _1604_/A _0893_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[5] sky130_fd_sc_hd__ebufn_8
XANTENNA__1354__C _1354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1397_ _1404_/CLK _1397_/D vssd1 vssd1 vccd1 vccd1 _1605_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0730__A _1141_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1320_ _1320_/A vssd1 vssd1 vccd1 vccd1 _1392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1182_ peripheralBus_data[6] _1144_/A _1181_/X _1155_/A vssd1 vssd1 vccd1 vccd1 _1183_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1251_ _1247_/X _1250_/Y _1222_/A vssd1 vssd1 vccd1 vccd1 _1381_/D sky130_fd_sc_hd__a21oi_1
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0815__A _0931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0966_ _0994_/A vssd1 vssd1 vccd1 vccd1 _0977_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_0897_ _0897_/A vssd1 vssd1 vccd1 vccd1 _0897_/X sky130_fd_sc_hd__clkbuf_1
X_1518_ _1518_/A _0992_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[15] sky130_fd_sc_hd__ebufn_8
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0820_ _0823_/A _0823_/B _0854_/C _0857_/D vssd1 vssd1 vccd1 vccd1 _0821_/A sky130_fd_sc_hd__or4_1
X_1423__55 vssd1 vssd1 vccd1 vccd1 _1423__55/HI _1529_/A sky130_fd_sc_hd__conb_1
X_0751_ _0867_/A vssd1 vssd1 vccd1 vccd1 _1123_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1303_ _1567_/A _1574_/A _1604_/A vssd1 vssd1 vccd1 vccd1 _1303_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1165_ _1506_/A _1164_/X _1175_/S vssd1 vssd1 vccd1 vccd1 _1165_/X sky130_fd_sc_hd__mux2_1
X_1096_ _1096_/A vssd1 vssd1 vccd1 vccd1 _1096_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1234_ _1378_/Q _1535_/A vssd1 vssd1 vccd1 vccd1 _1234_/Y sky130_fd_sc_hd__nand2_1
X_0949_ _0949_/A vssd1 vssd1 vccd1 vccd1 _0949_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1225__S _1225_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0803_ _0803_/A vssd1 vssd1 vccd1 vccd1 _0803_/X sky130_fd_sc_hd__clkbuf_1
X_0734_ _0754_/B input3/X input2/X vssd1 vssd1 vccd1 vccd1 _0737_/B sky130_fd_sc_hd__or3_1
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1079_ _1107_/A vssd1 vssd1 vccd1 vccd1 _1091_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1148_ _1148_/A vssd1 vssd1 vccd1 vccd1 _1359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1217_ _1217_/A vssd1 vssd1 vccd1 vccd1 _1371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1384__CLK _1396_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1493__125 vssd1 vssd1 vccd1 vccd1 _1493__125/HI _1623_/A sky130_fd_sc_hd__conb_1
XFILLER_6_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1002_ _1018_/A vssd1 vssd1 vccd1 vccd1 _1015_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1459__91 vssd1 vssd1 vccd1 vccd1 _1459__91/HI _1581_/A sky130_fd_sc_hd__conb_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1477__109 vssd1 vssd1 vccd1 vccd1 _1477__109/HI _1607_/A sky130_fd_sc_hd__conb_1
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput33 _1132_/X vssd1 vssd1 vccd1 vccd1 spi_cs[0] sky130_fd_sc_hd__buf_2
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input23_A peripheralBus_address[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1620_ _1620_/A _0824_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[21] sky130_fd_sc_hd__ebufn_8
X_1551_ _1551_/A _1082_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[16] sky130_fd_sc_hd__ebufn_8
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0982_ _0982_/A vssd1 vssd1 vccd1 vccd1 _0982_/X sky130_fd_sc_hd__clkbuf_1
X_1499__131 vssd1 vssd1 vccd1 vccd1 _1499__131/HI _1629_/A sky130_fd_sc_hd__conb_1
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1534_ _1534_/A _1040_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[31] sky130_fd_sc_hd__ebufn_8
X_1603_ _1603_/A _0890_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[4] sky130_fd_sc_hd__ebufn_8
XFILLER_27_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1396_ _1396_/CLK _1396_/D vssd1 vssd1 vccd1 vccd1 _1604_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1429__61 vssd1 vssd1 vccd1 vccd1 _1429__61/HI _1543_/A sky130_fd_sc_hd__conb_1
XFILLER_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1181_ _1509_/A _1180_/X _1193_/S vssd1 vssd1 vccd1 vccd1 _1181_/X sky130_fd_sc_hd__mux2_1
X_1250_ _1381_/Q _1250_/B vssd1 vssd1 vccd1 vccd1 _1250_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0965_ _0993_/A vssd1 vssd1 vccd1 vccd1 _0977_/A sky130_fd_sc_hd__clkbuf_1
X_0896_ _0904_/A _0904_/B _0898_/C _0902_/D vssd1 vssd1 vccd1 vccd1 _0897_/A sky130_fd_sc_hd__or4_1
X_1517_ _1517_/A _0990_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[14] sky130_fd_sc_hd__ebufn_8
X_1379_ _1404_/CLK _1379_/D vssd1 vssd1 vccd1 vccd1 _1379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0750_ _1258_/C vssd1 vssd1 vccd1 vccd1 _0867_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1233_ _1378_/Q _1535_/A vssd1 vssd1 vccd1 vccd1 _1233_/X sky130_fd_sc_hd__or2_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1302_ _1302_/A vssd1 vssd1 vccd1 vccd1 _1389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1164_ _1507_/A _1505_/A _1196_/S vssd1 vssd1 vccd1 vccd1 _1164_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1095_ _1105_/A _1105_/B _1099_/C _1099_/D vssd1 vssd1 vccd1 vccd1 _1096_/A sky130_fd_sc_hd__or4_1
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0948_ _0948_/A _0948_/B _0958_/C _0954_/D vssd1 vssd1 vccd1 vccd1 _0949_/A sky130_fd_sc_hd__or4_2
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0879_ _0879_/A vssd1 vssd1 vccd1 vccd1 _0879_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0802_ _0808_/A _0808_/B _0808_/C _0813_/D vssd1 vssd1 vccd1 vccd1 _0803_/A sky130_fd_sc_hd__or4_1
X_0733_ _0755_/B vssd1 vssd1 vccd1 vccd1 _0737_/A sky130_fd_sc_hd__inv_2
XFILLER_37_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1216_ _1269_/A _1216_/B vssd1 vssd1 vccd1 vccd1 _1217_/A sky130_fd_sc_hd__and2_1
XFILLER_52_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1147_ _1147_/A _1147_/B vssd1 vssd1 vccd1 vccd1 _1148_/A sky130_fd_sc_hd__and2_1
XFILLER_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1078_ _1078_/A vssd1 vssd1 vccd1 vccd1 _1078_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1001_ _1001_/A vssd1 vssd1 vccd1 vccd1 _1015_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_34_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput34 _1130_/X vssd1 vssd1 vccd1 vccd1 spi_cs[1] sky130_fd_sc_hd__buf_2
XFILLER_48_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input16_A peripheralBus_address[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1501__133 vssd1 vssd1 vccd1 vccd1 _1501__133/HI spi_en[0] sky130_fd_sc_hd__conb_1
X_1550_ _1550_/A _1078_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[15] sky130_fd_sc_hd__ebufn_8
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1374__CLK _1378_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0834__A _1143_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input8_A peripheralBus_address[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1397__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0981_ _0991_/A _0991_/B _0985_/C _1123_/D vssd1 vssd1 vccd1 vccd1 _0982_/A sky130_fd_sc_hd__or4_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1602_ _1602_/A _0888_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[3] sky130_fd_sc_hd__ebufn_8
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1533_ _1533_/A _1036_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[30] sky130_fd_sc_hd__ebufn_8
X_1395_ _1404_/CLK _1395_/D vssd1 vssd1 vccd1 vccd1 _1603_/A sky130_fd_sc_hd__dfxtp_2
X_1444__76 vssd1 vssd1 vccd1 vccd1 _1444__76/HI _1558_/A sky130_fd_sc_hd__conb_1
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1180_ _1510_/A _1508_/A _1186_/S vssd1 vssd1 vccd1 vccd1 _1180_/X sky130_fd_sc_hd__mux2_1
X_0964_ _0964_/A vssd1 vssd1 vccd1 vccd1 _0964_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1516_ _1516_/A _0986_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[13] sky130_fd_sc_hd__ebufn_8
X_0895_ _0921_/A vssd1 vssd1 vccd1 vccd1 _0904_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1378_ _1378_/CLK _1378_/D vssd1 vssd1 vccd1 vccd1 _1378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1232_ _1380_/Q vssd1 vssd1 vccd1 vccd1 _1236_/A sky130_fd_sc_hd__inv_2
X_1301_ _1325_/A _1301_/B vssd1 vssd1 vccd1 vccd1 _1302_/A sky130_fd_sc_hd__and2_1
XFILLER_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1163_ _1163_/A vssd1 vssd1 vccd1 vccd1 _1361_/D sky130_fd_sc_hd__clkbuf_1
X_1094_ _1108_/A vssd1 vssd1 vccd1 vccd1 _1105_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0842__A _0867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1414__46 vssd1 vssd1 vccd1 vccd1 _1414__46/HI _1520_/A sky130_fd_sc_hd__conb_1
X_0947_ _0947_/A vssd1 vssd1 vccd1 vccd1 _0947_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0878_ _0878_/A _0878_/B _0884_/C _0889_/D vssd1 vssd1 vccd1 vccd1 _0879_/A sky130_fd_sc_hd__or4_1
XFILLER_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0801_ _0931_/A vssd1 vssd1 vccd1 vccd1 _0813_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0732_ _1123_/B vssd1 vssd1 vccd1 vccd1 _0847_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1146_ _1155_/A _1140_/X _1144_/X _1145_/X vssd1 vssd1 vccd1 vccd1 _1147_/B sky130_fd_sc_hd__a22o_1
XFILLER_37_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1215_ peripheralBus_data[3] _1538_/A _1228_/S vssd1 vssd1 vccd1 vccd1 _1216_/B sky130_fd_sc_hd__mux2_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1077_ _1077_/A _1077_/B _1085_/C _1085_/D vssd1 vssd1 vccd1 vccd1 _1078_/A sky130_fd_sc_hd__or4_1
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1000_ _1000_/A vssd1 vssd1 vccd1 vccd1 _1000_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1129_ _1542_/A _1128_/A _1541_/A vssd1 vssd1 vccd1 vccd1 _1129_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_33_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput35 _1390_/Q vssd1 vssd1 vccd1 vccd1 spi_mosi[0] sky130_fd_sc_hd__buf_2
XANTENNA__0908__C _0912_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1483__115 vssd1 vssd1 vccd1 vccd1 _1483__115/HI _1613_/A sky130_fd_sc_hd__conb_1
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0910__D _1043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0935__A _0993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0980_ _0994_/A vssd1 vssd1 vccd1 vccd1 _0991_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1532_ _1532_/A _1034_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[29] sky130_fd_sc_hd__ebufn_8
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1601_ _1601_/A _0885_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[2] sky130_fd_sc_hd__ebufn_8
X_1394_ _1396_/CLK _1394_/D vssd1 vssd1 vccd1 vccd1 _1602_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1284__A1 peripheralBus_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1284__B2 _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0963_ _0963_/A _0963_/B _0972_/C _0969_/D vssd1 vssd1 vccd1 vccd1 _0964_/A sky130_fd_sc_hd__or4_1
X_0894_ _0920_/A vssd1 vssd1 vccd1 vccd1 _0904_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1515_ _1515_/A _0984_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[12] sky130_fd_sc_hd__ebufn_8
X_1377_ _1378_/CLK _1377_/D vssd1 vssd1 vccd1 vccd1 _1377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1387__CLK _1396_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1489__121 vssd1 vssd1 vccd1 vccd1 _1489__121/HI _1619_/A sky130_fd_sc_hd__conb_1
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1162_ _1177_/A _1162_/B vssd1 vssd1 vccd1 vccd1 _1163_/A sky130_fd_sc_hd__and2_1
XFILLER_49_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1300_ _1185_/X _1259_/A _1299_/X _1253_/X vssd1 vssd1 vccd1 vccd1 _1301_/B sky130_fd_sc_hd__a22o_1
X_1231_ _1334_/A vssd1 vssd1 vccd1 vccd1 _1348_/A sky130_fd_sc_hd__buf_2
XFILLER_60_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1093_ _1107_/A vssd1 vssd1 vccd1 vccd1 _1105_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0946_ _0948_/A _0948_/B _0958_/C _0946_/D vssd1 vssd1 vccd1 vccd1 _0947_/A sky130_fd_sc_hd__or4_1
X_0877_ _0891_/A vssd1 vssd1 vccd1 vccd1 _0889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1402__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0731_ _1108_/A vssd1 vssd1 vccd1 vccd1 _1123_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_0800_ _1258_/C vssd1 vssd1 vccd1 vccd1 _0931_/A sky130_fd_sc_hd__buf_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1145_ peripheralBus_data[0] vssd1 vssd1 vccd1 vccd1 _1145_/X sky130_fd_sc_hd__clkbuf_4
X_1214_ _1337_/A vssd1 vssd1 vccd1 vccd1 _1269_/A sky130_fd_sc_hd__buf_2
XFILLER_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1076_ _1076_/A vssd1 vssd1 vccd1 vccd1 _1076_/X sky130_fd_sc_hd__clkbuf_1
X_0929_ _0932_/A _0932_/B _0942_/C _0929_/D vssd1 vssd1 vccd1 vccd1 _0930_/A sky130_fd_sc_hd__or4_1
XFILLER_29_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1009__A _1141_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1059_ _1087_/A vssd1 vssd1 vccd1 vccd1 _1071_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1128_ _1128_/A _1128_/B vssd1 vssd1 vccd1 vccd1 _1128_/Y sky130_fd_sc_hd__nand2_2
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput36 _1367_/Q vssd1 vssd1 vccd1 vccd1 spi_mosi[1] sky130_fd_sc_hd__buf_2
X_1465__97 vssd1 vssd1 vccd1 vccd1 _1465__97/HI _1587_/A sky130_fd_sc_hd__conb_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input21_A peripheralBus_address[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0951__A _0994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1531_ _1531_/A _1030_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[28] sky130_fd_sc_hd__ebufn_8
XFILLER_4_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1600_ _1600_/A _0883_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[1] sky130_fd_sc_hd__ebufn_8
X_1393_ _1404_/CLK _1393_/D vssd1 vssd1 vccd1 vccd1 _1601_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1435__67 vssd1 vssd1 vccd1 vccd1 _1435__67/HI _1549_/A sky130_fd_sc_hd__conb_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0962_ _0962_/A vssd1 vssd1 vccd1 vccd1 _0962_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0893_ _0893_/A vssd1 vssd1 vccd1 vccd1 _0893_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1514_ _1514_/A _0978_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[11] sky130_fd_sc_hd__ebufn_8
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1376_ _1378_/CLK _1376_/D vssd1 vssd1 vccd1 vccd1 _1376_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0856__A _0928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1161_ peripheralBus_data[2] _1144_/X _1160_/X _1155_/X vssd1 vssd1 vccd1 vccd1 _1162_/B
+ sky130_fd_sc_hd__a22o_1
X_1092_ _1092_/A vssd1 vssd1 vccd1 vccd1 _1092_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1230_ _1230_/A vssd1 vssd1 vccd1 vccd1 _1375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0945_ _1001_/A vssd1 vssd1 vccd1 vccd1 _0958_/C sky130_fd_sc_hd__buf_2
X_0876_ _0876_/A vssd1 vssd1 vccd1 vccd1 _0876_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1359_ _1378_/CLK _1359_/D vssd1 vssd1 vccd1 vccd1 _1503_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1405__37 vssd1 vssd1 vccd1 vccd1 _1405__37/HI _1511_/A sky130_fd_sc_hd__conb_1
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1210__A _1224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0730_ _1141_/B vssd1 vssd1 vccd1 vccd1 _1108_/A sky130_fd_sc_hd__buf_2
XANTENNA__1166__A1 peripheralBus_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1377__CLK _1378_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1213_ _1213_/A vssd1 vssd1 vccd1 vccd1 _1370_/D sky130_fd_sc_hd__clkbuf_1
X_1144_ _1144_/A vssd1 vssd1 vccd1 vccd1 _1144_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1075_ _1077_/A _1077_/B _1085_/C _1085_/D vssd1 vssd1 vccd1 vccd1 _1076_/A sky130_fd_sc_hd__or4_1
XFILLER_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0859_ _0861_/A _0861_/B _0861_/C _0873_/D vssd1 vssd1 vccd1 vccd1 _0860_/A sky130_fd_sc_hd__or4_1
X_0928_ _0928_/A vssd1 vssd1 vccd1 vccd1 _0942_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1058_ _1058_/A vssd1 vssd1 vccd1 vccd1 _1058_/X sky130_fd_sc_hd__clkbuf_1
X_1127_ _1403_/Q _1402_/Q vssd1 vssd1 vccd1 vccd1 _1128_/B sky130_fd_sc_hd__nor2_2
XFILLER_21_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0949__A _0949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input14_A peripheralBus_address[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 _1367_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1530_ _1530_/A _1028_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[27] sky130_fd_sc_hd__ebufn_8
XANTENNA__1211__A0 peripheralBus_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1392_ _1404_/CLK _1392_/D vssd1 vssd1 vccd1 vccd1 _1600_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A peripheralBus_address[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0961_ _0963_/A _0963_/B _0972_/C _0969_/D vssd1 vssd1 vccd1 vccd1 _0962_/A sky130_fd_sc_hd__or4_1
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1473__105 vssd1 vssd1 vccd1 vccd1 _1473__105/HI _1595_/A sky130_fd_sc_hd__conb_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0892_ _0892_/A _0892_/B _0898_/C _0902_/D vssd1 vssd1 vccd1 vccd1 _0893_/A sky130_fd_sc_hd__or4_1
XFILLER_4_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1375_ _1404_/CLK _1375_/D vssd1 vssd1 vccd1 vccd1 _1542_/A sky130_fd_sc_hd__dfxtp_1
X_1513_ _1513_/A _0976_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[10] sky130_fd_sc_hd__ebufn_8
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1160_ _1505_/A _1159_/X _1175_/S vssd1 vssd1 vccd1 vccd1 _1160_/X sky130_fd_sc_hd__mux2_1
X_1091_ _1091_/A _1091_/B _1099_/C _1099_/D vssd1 vssd1 vccd1 vccd1 _1092_/A sky130_fd_sc_hd__or4_1
XFILLER_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0944_ _1258_/B vssd1 vssd1 vccd1 vccd1 _1001_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0875_ _0878_/A _0878_/B _0912_/C _0915_/D vssd1 vssd1 vccd1 vccd1 _0876_/A sky130_fd_sc_hd__or4_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0867__A _0867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1358_ _1354_/Y _1357_/Y _1147_/A vssd1 vssd1 vccd1 vccd1 _1404_/D sky130_fd_sc_hd__o21a_1
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1289_ peripheralBus_data[5] _1259_/A _1288_/X _1253_/X vssd1 vssd1 vccd1 vccd1 _1290_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1212_ _1222_/A _1212_/B vssd1 vssd1 vccd1 vccd1 _1213_/A sky130_fd_sc_hd__or2_1
XFILLER_1_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1074_ _1088_/A vssd1 vssd1 vccd1 vccd1 _1085_/D sky130_fd_sc_hd__clkbuf_1
X_1143_ _1143_/A _1258_/B _1143_/C _1353_/C vssd1 vssd1 vccd1 vccd1 _1144_/A sky130_fd_sc_hd__nor4_4
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0927_ _0927_/A vssd1 vssd1 vccd1 vccd1 _0927_/X sky130_fd_sc_hd__clkbuf_1
X_1479__111 vssd1 vssd1 vccd1 vccd1 _1479__111/HI _1609_/A sky130_fd_sc_hd__conb_1
X_0858_ _0858_/A vssd1 vssd1 vccd1 vccd1 _0858_/X sky130_fd_sc_hd__clkbuf_1
X_0789_ _0793_/A _0793_/B _0789_/C _0818_/D vssd1 vssd1 vccd1 vccd1 _0790_/A sky130_fd_sc_hd__or4_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1126_ _1250_/B _1379_/Q vssd1 vssd1 vccd1 vccd1 _1128_/A sky130_fd_sc_hd__nor2_2
X_1057_ _1063_/A _1063_/B _1057_/C _1057_/D vssd1 vssd1 vccd1 vccd1 _1058_/A sky130_fd_sc_hd__or4_1
XFILLER_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1216__A _1269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0965__A _0993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
X_1456__88 vssd1 vssd1 vccd1 vccd1 _1456__88/HI _1578_/A sky130_fd_sc_hd__conb_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1109_ _1117_/A _1117_/B _1113_/C _1113_/D vssd1 vssd1 vccd1 vccd1 _1110_/A sky130_fd_sc_hd__or4_1
XFILLER_26_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1391_ _1404_/CLK _1391_/D vssd1 vssd1 vccd1 vccd1 _1599_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1589_ _1589_/A _0807_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[22] sky130_fd_sc_hd__ebufn_8
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0946__C _0958_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1426__58 vssd1 vssd1 vccd1 vccd1 _1426__58/HI _1532_/A sky130_fd_sc_hd__conb_1
XFILLER_43_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0960_ _1001_/A vssd1 vssd1 vccd1 vccd1 _0972_/C sky130_fd_sc_hd__buf_2
XANTENNA__1196__A0 _1145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1512_ _1512_/A _0973_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[9] sky130_fd_sc_hd__ebufn_8
X_0891_ _0891_/A vssd1 vssd1 vccd1 vccd1 _0902_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1374_ _1378_/CLK _1374_/D vssd1 vssd1 vccd1 vccd1 _1541_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1440__72 vssd1 vssd1 vccd1 vccd1 _1440__72/HI _1554_/A sky130_fd_sc_hd__conb_1
XANTENNA__1187__A0 _1510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 _1378_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1224__A _1224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1496__128 vssd1 vssd1 vccd1 vccd1 _1496__128/HI _1626_/A sky130_fd_sc_hd__conb_1
XFILLER_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1090_ _1090_/A vssd1 vssd1 vccd1 vccd1 _1090_/X sky130_fd_sc_hd__clkbuf_1
X_0943_ _0943_/A vssd1 vssd1 vccd1 vccd1 _0943_/X sky130_fd_sc_hd__clkbuf_1
X_0874_ _0874_/A vssd1 vssd1 vccd1 vccd1 _0874_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1357_ _1357_/A _1357_/B vssd1 vssd1 vccd1 vccd1 _1357_/Y sky130_fd_sc_hd__nor2_1
X_1288_ _1572_/A _1287_/X _1288_/S vssd1 vssd1 vccd1 vccd1 _1288_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1219__A _1269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1211_ peripheralBus_data[2] _1537_/A _1225_/S vssd1 vssd1 vccd1 vccd1 _1212_/B sky130_fd_sc_hd__mux2_1
XFILLER_27_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1142_ _1313_/C vssd1 vssd1 vccd1 vccd1 _1353_/C sky130_fd_sc_hd__buf_2
XFILLER_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1073_ _1087_/A vssd1 vssd1 vccd1 vccd1 _1085_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_1_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0857_ _0861_/A _0861_/B _0912_/C _0857_/D vssd1 vssd1 vccd1 vccd1 _0858_/A sky130_fd_sc_hd__or4_1
X_0926_ _0932_/A _0932_/B _0926_/C _0929_/D vssd1 vssd1 vccd1 vccd1 _0927_/A sky130_fd_sc_hd__or4_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0788_ _0788_/A vssd1 vssd1 vccd1 vccd1 _0788_/X sky130_fd_sc_hd__clkbuf_1
X_1410__42 vssd1 vssd1 vccd1 vccd1 _1410__42/HI _1516_/A sky130_fd_sc_hd__conb_1
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0954__C _0958_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1125_ _1380_/Q vssd1 vssd1 vccd1 vccd1 _1250_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1056_ _1056_/A vssd1 vssd1 vccd1 vccd1 _1056_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0909_ _0909_/A vssd1 vssd1 vccd1 vccd1 _0909_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1108_ _1108_/A vssd1 vssd1 vccd1 vccd1 _1117_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_38_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1039_ _1049_/A _1049_/B _1123_/C _1043_/D vssd1 vssd1 vccd1 vccd1 _1040_/A sky130_fd_sc_hd__or4_1
XANTENNA__1052__A _1066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0891__A _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1390_ _1396_/CLK _1390_/D vssd1 vssd1 vccd1 vccd1 _1390_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__0861__D _0873_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1588_ _1588_/A _0805_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[21] sky130_fd_sc_hd__ebufn_8
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0886__A _1258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1510__A _1510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0890_ _0890_/A vssd1 vssd1 vccd1 vccd1 _0890_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1196__A1 _1185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1511_ _1511_/A _0970_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[8] sky130_fd_sc_hd__ebufn_8
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1373_ _1378_/CLK _1373_/D vssd1 vssd1 vccd1 vccd1 _1540_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1150__A _1337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0942_ _0948_/A _0948_/B _0942_/C _0946_/D vssd1 vssd1 vccd1 vccd1 _0943_/A sky130_fd_sc_hd__or4_1
X_0873_ _0878_/A _0878_/B _0884_/C _0873_/D vssd1 vssd1 vccd1 vccd1 _0874_/A sky130_fd_sc_hd__or4_1
XFILLER_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1287_ _1573_/A _1571_/A _1298_/S vssd1 vssd1 vccd1 vccd1 _1287_/X sky130_fd_sc_hd__mux2_1
X_1356_ _1357_/B _1343_/C _1128_/B _1222_/A vssd1 vssd1 vccd1 vccd1 _1403_/D sky130_fd_sc_hd__a211oi_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1145__A peripheralBus_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1072_ _1072_/A vssd1 vssd1 vccd1 vccd1 _1072_/X sky130_fd_sc_hd__clkbuf_1
X_1141_ _1141_/A _1141_/B vssd1 vssd1 vccd1 vccd1 _1313_/C sky130_fd_sc_hd__nand2_1
X_1210_ _1224_/A vssd1 vssd1 vccd1 vccd1 _1222_/A sky130_fd_sc_hd__buf_2
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_clk clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 _1404_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_18_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0787_ _0793_/A _0793_/B _0789_/C _0818_/D vssd1 vssd1 vccd1 vccd1 _0788_/A sky130_fd_sc_hd__or4_1
X_0925_ _0925_/A vssd1 vssd1 vccd1 vccd1 _0925_/X sky130_fd_sc_hd__clkbuf_1
X_0856_ _0928_/A vssd1 vssd1 vccd1 vccd1 _0912_/C sky130_fd_sc_hd__buf_2
X_1339_ _1403_/Q vssd1 vssd1 vccd1 vccd1 _1357_/B sky130_fd_sc_hd__inv_2
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0954__D _0954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0979__A _0993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1390__CLK _1396_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1025__D _1029_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1124_ _1124_/A vssd1 vssd1 vccd1 vccd1 _1124_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1041__C _1043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1055_ _1063_/A _1063_/B _1057_/C _1057_/D vssd1 vssd1 vccd1 vccd1 _1056_/A sky130_fd_sc_hd__or4_1
XFILLER_25_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0839_ _0839_/A vssd1 vssd1 vccd1 vccd1 _0839_/X sky130_fd_sc_hd__clkbuf_1
X_0908_ _0918_/A _0918_/B _0912_/C _0915_/D vssd1 vssd1 vccd1 vccd1 _0909_/A sky130_fd_sc_hd__or4_1
XFILLER_56_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1469__101 vssd1 vssd1 vccd1 vccd1 _1469__101/HI _1591_/A sky130_fd_sc_hd__conb_1
XFILLER_30_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0859__D _0873_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0875__C _0912_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1447__79 vssd1 vssd1 vccd1 vccd1 _1447__79/HI _1561_/A sky130_fd_sc_hd__conb_1
X_1107_ _1107_/A vssd1 vssd1 vccd1 vccd1 _1117_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_42_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1038_ _1066_/A vssd1 vssd1 vccd1 vccd1 _1049_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_26_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1461__93 vssd1 vssd1 vccd1 vccd1 _1461__93/HI _1583_/A sky130_fd_sc_hd__conb_1
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1587_ _1587_/A _0803_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[20] sky130_fd_sc_hd__ebufn_8
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1328__A _1337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input12_A peripheralBus_address[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1510_ _1510_/A _0968_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[7] sky130_fd_sc_hd__ebufn_8
XFILLER_4_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1372_ _1378_/CLK _1372_/D vssd1 vssd1 vccd1 vccd1 _1539_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1417__49 vssd1 vssd1 vccd1 vccd1 _1417__49/HI _1523_/A sky130_fd_sc_hd__conb_1
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input4_A peripheralBus_address[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1431__63 vssd1 vssd1 vccd1 vccd1 _1431__63/HI _1545_/A sky130_fd_sc_hd__conb_1
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0941_ _0941_/A vssd1 vssd1 vccd1 vccd1 _0941_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0872_ _0872_/A vssd1 vssd1 vccd1 vccd1 _0872_/X sky130_fd_sc_hd__clkbuf_1
X_1355_ _1352_/X _1354_/Y _1147_/A vssd1 vssd1 vccd1 vccd1 _1402_/D sky130_fd_sc_hd__o21a_1
XFILLER_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1286_ _1286_/A vssd1 vssd1 vccd1 vccd1 _1386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1140_ _1503_/A _1138_/X _1193_/S vssd1 vssd1 vccd1 vccd1 _1140_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1071_ _1077_/A _1077_/B _1071_/C _1071_/D vssd1 vssd1 vccd1 vccd1 _1072_/A sky130_fd_sc_hd__or4_1
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0924_ _0932_/A _0932_/B _0926_/C _0929_/D vssd1 vssd1 vccd1 vccd1 _0925_/A sky130_fd_sc_hd__or4_1
X_0855_ _0855_/A vssd1 vssd1 vccd1 vccd1 _0855_/X sky130_fd_sc_hd__clkbuf_1
X_0786_ _0786_/A vssd1 vssd1 vccd1 vccd1 _0786_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1486__118 vssd1 vssd1 vccd1 vccd1 _1486__118/HI _1616_/A sky130_fd_sc_hd__conb_1
XFILLER_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1338_ _1338_/A vssd1 vssd1 vccd1 vccd1 _1398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1269_ _1269_/A _1269_/B vssd1 vssd1 vccd1 vccd1 _1270_/A sky130_fd_sc_hd__and2_1
XFILLER_3_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1123_ _1123_/A _1123_/B _1123_/C _1123_/D vssd1 vssd1 vccd1 vccd1 _1124_/A sky130_fd_sc_hd__or4_1
XFILLER_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1054_ _1054_/A vssd1 vssd1 vccd1 vccd1 _1054_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0907_ _0921_/A vssd1 vssd1 vccd1 vccd1 _0918_/B sky130_fd_sc_hd__clkbuf_1
X_0838_ _0845_/A _0845_/B _0840_/C _0845_/D vssd1 vssd1 vccd1 vccd1 _0839_/A sky130_fd_sc_hd__or4_1
X_0769_ _0769_/A vssd1 vssd1 vccd1 vccd1 _0769_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1066__A _1066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_clk clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 _1396_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_47_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1106_ _1106_/A vssd1 vssd1 vccd1 vccd1 _1106_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1037_ _1065_/A vssd1 vssd1 vccd1 vccd1 _1049_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1380__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1586_ _1586_/A _0794_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[19] sky130_fd_sc_hd__ebufn_8
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1371_ _1378_/CLK _1371_/D vssd1 vssd1 vccd1 vccd1 _1538_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ _1569_/A _0916_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[2] sky130_fd_sc_hd__ebufn_8
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0940_ _0948_/A _0948_/B _0942_/C _0946_/D vssd1 vssd1 vccd1 vccd1 _0941_/A sky130_fd_sc_hd__or4_1
XFILLER_9_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0871_ _0878_/A _0878_/B _0912_/C _0915_/D vssd1 vssd1 vccd1 vccd1 _0872_/A sky130_fd_sc_hd__or4_1
X_1285_ _1295_/A _1285_/B vssd1 vssd1 vccd1 vccd1 _1286_/A sky130_fd_sc_hd__and2_1
X_1354_ _1403_/Q _1402_/Q _1354_/C vssd1 vssd1 vccd1 vccd1 _1354_/Y sky130_fd_sc_hd__nor3_1
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0793__D _0793_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1308__A0 peripheralBus_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1070_ _1070_/A vssd1 vssd1 vccd1 vccd1 _1070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0854_ _0861_/A _0861_/B _0854_/C _0857_/D vssd1 vssd1 vccd1 vccd1 _0855_/A sky130_fd_sc_hd__or4_1
XANTENNA__1244__C1 _1147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0923_ _0923_/A vssd1 vssd1 vccd1 vccd1 _0923_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0785_ _0793_/A _0793_/B _0789_/C _0818_/D vssd1 vssd1 vccd1 vccd1 _0786_/A sky130_fd_sc_hd__or4_1
X_1268_ peripheralBus_data[1] _1259_/X _1266_/X _1357_/A vssd1 vssd1 vccd1 vccd1 _1269_/B
+ sky130_fd_sc_hd__a22o_1
X_1337_ _1337_/A _1337_/B vssd1 vssd1 vccd1 vccd1 _1338_/A sky130_fd_sc_hd__and2_1
X_1199_ _1199_/A vssd1 vssd1 vccd1 vccd1 _1367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1122_ _1122_/A vssd1 vssd1 vccd1 vccd1 _1122_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1053_ _1063_/A _1063_/B _1057_/C _1057_/D vssd1 vssd1 vccd1 vccd1 _1054_/A sky130_fd_sc_hd__or4_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0837_ _0837_/A vssd1 vssd1 vccd1 vccd1 _0837_/X sky130_fd_sc_hd__clkbuf_1
X_0906_ _0920_/A vssd1 vssd1 vccd1 vccd1 _0918_/A sky130_fd_sc_hd__clkbuf_1
X_0768_ _0775_/A _0775_/B _1123_/D _0775_/D vssd1 vssd1 vccd1 vccd1 _0769_/A sky130_fd_sc_hd__or4_1
XFILLER_56_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1105_ _1105_/A _1105_/B _1113_/C _1113_/D vssd1 vssd1 vccd1 vccd1 _1106_/A sky130_fd_sc_hd__or4_1
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1036_ _1036_/A vssd1 vssd1 vccd1 vccd1 _1036_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1452__84 vssd1 vssd1 vccd1 vccd1 _1452__84/HI _1566_/A sky130_fd_sc_hd__conb_1
XFILLER_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1585_ _1585_/A _0782_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[18] sky130_fd_sc_hd__ebufn_8
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1019_ _1021_/A _1021_/B _1029_/C _1029_/D vssd1 vssd1 vccd1 vccd1 _1020_/A sky130_fd_sc_hd__or4_1
XFILLER_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1370_ _1378_/CLK _1370_/D vssd1 vssd1 vccd1 vccd1 _1537_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1370__CLK _1378_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ _1568_/A _0913_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[1] sky130_fd_sc_hd__ebufn_8
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0870_ _0931_/A vssd1 vssd1 vccd1 vccd1 _0915_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_1422__54 vssd1 vssd1 vccd1 vccd1 _1422__54/HI _1528_/A sky130_fd_sc_hd__conb_1
XANTENNA__1393__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1353_ _1353_/A _1353_/B _1353_/C _1353_/D vssd1 vssd1 vccd1 vccd1 _1354_/C sky130_fd_sc_hd__or4_2
X_1284_ peripheralBus_data[4] _1259_/A _1283_/X _1357_/A vssd1 vssd1 vccd1 vccd1 _1285_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0999_ _1005_/A _1005_/B _0999_/C _0999_/D vssd1 vssd1 vccd1 vccd1 _1000_/A sky130_fd_sc_hd__or4_1
XFILLER_27_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1308__A1 peripheralBus_data[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0853_ _0853_/A vssd1 vssd1 vccd1 vccd1 _0853_/X sky130_fd_sc_hd__clkbuf_2
X_0922_ _0932_/A _0932_/B _0926_/C _0929_/D vssd1 vssd1 vccd1 vccd1 _0923_/A sky130_fd_sc_hd__or4_1
X_0784_ _0891_/A vssd1 vssd1 vccd1 vccd1 _0818_/D sky130_fd_sc_hd__clkbuf_2
X_1198_ _1208_/A _1198_/B vssd1 vssd1 vccd1 vccd1 _1199_/A sky130_fd_sc_hd__and2_1
Xinput1 peripheralBus_address[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
X_1267_ _1267_/A vssd1 vssd1 vccd1 vccd1 _1357_/A sky130_fd_sc_hd__clkbuf_4
X_1336_ _1185_/X _1606_/A _1336_/S vssd1 vssd1 vccd1 vccd1 _1337_/B sky130_fd_sc_hd__mux2_1
XFILLER_51_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1121_ _1123_/A _1123_/B _1121_/C _1121_/D vssd1 vssd1 vccd1 vccd1 _1122_/A sky130_fd_sc_hd__or4_1
X_1052_ _1066_/A vssd1 vssd1 vccd1 vccd1 _1063_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_25_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1492__124 vssd1 vssd1 vccd1 vccd1 _1492__124/HI _1622_/A sky130_fd_sc_hd__conb_1
X_0836_ _0847_/A _0847_/B _1043_/C _0954_/D vssd1 vssd1 vccd1 vccd1 _0837_/A sky130_fd_sc_hd__or4_1
X_0767_ _0767_/A vssd1 vssd1 vccd1 vccd1 _0767_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0905_ _0905_/A vssd1 vssd1 vccd1 vccd1 _0905_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1319_ _1325_/A _1319_/B vssd1 vssd1 vccd1 vccd1 _1320_/A sky130_fd_sc_hd__and2_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1458__90 vssd1 vssd1 vccd1 vccd1 _1458__90/HI _1580_/A sky130_fd_sc_hd__conb_1
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input28_A spi_miso[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1476__108 vssd1 vssd1 vccd1 vccd1 _1476__108/HI _1598_/A sky130_fd_sc_hd__conb_1
XFILLER_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1104_ _1104_/A vssd1 vssd1 vccd1 vccd1 _1104_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1035_ _1035_/A _1035_/B _1123_/C _1043_/D vssd1 vssd1 vccd1 vccd1 _1036_/A sky130_fd_sc_hd__or4_1
XFILLER_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0819_ _0819_/A vssd1 vssd1 vccd1 vccd1 _0819_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1584_ _1584_/A _0774_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[17] sky130_fd_sc_hd__ebufn_8
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1018_ _1018_/A vssd1 vssd1 vccd1 vccd1 _1029_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1428__60 vssd1 vssd1 vccd1 vccd1 _1428__60/HI _1534_/A sky130_fd_sc_hd__conb_1
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1498__130 vssd1 vssd1 vccd1 vccd1 _1498__130/HI _1628_/A sky130_fd_sc_hd__conb_1
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1567_ _1567_/A _0909_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[0] sky130_fd_sc_hd__ebufn_8
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input10_A peripheralBus_address[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1283_ _1571_/A _1282_/X _1288_/S vssd1 vssd1 vccd1 vccd1 _1283_/X sky130_fd_sc_hd__mux2_1
X_1352_ _1403_/Q _1343_/C _1402_/Q vssd1 vssd1 vccd1 vccd1 _1352_/X sky130_fd_sc_hd__o21a_1
X_0998_ _0998_/A vssd1 vssd1 vccd1 vccd1 _0998_/X sky130_fd_sc_hd__clkbuf_1
X_1619_ _1619_/A _0819_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[20] sky130_fd_sc_hd__ebufn_8
XFILLER_59_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input2_A peripheralBus_address[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0921_ _0921_/A vssd1 vssd1 vccd1 vccd1 _0932_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_0852_ _0861_/A _0861_/B _0861_/C _0873_/D vssd1 vssd1 vccd1 vccd1 _0853_/A sky130_fd_sc_hd__or4_1
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0783_ _1202_/B vssd1 vssd1 vccd1 vccd1 _0891_/A sky130_fd_sc_hd__buf_2
XANTENNA__1180__A0 _1510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1404_ _1404_/CLK _1404_/D vssd1 vssd1 vccd1 vccd1 _1404_/Q sky130_fd_sc_hd__dfxtp_1
X_1335_ _1335_/A vssd1 vssd1 vccd1 vccd1 _1397_/D sky130_fd_sc_hd__clkbuf_1
X_1197_ _1155_/A _1195_/X _1196_/X _1144_/X vssd1 vssd1 vccd1 vccd1 _1198_/B sky130_fd_sc_hd__a22o_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 peripheralBus_address[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
X_1266_ _1568_/A _1264_/X _1288_/S vssd1 vssd1 vccd1 vccd1 _1266_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1383__CLK _1396_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1120_ _1120_/A vssd1 vssd1 vccd1 vccd1 _1120_/X sky130_fd_sc_hd__clkbuf_1
X_1051_ _1065_/A vssd1 vssd1 vccd1 vccd1 _1063_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0904_ _0904_/A _0904_/B _0910_/C _1043_/C vssd1 vssd1 vccd1 vccd1 _0905_/A sky130_fd_sc_hd__or4_1
X_0835_ _1121_/D vssd1 vssd1 vccd1 vccd1 _0954_/D sky130_fd_sc_hd__clkbuf_2
X_0766_ _0775_/A _0775_/B _1123_/D _0775_/D vssd1 vssd1 vccd1 vccd1 _0767_/A sky130_fd_sc_hd__or4_1
X_1318_ peripheralBus_data[1] _1600_/A _1336_/S vssd1 vssd1 vccd1 vccd1 _1319_/B sky130_fd_sc_hd__mux2_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1249_ _1236_/A _1236_/C _1128_/A _1222_/A vssd1 vssd1 vccd1 vccd1 _1380_/D sky130_fd_sc_hd__a211oi_1
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1103_ _1105_/A _1105_/B _1113_/C _1113_/D vssd1 vssd1 vccd1 vccd1 _1104_/A sky130_fd_sc_hd__or4_1
XFILLER_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1034_ _1034_/A vssd1 vssd1 vccd1 vccd1 _1034_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1500__132 vssd1 vssd1 vccd1 vccd1 _1500__132/HI _1630_/A sky130_fd_sc_hd__conb_1
X_0818_ _0823_/A _0823_/B _0840_/C _0818_/D vssd1 vssd1 vccd1 vccd1 _0819_/A sky130_fd_sc_hd__or4_1
X_0749_ _0749_/A vssd1 vssd1 vccd1 vccd1 _0749_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1583_ _1583_/A _0763_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[16] sky130_fd_sc_hd__ebufn_8
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1017_ _1353_/B vssd1 vssd1 vccd1 vccd1 _1029_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_34_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1443__75 vssd1 vssd1 vccd1 vccd1 _1443__75/HI _1557_/A sky130_fd_sc_hd__conb_1
XFILLER_57_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1566_ _1566_/A _1120_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[31] sky130_fd_sc_hd__ebufn_8
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1351_ _1401_/Q _1343_/X _1350_/Y _1147_/A vssd1 vssd1 vccd1 vccd1 _1401_/D sky130_fd_sc_hd__o211a_1
X_1282_ _1572_/A _1570_/A _1298_/S vssd1 vssd1 vccd1 vccd1 _1282_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1618_ _1618_/A _0799_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[19] sky130_fd_sc_hd__ebufn_8
X_0997_ _1005_/A _1005_/B _0999_/C _0999_/D vssd1 vssd1 vccd1 vccd1 _0998_/A sky130_fd_sc_hd__or4_1
X_1413__45 vssd1 vssd1 vccd1 vccd1 _1413__45/HI _1519_/A sky130_fd_sc_hd__conb_1
X_1549_ _1549_/A _1076_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[14] sky130_fd_sc_hd__ebufn_8
XANTENNA__0726__A _1141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0920_ _0920_/A vssd1 vssd1 vccd1 vccd1 _0932_/A sky130_fd_sc_hd__clkbuf_1
X_0851_ _0891_/A vssd1 vssd1 vccd1 vccd1 _0873_/D sky130_fd_sc_hd__clkbuf_2
X_0782_ _0782_/A vssd1 vssd1 vccd1 vccd1 _0782_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1265_ _1305_/S vssd1 vssd1 vccd1 vccd1 _1288_/S sky130_fd_sc_hd__clkbuf_2
X_1403_ _1404_/CLK _1403_/D vssd1 vssd1 vccd1 vccd1 _1403_/Q sky130_fd_sc_hd__dfxtp_1
X_1334_ _1334_/A _1334_/B vssd1 vssd1 vccd1 vccd1 _1335_/A sky130_fd_sc_hd__or2_1
X_1196_ _1145_/X _1185_/X _1196_/S vssd1 vssd1 vccd1 vccd1 _1196_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput3 peripheralBus_address[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1171__A1 peripheralBus_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output34_A _1130_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1050_ _1050_/A vssd1 vssd1 vccd1 vccd1 _1050_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0834_ _1143_/C vssd1 vssd1 vccd1 vccd1 _1121_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0903_ _0903_/A vssd1 vssd1 vccd1 vccd1 _0903_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0765_ _1123_/B vssd1 vssd1 vccd1 vccd1 _0775_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1317_ _1317_/A vssd1 vssd1 vccd1 vccd1 _1391_/D sky130_fd_sc_hd__clkbuf_1
X_1248_ _1245_/Y _1247_/X _1348_/A vssd1 vssd1 vccd1 vccd1 _1379_/D sky130_fd_sc_hd__a21oi_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1179_ _1337_/A vssd1 vssd1 vccd1 vccd1 _1208_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1449__81 vssd1 vssd1 vccd1 vccd1 _1449__81/HI _1563_/A sky130_fd_sc_hd__conb_1
XFILLER_62_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0914__A _0928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1102_ _1143_/C vssd1 vssd1 vccd1 vccd1 _1113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1033_ _1035_/A _1035_/B _1123_/C _1043_/D vssd1 vssd1 vccd1 vccd1 _1034_/A sky130_fd_sc_hd__or4_1
X_0817_ _0817_/A vssd1 vssd1 vccd1 vccd1 _0817_/X sky130_fd_sc_hd__clkbuf_1
X_0748_ _0847_/A _0847_/B _0847_/C _0793_/D vssd1 vssd1 vccd1 vccd1 _0749_/A sky130_fd_sc_hd__or4_1
XANTENNA__1373__CLK _1378_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1482__114 vssd1 vssd1 vccd1 vccd1 _1482__114/HI _1612_/A sky130_fd_sc_hd__conb_1
XFILLER_7_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1582_ _1582_/A _0749_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[15] sky130_fd_sc_hd__ebufn_8
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1396__CLK _1396_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1016_ _1016_/A vssd1 vssd1 vccd1 vccd1 _1016_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1419__51 vssd1 vssd1 vccd1 vccd1 _1419__51/HI _1525_/A sky130_fd_sc_hd__conb_1
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1295__A _1295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1565_ _1565_/A _1118_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[30] sky130_fd_sc_hd__ebufn_8
XFILLER_39_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1488__120 vssd1 vssd1 vccd1 vccd1 _1488__120/HI _1618_/A sky130_fd_sc_hd__conb_1
X_1281_ _1281_/A vssd1 vssd1 vccd1 vccd1 _1385_/D sky130_fd_sc_hd__clkbuf_1
X_1350_ _1401_/Q _1349_/Y _1343_/X vssd1 vssd1 vccd1 vccd1 _1350_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0996_ _0996_/A vssd1 vssd1 vccd1 vccd1 _0996_/X sky130_fd_sc_hd__clkbuf_1
X_1617_ _1617_/A _0790_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[18] sky130_fd_sc_hd__ebufn_8
XFILLER_8_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1548_ _1548_/A _1072_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[13] sky130_fd_sc_hd__ebufn_8
XFILLER_6_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0917__A _0931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0850_ _0850_/A vssd1 vssd1 vccd1 vccd1 _0861_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0781_ _0793_/A _0793_/B _0847_/C _0793_/D vssd1 vssd1 vccd1 vccd1 _0782_/A sky130_fd_sc_hd__or4_1
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1402_ _1404_/CLK _1402_/D vssd1 vssd1 vccd1 vccd1 _1402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput4 peripheralBus_address[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
X_1264_ _1569_/A _1567_/A _1308_/S vssd1 vssd1 vccd1 vccd1 _1264_/X sky130_fd_sc_hd__mux2_1
X_1333_ peripheralBus_data[6] _1605_/A _1333_/S vssd1 vssd1 vccd1 vccd1 _1334_/B sky130_fd_sc_hd__mux2_1
XFILLER_51_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1195_ _1367_/Q _1193_/X _1195_/S vssd1 vssd1 vccd1 vccd1 _1195_/X sky130_fd_sc_hd__mux2_1
X_0979_ _0993_/A vssd1 vssd1 vccd1 vccd1 _0991_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1171__A2 _1144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0833_ _1246_/A _1312_/B _1312_/C _0833_/D vssd1 vssd1 vccd1 vccd1 _1143_/C sky130_fd_sc_hd__or4_4
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0902_ _0904_/A _0904_/B _0910_/C _0902_/D vssd1 vssd1 vccd1 vccd1 _0903_/A sky130_fd_sc_hd__or4_1
X_0764_ _1123_/A vssd1 vssd1 vccd1 vccd1 _0775_/A sky130_fd_sc_hd__clkbuf_1
X_1178_ _1178_/A vssd1 vssd1 vccd1 vccd1 _1364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1247_ _1250_/B _1379_/Q _1247_/C vssd1 vssd1 vccd1 vccd1 _1247_/X sky130_fd_sc_hd__or3_1
X_1316_ _1325_/A _1316_/B vssd1 vssd1 vccd1 vccd1 _1317_/A sky130_fd_sc_hd__and2_1
XFILLER_64_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1464__96 vssd1 vssd1 vccd1 vccd1 _1464__96/HI _1586_/A sky130_fd_sc_hd__conb_1
XFILLER_11_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1101_ _1202_/B vssd1 vssd1 vccd1 vccd1 _1113_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1032_ _1088_/A vssd1 vssd1 vccd1 vccd1 _1043_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0816_ _0823_/A _0823_/B _0854_/C _0857_/D vssd1 vssd1 vccd1 vccd1 _0817_/A sky130_fd_sc_hd__or4_1
X_0747_ _0910_/C vssd1 vssd1 vccd1 vccd1 _0793_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_37_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0750__A _1258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input26_A peripheralBus_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1581_ _1581_/A _1124_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[14] sky130_fd_sc_hd__ebufn_8
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1015_ _1021_/A _1021_/B _1015_/C _1015_/D vssd1 vssd1 vccd1 vccd1 _1016_/A sky130_fd_sc_hd__or4_1
XFILLER_22_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1434__66 vssd1 vssd1 vccd1 vccd1 _1434__66/HI _1548_/A sky130_fd_sc_hd__conb_1
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1274__B2 _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1274__A1 peripheralBus_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1564_ _1564_/A _1116_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[29] sky130_fd_sc_hd__ebufn_8
XFILLER_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1386__CLK _1396_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1280_ _1295_/A _1280_/B vssd1 vssd1 vccd1 vccd1 _1281_/A sky130_fd_sc_hd__and2_1
XFILLER_63_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0995_ _1005_/A _1005_/B _0999_/C _0999_/D vssd1 vssd1 vccd1 vccd1 _0996_/A sky130_fd_sc_hd__or4_1
X_1616_ _1616_/A _0788_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[17] sky130_fd_sc_hd__ebufn_8
X_1547_ _1547_/A _1070_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[12] sky130_fd_sc_hd__ebufn_8
XFILLER_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0780_ _0850_/A vssd1 vssd1 vccd1 vccd1 _0793_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1401_ _1404_/CLK _1401_/D vssd1 vssd1 vccd1 vccd1 _1401_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1401__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 peripheralBus_address[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
X_1194_ _1376_/Q _1377_/Q _1538_/A vssd1 vssd1 vccd1 vccd1 _1195_/S sky130_fd_sc_hd__mux2_1
X_1263_ _1604_/A vssd1 vssd1 vccd1 vccd1 _1308_/S sky130_fd_sc_hd__buf_2
X_1332_ _1332_/A vssd1 vssd1 vccd1 vccd1 _1396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0978_ _0978_/A vssd1 vssd1 vccd1 vccd1 _0978_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0928__A _0928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0763_ _0763_/A vssd1 vssd1 vccd1 vccd1 _0763_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0832_ input4/X input7/X input6/X vssd1 vssd1 vccd1 vccd1 _0833_/D sky130_fd_sc_hd__or3_1
X_0901_ _0901_/A vssd1 vssd1 vccd1 vccd1 _0901_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1315_ _1145_/X _1599_/A _1336_/S vssd1 vssd1 vccd1 vccd1 _1316_/B sky130_fd_sc_hd__mux2_1
X_1177_ _1177_/A _1177_/B vssd1 vssd1 vccd1 vccd1 _1178_/A sky130_fd_sc_hd__and2_1
XFILLER_56_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1246_ _1246_/A _1353_/B _1353_/C _1246_/D vssd1 vssd1 vccd1 vccd1 _1247_/C sky130_fd_sc_hd__or4_2
XFILLER_2_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1100_ _1100_/A vssd1 vssd1 vccd1 vccd1 _1100_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1031_ _1143_/C vssd1 vssd1 vccd1 vccd1 _1088_/A sky130_fd_sc_hd__clkbuf_2
X_0815_ _0931_/A vssd1 vssd1 vccd1 vccd1 _0857_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_0746_ _1258_/C vssd1 vssd1 vccd1 vccd1 _0910_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1229_ _1269_/A _1229_/B vssd1 vssd1 vccd1 vccd1 _1230_/A sky130_fd_sc_hd__and2_1
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input19_A peripheralBus_address[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1102__A _1143_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1580_ _1580_/A _0982_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[13] sky130_fd_sc_hd__ebufn_8
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1014_ _1014_/A vssd1 vssd1 vccd1 vccd1 _1014_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0851__A _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0729_ _0729_/A vssd1 vssd1 vccd1 vccd1 _1141_/B sky130_fd_sc_hd__inv_2
XFILLER_57_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0936__A _1141_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1563_ _1563_/A _1114_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[28] sky130_fd_sc_hd__ebufn_8
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1007__A _1141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1472__104 vssd1 vssd1 vccd1 vccd1 _1472__104/HI _1594_/A sky130_fd_sc_hd__conb_1
XFILLER_13_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0994_ _0994_/A vssd1 vssd1 vccd1 vccd1 _1005_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1615_ _1615_/A _0786_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[16] sky130_fd_sc_hd__ebufn_8
X_1546_ _1546_/A _1068_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[11] sky130_fd_sc_hd__ebufn_8
XFILLER_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1400_ _1404_/CLK _1400_/D vssd1 vssd1 vccd1 vccd1 _1400_/Q sky130_fd_sc_hd__dfxtp_1
X_1331_ _1334_/A _1331_/B vssd1 vssd1 vccd1 vccd1 _1332_/A sky130_fd_sc_hd__or2_1
X_1193_ _1191_/X _1192_/X _1193_/S vssd1 vssd1 vccd1 vccd1 _1193_/X sky130_fd_sc_hd__mux2_1
Xinput6 peripheralBus_address[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
X_1262_ _1262_/A vssd1 vssd1 vccd1 vccd1 _1382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1376__CLK _1378_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0977_ _0977_/A _0977_/B _0985_/C _0985_/D vssd1 vssd1 vccd1 vccd1 _0978_/A sky130_fd_sc_hd__or4_1
X_1529_ _1529_/A _1026_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[26] sky130_fd_sc_hd__ebufn_8
XANTENNA__1156__A1 peripheralBus_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1478__110 vssd1 vssd1 vccd1 vccd1 _1478__110/HI _1608_/A sky130_fd_sc_hd__conb_1
XFILLER_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0944__A _1258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0900_ _0904_/A _0904_/B _0910_/C _0902_/D vssd1 vssd1 vccd1 vccd1 _0901_/A sky130_fd_sc_hd__or4_1
X_0762_ _0847_/A _0847_/B _0847_/C _0793_/D vssd1 vssd1 vccd1 vccd1 _0763_/A sky130_fd_sc_hd__or4_1
X_0831_ input5/X vssd1 vssd1 vccd1 vccd1 _1246_/A sky130_fd_sc_hd__inv_2
XANTENNA__1399__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1314_ _1333_/S vssd1 vssd1 vccd1 vccd1 _1336_/S sky130_fd_sc_hd__buf_2
X_1176_ peripheralBus_data[5] _1144_/A _1175_/X _1155_/X vssd1 vssd1 vccd1 vccd1 _1177_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1245_ _1250_/B _1236_/C _1379_/Q vssd1 vssd1 vccd1 vccd1 _1245_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1030_ _1030_/A vssd1 vssd1 vccd1 vccd1 _1030_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0814_ _0814_/A vssd1 vssd1 vccd1 vccd1 _0814_/X sky130_fd_sc_hd__clkbuf_1
Xinput20 peripheralBus_address[5] vssd1 vssd1 vccd1 vccd1 _0753_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1455__87 vssd1 vssd1 vccd1 vccd1 _1455__87/HI _1577_/A sky130_fd_sc_hd__conb_1
X_0745_ _1353_/A _1312_/B _1312_/C _0745_/D vssd1 vssd1 vccd1 vccd1 _1258_/C sky130_fd_sc_hd__or4_4
X_1228_ _1185_/X _1542_/A _1228_/S vssd1 vssd1 vccd1 vccd1 _1229_/B sky130_fd_sc_hd__mux2_1
X_1159_ _1506_/A _1504_/A _1196_/S vssd1 vssd1 vccd1 vccd1 _1159_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1013_ _1021_/A _1021_/B _1015_/C _1015_/D vssd1 vssd1 vccd1 vccd1 _1014_/A sky130_fd_sc_hd__or4_1
XFILLER_19_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0728_ _1123_/A vssd1 vssd1 vccd1 vccd1 _0847_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1203__A _1225_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1425__57 vssd1 vssd1 vccd1 vccd1 _1425__57/HI _1531_/A sky130_fd_sc_hd__conb_1
XFILLER_33_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1562_ _1562_/A _1112_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[27] sky130_fd_sc_hd__ebufn_8
XFILLER_3_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1023__A _1065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0993_ _0993_/A vssd1 vssd1 vccd1 vccd1 _1005_/A sky130_fd_sc_hd__clkbuf_1
X_1495__127 vssd1 vssd1 vccd1 vccd1 _1495__127/HI _1625_/A sky130_fd_sc_hd__conb_1
X_1614_ _1614_/A _0776_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[15] sky130_fd_sc_hd__ebufn_8
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1545_ _1545_/A _1064_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[10] sky130_fd_sc_hd__ebufn_8
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1261_ _1269_/A _1261_/B vssd1 vssd1 vccd1 vccd1 _1262_/A sky130_fd_sc_hd__and2_1
X_1330_ peripheralBus_data[5] _1308_/S _1333_/S vssd1 vssd1 vccd1 vccd1 _1331_/B sky130_fd_sc_hd__mux2_1
X_1192_ _1504_/A _1509_/A _1540_/A vssd1 vssd1 vccd1 vccd1 _1192_/X sky130_fd_sc_hd__mux2_1
Xinput7 peripheralBus_address[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0976_ _0976_/A vssd1 vssd1 vccd1 vccd1 _0976_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1528_ _1528_/A _1022_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[25] sky130_fd_sc_hd__ebufn_8
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0830_ _1087_/A vssd1 vssd1 vccd1 vccd1 _1043_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0761_ _0761_/A vssd1 vssd1 vccd1 vccd1 _0761_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_1244_ _1378_/Q _1236_/X _1243_/Y _1147_/A vssd1 vssd1 vccd1 vccd1 _1378_/D sky130_fd_sc_hd__o211a_1
X_1313_ _1353_/A _1313_/B _1313_/C _1353_/D vssd1 vssd1 vccd1 vccd1 _1333_/S sky130_fd_sc_hd__or4_4
XFILLER_2_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1175_ _1508_/A _1174_/X _1175_/S vssd1 vssd1 vccd1 vccd1 _1175_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1031__A _1143_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0959_ _0959_/A vssd1 vssd1 vccd1 vccd1 _0959_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__0870__A _0931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1366__CLK _1378_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0813_ _0823_/A _0823_/B _0854_/C _0813_/D vssd1 vssd1 vccd1 vccd1 _0814_/A sky130_fd_sc_hd__or4_1
Xinput10 peripheralBus_address[18] vssd1 vssd1 vccd1 vccd1 _0743_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_14_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput21 peripheralBus_address[6] vssd1 vssd1 vccd1 vccd1 _0753_/D sky130_fd_sc_hd__clkbuf_1
X_0744_ input5/X input7/X input6/X vssd1 vssd1 vccd1 vccd1 _0745_/D sky130_fd_sc_hd__or3_1
X_1158_ _1158_/A vssd1 vssd1 vccd1 vccd1 _1360_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__0865__A _1141_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1227_ _1227_/A vssd1 vssd1 vccd1 vccd1 _1374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1089_ _1091_/A _1091_/B _1099_/C _1099_/D vssd1 vssd1 vccd1 vccd1 _1090_/A sky130_fd_sc_hd__or4_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1389__CLK _1396_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1012_ _1012_/A vssd1 vssd1 vccd1 vccd1 _1012_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0727_ _1107_/A vssd1 vssd1 vccd1 vccd1 _1123_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1268__B2 _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1268__A1 peripheralBus_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input24_A peripheralBus_address[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1630_ _1630_/A _0879_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[31] sky130_fd_sc_hd__ebufn_8
XANTENNA__1404__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1561_ _1561_/A _1110_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[26] sky130_fd_sc_hd__ebufn_8
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1214__A _1337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0992_ _0992_/A vssd1 vssd1 vccd1 vccd1 _0992_/X sky130_fd_sc_hd__clkbuf_1
X_1613_ _1613_/A _0772_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[14] sky130_fd_sc_hd__ebufn_8
X_1544_ _1544_/A _1062_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[9] sky130_fd_sc_hd__ebufn_8
XFILLER_8_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1191_ _1503_/A _1510_/A _1540_/A vssd1 vssd1 vccd1 vccd1 _1191_/X sky130_fd_sc_hd__mux2_1
Xinput8 peripheralBus_address[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
X_1260_ _1253_/X _1257_/X _1259_/X _1145_/X vssd1 vssd1 vccd1 vccd1 _1261_/B sky130_fd_sc_hd__a22o_1
XFILLER_51_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0975_ _0977_/A _0977_/B _0985_/C _0985_/D vssd1 vssd1 vccd1 vccd1 _0976_/A sky130_fd_sc_hd__or4_1
X_1527_ _1527_/A _1020_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[24] sky130_fd_sc_hd__ebufn_8
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1389_ _1396_/CLK _1389_/D vssd1 vssd1 vccd1 vccd1 _1574_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0760_ _0847_/A _0847_/B _1123_/D _0775_/D vssd1 vssd1 vccd1 vccd1 _0761_/A sky130_fd_sc_hd__or4_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1174_ _1509_/A _1507_/A _1186_/S vssd1 vssd1 vccd1 vccd1 _1174_/X sky130_fd_sc_hd__mux2_1
X_1312_ input5/X _1312_/B _1312_/C _1312_/D vssd1 vssd1 vccd1 vccd1 _1353_/D sky130_fd_sc_hd__or4_2
X_1243_ _1378_/Q _1242_/Y _1236_/X vssd1 vssd1 vccd1 vccd1 _1243_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0958_ _0963_/A _0963_/B _0958_/C _0969_/D vssd1 vssd1 vccd1 vccd1 _0959_/A sky130_fd_sc_hd__or4_1
X_0889_ _0892_/A _0892_/B _0898_/C _0889_/D vssd1 vssd1 vccd1 vccd1 _0890_/A sky130_fd_sc_hd__or4_1
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0748__D _0793_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0812_ _0928_/A vssd1 vssd1 vccd1 vccd1 _0854_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput11 peripheralBus_address[19] vssd1 vssd1 vccd1 vccd1 _0743_/B sky130_fd_sc_hd__clkbuf_1
X_0743_ input9/X _0743_/B _0743_/C input8/X vssd1 vssd1 vccd1 vccd1 _1312_/C sky130_fd_sc_hd__or4b_2
Xinput22 peripheralBus_address[7] vssd1 vssd1 vccd1 vccd1 _0753_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1468__100 vssd1 vssd1 vccd1 vccd1 _1468__100/HI _1590_/A sky130_fd_sc_hd__conb_1
XFILLER_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1157_ _1177_/A _1157_/B vssd1 vssd1 vccd1 vccd1 _1158_/A sky130_fd_sc_hd__and2_1
XFILLER_37_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1226_ _1334_/A _1226_/B vssd1 vssd1 vccd1 vccd1 _1227_/A sky130_fd_sc_hd__or2_1
X_1446__78 vssd1 vssd1 vccd1 vccd1 _1446__78/HI _1560_/A sky130_fd_sc_hd__conb_1
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1088_ _1088_/A vssd1 vssd1 vccd1 vccd1 _1099_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1460__92 vssd1 vssd1 vccd1 vccd1 _1460__92/HI _1582_/A sky130_fd_sc_hd__conb_1
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1011_ _1021_/A _1021_/B _1015_/C _1015_/D vssd1 vssd1 vccd1 vccd1 _1012_/A sky130_fd_sc_hd__or4_1
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0966__A _0994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0726_ _1141_/A vssd1 vssd1 vccd1 vccd1 _1107_/A sky130_fd_sc_hd__buf_2
XANTENNA__1037__A _1065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1209_ _1209_/A vssd1 vssd1 vccd1 vccd1 _1369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input17_A peripheralBus_address[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0952__C _0958_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1560_ _1560_/A _1106_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[25] sky130_fd_sc_hd__ebufn_8
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1416__48 vssd1 vssd1 vccd1 vccd1 _1416__48/HI _1522_/A sky130_fd_sc_hd__conb_1
XANTENNA__1379__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input9_A peripheralBus_address[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1430__62 vssd1 vssd1 vccd1 vccd1 _1430__62/HI _1544_/A sky130_fd_sc_hd__conb_1
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0991_ _0991_/A _0991_/B _0999_/C _0999_/D vssd1 vssd1 vccd1 vccd1 _0992_/A sky130_fd_sc_hd__or4_1
XFILLER_8_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1612_ _1612_/A _0767_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[13] sky130_fd_sc_hd__ebufn_8
X_1543_ _1543_/A _1058_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[8] sky130_fd_sc_hd__ebufn_8
XFILLER_5_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0857__C _0912_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput9 peripheralBus_address[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
X_1190_ _1190_/A vssd1 vssd1 vccd1 vccd1 _1366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0974_ _1001_/A vssd1 vssd1 vccd1 vccd1 _0985_/C sky130_fd_sc_hd__clkbuf_1
X_1526_ _1526_/A _1016_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[23] sky130_fd_sc_hd__ebufn_8
XFILLER_35_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1388_ _1396_/CLK _1388_/D vssd1 vssd1 vccd1 vccd1 _1573_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1485__117 vssd1 vssd1 vccd1 vccd1 _1485__117/HI _1615_/A sky130_fd_sc_hd__conb_1
XFILLER_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1311_ _1311_/A vssd1 vssd1 vccd1 vccd1 _1390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1173_ _1173_/A vssd1 vssd1 vccd1 vccd1 _1363_/D sky130_fd_sc_hd__clkbuf_1
X_1242_ _1379_/Q _1236_/C _1250_/B vssd1 vssd1 vccd1 vccd1 _1242_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0957_ _1018_/A vssd1 vssd1 vccd1 vccd1 _0969_/D sky130_fd_sc_hd__clkbuf_2
X_0888_ _0888_/A vssd1 vssd1 vccd1 vccd1 _0888_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1509_ _1509_/A _0964_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[6] sky130_fd_sc_hd__ebufn_8
XANTENNA__1298__A0 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0811_ _0850_/A vssd1 vssd1 vccd1 vccd1 _0823_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_52_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0742_ _0742_/A _0742_/B _0742_/C _0742_/D vssd1 vssd1 vccd1 vccd1 _1312_/B sky130_fd_sc_hd__or4_4
Xinput12 peripheralBus_address[1] vssd1 vssd1 vccd1 vccd1 _0752_/A sky130_fd_sc_hd__clkbuf_1
Xinput23 peripheralBus_address[8] vssd1 vssd1 vccd1 vccd1 _0754_/B sky130_fd_sc_hd__clkbuf_1
X_1156_ peripheralBus_data[1] _1144_/X _1154_/X _1155_/X vssd1 vssd1 vccd1 vccd1 _1157_/B
+ sky130_fd_sc_hd__a22o_1
X_1087_ _1087_/A vssd1 vssd1 vccd1 vccd1 _1099_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1225_ peripheralBus_data[6] _1541_/A _1225_/S vssd1 vssd1 vccd1 vccd1 _1226_/B sky130_fd_sc_hd__mux2_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1204__A0 _1145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1010_ _1066_/A vssd1 vssd1 vccd1 vccd1 _1021_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1143__A _1143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output30_A _1128_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1208_ _1208_/A _1208_/B vssd1 vssd1 vccd1 vccd1 _1209_/A sky130_fd_sc_hd__and2_1
XFILLER_40_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1139_ _1377_/Q _1376_/Q _1538_/A vssd1 vssd1 vccd1 vccd1 _1193_/S sky130_fd_sc_hd__mux2_2
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0952__D _0954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0797__A _0867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0963__C _0972_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0990_ _0990_/A vssd1 vssd1 vccd1 vccd1 _0990_/X sky130_fd_sc_hd__clkbuf_1
X_1611_ _1611_/A _0769_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[12] sky130_fd_sc_hd__ebufn_8
XFILLER_8_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1542_ _1542_/A _1056_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[7] sky130_fd_sc_hd__ebufn_8
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0958__C _0958_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1369__CLK _1378_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0973_ _0973_/A vssd1 vssd1 vccd1 vccd1 _0973_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1525_ _1525_/A _1014_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[22] sky130_fd_sc_hd__ebufn_8
X_1387_ _1396_/CLK _1387_/D vssd1 vssd1 vccd1 vccd1 _1572_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1467__99 vssd1 vssd1 vccd1 vccd1 _1467__99/HI _1589_/A sky130_fd_sc_hd__conb_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1241_ _1348_/A _1241_/B vssd1 vssd1 vccd1 vccd1 _1377_/D sky130_fd_sc_hd__nor2_1
X_1310_ _1325_/A _1310_/B vssd1 vssd1 vccd1 vccd1 _1311_/A sky130_fd_sc_hd__and2_1
XFILLER_1_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1172_ _1177_/A _1172_/B vssd1 vssd1 vccd1 vccd1 _1173_/A sky130_fd_sc_hd__and2_1
XFILLER_52_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0956_ _1143_/C vssd1 vssd1 vccd1 vccd1 _1018_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0887_ _0892_/A _0892_/B _0898_/C _0889_/D vssd1 vssd1 vccd1 vccd1 _0888_/A sky130_fd_sc_hd__or4_1
XFILLER_55_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1508_ _1508_/A _0962_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[5] sky130_fd_sc_hd__ebufn_8
XFILLER_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1289__A1 peripheralBus_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0810_ _0849_/A vssd1 vssd1 vccd1 vccd1 _0823_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 peripheralBus_address[20] vssd1 vssd1 vccd1 vccd1 _0742_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0741_ input4/X vssd1 vssd1 vccd1 vccd1 _1353_/A sky130_fd_sc_hd__inv_2
Xinput24 peripheralBus_address[9] vssd1 vssd1 vccd1 vccd1 _0754_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_37_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1224_ _1224_/A vssd1 vssd1 vccd1 vccd1 _1334_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1155_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1155_/X sky130_fd_sc_hd__clkbuf_2
X_1086_ _1086_/A vssd1 vssd1 vccd1 vccd1 _1086_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0939_ _0939_/A vssd1 vssd1 vccd1 vccd1 _0939_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1437__69 vssd1 vssd1 vccd1 vccd1 _1437__69/HI _1551_/A sky130_fd_sc_hd__conb_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1143__B _1258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1451__83 vssd1 vssd1 vccd1 vccd1 _1451__83/HI _1565_/A sky130_fd_sc_hd__conb_1
XFILLER_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1207_ peripheralBus_data[1] _1536_/A _1228_/S vssd1 vssd1 vccd1 vccd1 _1208_/B sky130_fd_sc_hd__mux2_1
X_1138_ _1504_/A input29/X _1186_/S vssd1 vssd1 vccd1 vccd1 _1138_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1069_ _1077_/A _1077_/B _1071_/C _1071_/D vssd1 vssd1 vccd1 vccd1 _1070_/A sky130_fd_sc_hd__or4_1
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0993__A _0993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1407__39 vssd1 vssd1 vccd1 vccd1 _1407__39/HI _1513_/A sky130_fd_sc_hd__conb_1
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input22_A peripheralBus_address[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0963__D _0969_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1421__53 vssd1 vssd1 vccd1 vccd1 _1421__53/HI _1527_/A sky130_fd_sc_hd__conb_1
X_1610_ _1610_/A _0853_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[11] sky130_fd_sc_hd__ebufn_8
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1541_ _1541_/A _1054_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[6] sky130_fd_sc_hd__ebufn_8
XFILLER_5_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0873__D _0873_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0958__D _0969_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1307__A0 _1390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0972_ _0977_/A _0977_/B _0972_/C _0985_/D vssd1 vssd1 vccd1 vccd1 _0973_/A sky130_fd_sc_hd__or4_1
X_1524_ _1524_/A _1012_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[21] sky130_fd_sc_hd__ebufn_8
XANTENNA__1029__D _1029_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0868__D _0873_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1386_ _1396_/CLK _1386_/D vssd1 vssd1 vccd1 vccd1 _1571_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0969__C _0972_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1171_ peripheralBus_data[4] _1144_/A _1170_/X _1155_/X vssd1 vssd1 vccd1 vccd1 _1172_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1240_ _1236_/A _1377_/Q _1239_/Y _1236_/X vssd1 vssd1 vccd1 vccd1 _1241_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0955_ _0955_/A vssd1 vssd1 vccd1 vccd1 _0955_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0886_ _1258_/C vssd1 vssd1 vccd1 vccd1 _0898_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1507_ _1507_/A _0959_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[4] sky130_fd_sc_hd__ebufn_8
XANTENNA__1337__A _1337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1369_ _1378_/CLK _1369_/D vssd1 vssd1 vccd1 vccd1 _1536_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1491__123 vssd1 vssd1 vccd1 vccd1 _1491__123/HI _1621_/A sky130_fd_sc_hd__conb_1
XANTENNA__1359__CLK _1378_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 peripheralBus_address[21] vssd1 vssd1 vccd1 vccd1 _0742_/A sky130_fd_sc_hd__clkbuf_1
X_0740_ _1123_/C vssd1 vssd1 vccd1 vccd1 _0847_/C sky130_fd_sc_hd__clkbuf_2
Xinput25 peripheralBus_oe vssd1 vssd1 vccd1 vccd1 _0729_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1154_ _1504_/A _1152_/X _1175_/S vssd1 vssd1 vccd1 vccd1 _1154_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1223_ _1223_/A vssd1 vssd1 vccd1 vccd1 _1373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1085_ _1091_/A _1091_/B _1085_/C _1085_/D vssd1 vssd1 vccd1 vccd1 _1086_/A sky130_fd_sc_hd__or4_1
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0869_ _0869_/A vssd1 vssd1 vccd1 vccd1 _0869_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1475__107 vssd1 vssd1 vccd1 vccd1 _1475__107/HI _1597_/A sky130_fd_sc_hd__conb_1
X_0938_ _0948_/A _0948_/B _0942_/C _0946_/D vssd1 vssd1 vccd1 vccd1 _0939_/A sky130_fd_sc_hd__or4_1
XFILLER_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1143__C _1143_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1137_ _1540_/A vssd1 vssd1 vccd1 vccd1 _1186_/S sky130_fd_sc_hd__clkbuf_2
X_1206_ _1206_/A vssd1 vssd1 vccd1 vccd1 _1368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1068_ _1068_/A vssd1 vssd1 vccd1 vccd1 _1068_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input15_A peripheralBus_address[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1540_ _1540_/A _1122_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[5] sky130_fd_sc_hd__ebufn_8
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1392__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A peripheralBus_address[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0971_ _1018_/A vssd1 vssd1 vccd1 vccd1 _0985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1523_ _1523_/A _1006_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[20] sky130_fd_sc_hd__ebufn_8
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1385_ _1396_/CLK _1385_/D vssd1 vssd1 vccd1 vccd1 _1570_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1225__A0 peripheralBus_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0969__D _0969_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1170_ _1507_/A _1169_/X _1175_/S vssd1 vssd1 vccd1 vccd1 _1170_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0954_ _0963_/A _0963_/B _0958_/C _0954_/D vssd1 vssd1 vccd1 vccd1 _0955_/A sky130_fd_sc_hd__or4_1
XFILLER_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0885_ _0885_/A vssd1 vssd1 vccd1 vccd1 _0885_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1506_ _1506_/A _0955_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[3] sky130_fd_sc_hd__ebufn_8
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1368_ _1378_/CLK _1368_/D vssd1 vssd1 vccd1 vccd1 _1535_/A sky130_fd_sc_hd__dfxtp_1
X_1299_ _1574_/A _1298_/X _1305_/S vssd1 vssd1 vccd1 vccd1 _1299_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1207__A0 peripheralBus_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput15 peripheralBus_address[22] vssd1 vssd1 vccd1 vccd1 _0742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput26 peripheralBus_we vssd1 vssd1 vccd1 vccd1 _1141_/A sky130_fd_sc_hd__clkbuf_4
X_1153_ _1193_/S vssd1 vssd1 vccd1 vccd1 _1175_/S sky130_fd_sc_hd__clkbuf_2
X_1084_ _1084_/A vssd1 vssd1 vccd1 vccd1 _1084_/X sky130_fd_sc_hd__clkbuf_1
X_1222_ _1222_/A _1222_/B vssd1 vssd1 vccd1 vccd1 _1223_/A sky130_fd_sc_hd__or2_1
XFILLER_52_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0799_ _0799_/A vssd1 vssd1 vccd1 vccd1 _0799_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0937_ _0994_/A vssd1 vssd1 vccd1 vccd1 _0948_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_0868_ _0878_/A _0878_/B _0884_/C _0873_/D vssd1 vssd1 vccd1 vccd1 _0869_/A sky130_fd_sc_hd__or4_1
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1258__A _1267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0800__A _1258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1136_ _1143_/A vssd1 vssd1 vccd1 vccd1 _1155_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1205_ _1208_/A _1205_/B vssd1 vssd1 vccd1 vccd1 _1206_/A sky130_fd_sc_hd__and2_1
X_1067_ _1077_/A _1077_/B _1071_/C _1071_/D vssd1 vssd1 vccd1 vccd1 _1068_/A sky130_fd_sc_hd__or4_1
XFILLER_18_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1442__74 vssd1 vssd1 vccd1 vccd1 _1442__74/HI _1556_/A sky130_fd_sc_hd__conb_1
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1119_ _1123_/A _1123_/B _1121_/C _1121_/D vssd1 vssd1 vccd1 vccd1 _1120_/A sky130_fd_sc_hd__or4_1
XFILLER_29_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1412__44 vssd1 vssd1 vccd1 vccd1 _1412__44/HI _1518_/A sky130_fd_sc_hd__conb_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1599_ _1599_/A _0905_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[0] sky130_fd_sc_hd__ebufn_8
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0970_ _0970_/A vssd1 vssd1 vccd1 vccd1 _0970_/X sky130_fd_sc_hd__clkbuf_1
X_1522_ _1522_/A _1004_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[19] sky130_fd_sc_hd__ebufn_8
X_1384_ _1396_/CLK _1384_/D vssd1 vssd1 vccd1 vccd1 _1569_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1382__CLK _1396_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0953_ _0953_/A vssd1 vssd1 vccd1 vccd1 _0953_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0884_ _0892_/A _0892_/B _0884_/C _0889_/D vssd1 vssd1 vccd1 vccd1 _0885_/A sky130_fd_sc_hd__or4_1
X_1367_ _1367_/CLK _1367_/D vssd1 vssd1 vccd1 vccd1 _1367_/Q sky130_fd_sc_hd__dfxtp_1
X_1505_ _1505_/A _0953_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[2] sky130_fd_sc_hd__ebufn_8
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1298_ input28/X _1573_/A _1298_/S vssd1 vssd1 vccd1 vccd1 _1298_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1448__80 vssd1 vssd1 vccd1 vccd1 _1448__80/HI _1562_/A sky130_fd_sc_hd__conb_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput27 rst vssd1 vssd1 vccd1 vccd1 _1224_/A sky130_fd_sc_hd__buf_2
Xinput16 peripheralBus_address[23] vssd1 vssd1 vccd1 vccd1 _0742_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_52_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1221_ peripheralBus_data[5] _1196_/S _1225_/S vssd1 vssd1 vccd1 vccd1 _1222_/B sky130_fd_sc_hd__mux2_1
XFILLER_35_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1152_ _1505_/A _1503_/A _1196_/S vssd1 vssd1 vccd1 vccd1 _1152_/X sky130_fd_sc_hd__mux2_1
X_1083_ _1091_/A _1091_/B _1085_/C _1085_/D vssd1 vssd1 vccd1 vccd1 _1084_/A sky130_fd_sc_hd__or4_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0936_ _1141_/B vssd1 vssd1 vccd1 vccd1 _0994_/A sky130_fd_sc_hd__buf_2
XFILLER_20_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0798_ _0808_/A _0808_/B _0840_/C _0818_/D vssd1 vssd1 vccd1 vccd1 _0799_/A sky130_fd_sc_hd__or4_1
X_0867_ _0867_/A vssd1 vssd1 vccd1 vccd1 _0884_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1258__B _1258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1204_ _1145_/X _1535_/A _1228_/S vssd1 vssd1 vccd1 vccd1 _1205_/B sky130_fd_sc_hd__mux2_1
XANTENNA__1355__B1 _1147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1066_ _1066_/A vssd1 vssd1 vccd1 vccd1 _1077_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1481__113 vssd1 vssd1 vccd1 vccd1 _1481__113/HI _1611_/A sky130_fd_sc_hd__conb_1
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1135_ _1381_/Q vssd1 vssd1 vccd1 vccd1 _1143_/A sky130_fd_sc_hd__clkinv_2
X_0919_ _0919_/A vssd1 vssd1 vccd1 vccd1 _0919_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1418__50 vssd1 vssd1 vccd1 vccd1 _1418__50/HI _1524_/A sky130_fd_sc_hd__conb_1
XFILLER_33_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1269__A _1269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1179__A _1337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1118_ _1118_/A vssd1 vssd1 vccd1 vccd1 _1118_/X sky130_fd_sc_hd__clkbuf_1
X_1049_ _1049_/A _1049_/B _1057_/C _1057_/D vssd1 vssd1 vccd1 vccd1 _1050_/A sky130_fd_sc_hd__or4_1
XFILLER_21_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1598_ _1598_/A _0876_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[31] sky130_fd_sc_hd__ebufn_8
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input20_A peripheralBus_address[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1221__S _1225_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1521_ _1521_/A _1000_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[18] sky130_fd_sc_hd__ebufn_8
X_1383_ _1396_/CLK _1383_/D vssd1 vssd1 vccd1 vccd1 _1568_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1161__A1 peripheralBus_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0952_ _0963_/A _0963_/B _0958_/C _0954_/D vssd1 vssd1 vccd1 vccd1 _0953_/A sky130_fd_sc_hd__or4_1
XFILLER_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1504_ _1504_/A _0949_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[1] sky130_fd_sc_hd__ebufn_8
X_0883_ _0883_/A vssd1 vssd1 vccd1 vccd1 _0883_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1366_ _1378_/CLK _1366_/D vssd1 vssd1 vccd1 vccd1 _1510_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1297_ _1297_/A vssd1 vssd1 vccd1 vccd1 _1325_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1463__95 vssd1 vssd1 vccd1 vccd1 _1463__95/HI _1585_/A sky130_fd_sc_hd__conb_1
Xinput28 spi_miso[0] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_2
Xinput17 peripheralBus_address[2] vssd1 vssd1 vccd1 vccd1 _0755_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1151_ _1540_/A vssd1 vssd1 vccd1 vccd1 _1196_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1220_ _1220_/A vssd1 vssd1 vccd1 vccd1 _1372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1082_ _1082_/A vssd1 vssd1 vccd1 vccd1 _1082_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0935_ _0993_/A vssd1 vssd1 vccd1 vccd1 _0948_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0866_ _0921_/A vssd1 vssd1 vccd1 vccd1 _0878_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_0797_ _0867_/A vssd1 vssd1 vccd1 vccd1 _0840_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_1349_ _1402_/Q _1343_/C _1403_/Q vssd1 vssd1 vccd1 vccd1 _1349_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1258__C _1258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1372__CLK _1378_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1290__A _1295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1203_ _1225_/S vssd1 vssd1 vccd1 vccd1 _1228_/S sky130_fd_sc_hd__clkbuf_2
X_1134_ _1297_/A vssd1 vssd1 vccd1 vccd1 _1147_/A sky130_fd_sc_hd__buf_2
X_1065_ _1065_/A vssd1 vssd1 vccd1 vccd1 _1077_/A sky130_fd_sc_hd__clkbuf_1
X_0849_ _0849_/A vssd1 vssd1 vccd1 vccd1 _0861_/A sky130_fd_sc_hd__clkbuf_1
X_0918_ _0918_/A _0918_/B _0926_/C _0929_/D vssd1 vssd1 vccd1 vccd1 _0919_/A sky130_fd_sc_hd__or4_1
XANTENNA__1395__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1433__65 vssd1 vssd1 vccd1 vccd1 _1433__65/HI _1547_/A sky130_fd_sc_hd__conb_1
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1285__A _1295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1117_ _1117_/A _1117_/B _1121_/C _1121_/D vssd1 vssd1 vccd1 vccd1 _1118_/A sky130_fd_sc_hd__or4_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1048_ _1048_/A vssd1 vssd1 vccd1 vccd1 _1048_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0822__A _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1597_ _1597_/A _0872_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[30] sky130_fd_sc_hd__ebufn_8
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input13_A peripheralBus_address[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1228__A0 _1185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1520_ _1520_/A _0998_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[17] sky130_fd_sc_hd__ebufn_8
X_1382_ _1396_/CLK _1382_/D vssd1 vssd1 vccd1 vccd1 _1567_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input5_A peripheralBus_address[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0951_ _0994_/A vssd1 vssd1 vccd1 vccd1 _0963_/B sky130_fd_sc_hd__clkbuf_1
X_0882_ _0892_/A _0892_/B _0884_/C _0889_/D vssd1 vssd1 vccd1 vccd1 _0883_/A sky130_fd_sc_hd__or4_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1503_ _1503_/A _0848_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[0] sky130_fd_sc_hd__ebufn_8
X_1365_ _1367_/CLK _1365_/D vssd1 vssd1 vccd1 vccd1 _1509_/A sky130_fd_sc_hd__dfxtp_2
X_1296_ _1296_/A vssd1 vssd1 vccd1 vccd1 _1388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 peripheralBus_address[3] vssd1 vssd1 vccd1 vccd1 _0755_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput29 spi_miso[1] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1150_ _1337_/A vssd1 vssd1 vccd1 vccd1 _1177_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1439__71 vssd1 vssd1 vccd1 vccd1 _1439__71/HI _1553_/A sky130_fd_sc_hd__conb_1
X_1081_ _1091_/A _1091_/B _1085_/C _1085_/D vssd1 vssd1 vccd1 vccd1 _1082_/A sky130_fd_sc_hd__or4_1
X_0934_ _1141_/A vssd1 vssd1 vccd1 vccd1 _0993_/A sky130_fd_sc_hd__buf_2
X_0865_ _1141_/B vssd1 vssd1 vccd1 vccd1 _0921_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0796_ _0850_/A vssd1 vssd1 vccd1 vccd1 _0808_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1348_ _1348_/A _1348_/B vssd1 vssd1 vccd1 vccd1 _1400_/D sky130_fd_sc_hd__nor2_1
X_1279_ peripheralBus_data[3] _1259_/X _1278_/X _1357_/A vssd1 vssd1 vccd1 vccd1 _1280_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1202_ _1246_/A _1202_/B _1353_/C _1246_/D vssd1 vssd1 vccd1 vccd1 _1225_/S sky130_fd_sc_hd__or4_4
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1064_ _1064_/A vssd1 vssd1 vccd1 vccd1 _1064_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1133_ _1224_/A vssd1 vssd1 vccd1 vccd1 _1297_/A sky130_fd_sc_hd__inv_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0779_ _1108_/A vssd1 vssd1 vccd1 vccd1 _0850_/A sky130_fd_sc_hd__clkbuf_2
X_0848_ _0848_/A vssd1 vssd1 vccd1 vccd1 _0848_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0917_ _0931_/A vssd1 vssd1 vccd1 vccd1 _0929_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1409__41 vssd1 vssd1 vccd1 vccd1 _1409__41/HI _1515_/A sky130_fd_sc_hd__conb_1
XFILLER_30_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1116_ _1116_/A vssd1 vssd1 vccd1 vccd1 _1116_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1047_ _1049_/A _1049_/B _1057_/C _1057_/D vssd1 vssd1 vccd1 vccd1 _1048_/A sky130_fd_sc_hd__or4_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1255__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1471__103 vssd1 vssd1 vccd1 vccd1 _1471__103/HI _1593_/A sky130_fd_sc_hd__conb_1
XFILLER_62_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1385__CLK _1396_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1596_ _1596_/A _0858_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[29] sky130_fd_sc_hd__ebufn_8
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1381_ _1404_/CLK _1381_/D vssd1 vssd1 vccd1 vccd1 _1381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ _1579_/A _0947_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[12] sky130_fd_sc_hd__ebufn_8
XANTENNA__1400__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0950_ _0993_/A vssd1 vssd1 vccd1 vccd1 _0963_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_9_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0881_ _0921_/A vssd1 vssd1 vccd1 vccd1 _0892_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1364_ _1367_/CLK _1364_/D vssd1 vssd1 vccd1 vccd1 _1508_/A sky130_fd_sc_hd__dfxtp_1
X_1295_ _1295_/A _1295_/B vssd1 vssd1 vccd1 vccd1 _1296_/A sky130_fd_sc_hd__and2_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0738__A _1258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput19 peripheralBus_address[4] vssd1 vssd1 vccd1 vccd1 _0753_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_10_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1080_ _1108_/A vssd1 vssd1 vccd1 vccd1 _1091_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0795_ _0849_/A vssd1 vssd1 vccd1 vccd1 _0808_/A sky130_fd_sc_hd__clkbuf_1
X_1454__86 vssd1 vssd1 vccd1 vccd1 _1454__86/HI _1576_/A sky130_fd_sc_hd__conb_1
XANTENNA__1358__B1 _1147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0933_ _0933_/A vssd1 vssd1 vccd1 vccd1 _0933_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0864_ _0920_/A vssd1 vssd1 vccd1 vccd1 _0878_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1347_ _1357_/B _1400_/Q _1346_/Y _1343_/X vssd1 vssd1 vccd1 vccd1 _1348_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1278_ _1570_/A _1277_/X _1288_/S vssd1 vssd1 vccd1 vccd1 _1278_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0931__A _0931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1201_ input4/X _1312_/B _1312_/C _1312_/D vssd1 vssd1 vccd1 vccd1 _1246_/D sky130_fd_sc_hd__or4_2
XFILLER_2_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1063_ _1063_/A _1063_/B _1071_/C _1071_/D vssd1 vssd1 vccd1 vccd1 _1064_/A sky130_fd_sc_hd__or4_1
X_1132_ _1606_/A _1128_/B _1131_/Y vssd1 vssd1 vccd1 vccd1 _1132_/X sky130_fd_sc_hd__o21a_1
XFILLER_18_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0916_ _0916_/A vssd1 vssd1 vccd1 vccd1 _0916_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0778_ _0849_/A vssd1 vssd1 vccd1 vccd1 _0793_/A sky130_fd_sc_hd__clkbuf_1
X_0847_ _0847_/A _0847_/B _0847_/C _0954_/D vssd1 vssd1 vccd1 vccd1 _0848_/A sky130_fd_sc_hd__or4_1
XFILLER_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0751__A _0867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1424__56 vssd1 vssd1 vccd1 vccd1 _1424__56/HI _1530_/A sky130_fd_sc_hd__conb_1
XFILLER_38_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1115_ _1117_/A _1117_/B _1121_/C _1121_/D vssd1 vssd1 vccd1 vccd1 _1116_/A sky130_fd_sc_hd__or4_1
X_1046_ _1088_/A vssd1 vssd1 vccd1 vccd1 _1057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0746__A _1258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0912__C _0912_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1191__A1 _1510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1595_ _1595_/A _0855_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[28] sky130_fd_sc_hd__ebufn_8
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1182__A1 peripheralBus_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1029_ _1035_/A _1035_/B _1029_/C _1029_/D vssd1 vssd1 vccd1 vccd1 _1030_/A sky130_fd_sc_hd__or4_1
X_1494__126 vssd1 vssd1 vccd1 vccd1 _1494__126/HI _1624_/A sky130_fd_sc_hd__conb_1
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1380_ _1404_/CLK _1380_/D vssd1 vssd1 vccd1 vccd1 _1380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1010__A _1066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1578_ _1578_/A _0943_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[11] sky130_fd_sc_hd__ebufn_8
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1375__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1146__B2 _1145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0934__A _1141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0880_ _0920_/A vssd1 vssd1 vccd1 vccd1 _0892_/A sky130_fd_sc_hd__clkbuf_1
X_1363_ _1367_/CLK _1363_/D vssd1 vssd1 vccd1 vccd1 _1507_/A sky130_fd_sc_hd__dfxtp_1
X_1294_ peripheralBus_data[6] _1259_/A _1293_/X _1253_/X vssd1 vssd1 vccd1 vccd1 _1295_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1398__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1300__A1 _1185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0904__D _1043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0932_ _0932_/A _0932_/B _0942_/C _0946_/D vssd1 vssd1 vccd1 vccd1 _0933_/A sky130_fd_sc_hd__or4_1
XFILLER_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0794_ _0794_/A vssd1 vssd1 vccd1 vccd1 _0794_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0863_ _1141_/A vssd1 vssd1 vccd1 vccd1 _0920_/A sky130_fd_sc_hd__clkbuf_2
X_1346_ _1603_/A vssd1 vssd1 vccd1 vccd1 _1346_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1277_ _1571_/A _1569_/A _1308_/S vssd1 vssd1 vccd1 vccd1 _1277_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1200_ input7/X input6/X vssd1 vssd1 vccd1 vccd1 _1312_/D sky130_fd_sc_hd__or2_1
XFILLER_2_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1062_ _1062_/A vssd1 vssd1 vccd1 vccd1 _1062_/X sky130_fd_sc_hd__clkbuf_1
X_1131_ _1606_/A _1128_/B _1605_/A vssd1 vssd1 vccd1 vccd1 _1131_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0915_ _0918_/A _0918_/B _0926_/C _0915_/D vssd1 vssd1 vccd1 vccd1 _0916_/A sky130_fd_sc_hd__or4_1
X_0846_ _0846_/A vssd1 vssd1 vccd1 vccd1 _0846_/X sky130_fd_sc_hd__clkbuf_1
X_0777_ _1107_/A vssd1 vssd1 vccd1 vccd1 _0849_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1329_ _1329_/A vssd1 vssd1 vccd1 vccd1 _1395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input29_A spi_miso[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1114_ _1114_/A vssd1 vssd1 vccd1 vccd1 _1114_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1045_ _1087_/A vssd1 vssd1 vccd1 vccd1 _1057_/C sky130_fd_sc_hd__clkbuf_1
X_0829_ _1202_/B vssd1 vssd1 vccd1 vccd1 _1087_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0937__A _0994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1594_ _1594_/A _0828_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[27] sky130_fd_sc_hd__ebufn_8
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1008__A _1065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1182__A2 _1144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1028_ _1028_/A vssd1 vssd1 vccd1 vccd1 _1028_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0757__A _1313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1577_ _1577_/A _0941_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[10] sky130_fd_sc_hd__ebufn_8
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1502__134 vssd1 vssd1 vccd1 vccd1 _1502__134/HI spi_en[1] sky130_fd_sc_hd__conb_1
XFILLER_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input11_A peripheralBus_address[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0950__A _0993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1362_ _1367_/CLK _1362_/D vssd1 vssd1 vccd1 vccd1 _1506_/A sky130_fd_sc_hd__dfxtp_1
X_1293_ _1573_/A _1292_/X _1305_/S vssd1 vssd1 vccd1 vccd1 _1293_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1629_ _1629_/A _0874_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[30] sky130_fd_sc_hd__ebufn_8
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input3_A peripheralBus_address[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0770__A _0867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0862_ _0862_/A vssd1 vssd1 vccd1 vccd1 _0862_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0931_ _0931_/A vssd1 vssd1 vccd1 vccd1 _0946_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0793_ _0793_/A _0793_/B _0808_/C _0793_/D vssd1 vssd1 vccd1 vccd1 _0794_/A sky130_fd_sc_hd__or4_1
X_1345_ _1348_/A _1345_/B vssd1 vssd1 vccd1 vccd1 _1399_/D sky130_fd_sc_hd__nor2_1
X_1276_ _1276_/A vssd1 vssd1 vccd1 vccd1 _1384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1294__A1 peripheralBus_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1445__77 vssd1 vssd1 vccd1 vccd1 _1445__77/HI _1559_/A sky130_fd_sc_hd__conb_1
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1130_ _1542_/A _1128_/A _1129_/Y vssd1 vssd1 vccd1 vccd1 _1130_/X sky130_fd_sc_hd__o21a_1
XFILLER_2_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1061_ _1063_/A _1063_/B _1071_/C _1071_/D vssd1 vssd1 vccd1 vccd1 _1062_/A sky130_fd_sc_hd__or4_1
XANTENNA__1388__CLK _1396_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0845_ _0845_/A _0845_/B _0861_/C _0845_/D vssd1 vssd1 vccd1 vccd1 _0846_/A sky130_fd_sc_hd__or4_1
X_0914_ _0928_/A vssd1 vssd1 vccd1 vccd1 _0926_/C sky130_fd_sc_hd__clkbuf_1
X_0776_ _0776_/A vssd1 vssd1 vccd1 vccd1 _0776_/X sky130_fd_sc_hd__clkbuf_1
X_1259_ _1259_/A vssd1 vssd1 vccd1 vccd1 _1259_/X sky130_fd_sc_hd__clkbuf_2
X_1328_ _1337_/A _1328_/B vssd1 vssd1 vccd1 vccd1 _1329_/A sky130_fd_sc_hd__and2_1
XFILLER_33_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1113_ _1117_/A _1117_/B _1113_/C _1113_/D vssd1 vssd1 vccd1 vccd1 _1114_/A sky130_fd_sc_hd__or4_1
XANTENNA__0836__C _1043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1044_ _1044_/A vssd1 vssd1 vccd1 vccd1 _1044_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0828_ _0828_/A vssd1 vssd1 vccd1 vccd1 _0828_/X sky130_fd_sc_hd__clkbuf_1
X_1415__47 vssd1 vssd1 vccd1 vccd1 _1415__47/HI _1521_/A sky130_fd_sc_hd__conb_1
X_0759_ _1121_/C vssd1 vssd1 vccd1 vccd1 _0775_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1403__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1593_ _1593_/A _0821_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[26] sky130_fd_sc_hd__ebufn_8
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1027_ _1035_/A _1035_/B _1029_/C _1029_/D vssd1 vssd1 vccd1 vccd1 _1028_/A sky130_fd_sc_hd__or4_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1024__A _1066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0863__A _1141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1330__A0 peripheralBus_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1321__A0 peripheralBus_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1576_ _1576_/A _0939_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[9] sky130_fd_sc_hd__ebufn_8
XFILLER_58_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1361_ _1367_/CLK _1361_/D vssd1 vssd1 vccd1 vccd1 _1505_/A sky130_fd_sc_hd__dfxtp_1
X_1292_ _1574_/A _1572_/A _1298_/S vssd1 vssd1 vccd1 vccd1 _1292_/X sky130_fd_sc_hd__mux2_1
X_1484__116 vssd1 vssd1 vccd1 vccd1 _1484__116/HI _1614_/A sky130_fd_sc_hd__conb_1
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1559_ _1559_/A _1104_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[24] sky130_fd_sc_hd__ebufn_8
X_1628_ _1628_/A _0869_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[29] sky130_fd_sc_hd__ebufn_8
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0861_ _0861_/A _0861_/B _0861_/C _0873_/D vssd1 vssd1 vccd1 vccd1 _0862_/A sky130_fd_sc_hd__or4_1
X_0792_ _0928_/A vssd1 vssd1 vccd1 vccd1 _0808_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0930_ _0930_/A vssd1 vssd1 vccd1 vccd1 _0930_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1344_ _1357_/B _1399_/Q _1603_/A _1343_/X vssd1 vssd1 vccd1 vccd1 _1345_/B sky130_fd_sc_hd__o2bb2a_1
X_1275_ _1295_/A _1275_/B vssd1 vssd1 vccd1 vccd1 _1276_/A sky130_fd_sc_hd__and2_1
XFILLER_51_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0956__A _1143_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1060_ _1088_/A vssd1 vssd1 vccd1 vccd1 _1071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output35_A _1390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0844_ _0844_/A vssd1 vssd1 vccd1 vccd1 _0844_/X sky130_fd_sc_hd__clkbuf_1
X_0775_ _0775_/A _0775_/B _0789_/C _0775_/D vssd1 vssd1 vccd1 vccd1 _0776_/A sky130_fd_sc_hd__or4_1
X_0913_ _0913_/A vssd1 vssd1 vccd1 vccd1 _0913_/X sky130_fd_sc_hd__clkbuf_1
X_1189_ _1208_/A _1189_/B vssd1 vssd1 vccd1 vccd1 _1190_/A sky130_fd_sc_hd__and2_1
X_1327_ peripheralBus_data[4] _1603_/A _1336_/S vssd1 vssd1 vccd1 vccd1 _1328_/B sky130_fd_sc_hd__mux2_1
X_1258_ _1267_/A _1258_/B _1258_/C _1353_/C vssd1 vssd1 vccd1 vccd1 _1259_/A sky130_fd_sc_hd__nor4_4
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1112_ _1112_/A vssd1 vssd1 vccd1 vccd1 _1112_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0836__D _0954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1043_ _1049_/A _1049_/B _1043_/C _1043_/D vssd1 vssd1 vccd1 vccd1 _1044_/A sky130_fd_sc_hd__or4_1
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0827_ _0845_/A _0845_/B _0854_/C _0857_/D vssd1 vssd1 vccd1 vccd1 _0828_/A sky130_fd_sc_hd__or4_1
X_0758_ _1202_/B vssd1 vssd1 vccd1 vccd1 _1121_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1176__A1 peripheralBus_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1378__CLK _1378_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1592_ _1592_/A _0817_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[25] sky130_fd_sc_hd__ebufn_8
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1026_ _1026_/A vssd1 vssd1 vccd1 vccd1 _1026_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1575_ _1575_/A _0933_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[8] sky130_fd_sc_hd__ebufn_8
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1009_ _1141_/B vssd1 vssd1 vccd1 vccd1 _1066_/A sky130_fd_sc_hd__buf_2
XFILLER_25_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0784__A _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1466__98 vssd1 vssd1 vccd1 vccd1 _1466__98/HI _1588_/A sky130_fd_sc_hd__conb_1
XFILLER_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1360_ _1367_/CLK _1360_/D vssd1 vssd1 vccd1 vccd1 _1504_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1291_ _1291_/A vssd1 vssd1 vccd1 vccd1 _1387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1627_ _1627_/A _0860_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[28] sky130_fd_sc_hd__ebufn_8
X_1558_ _1558_/A _1100_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[23] sky130_fd_sc_hd__ebufn_8
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1221__A0 peripheralBus_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0860_ _0860_/A vssd1 vssd1 vccd1 vccd1 _0860_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0791_ _1353_/B vssd1 vssd1 vccd1 vccd1 _0928_/A sky130_fd_sc_hd__buf_2
XFILLER_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1343_ _1357_/B _1402_/Q _1343_/C vssd1 vssd1 vccd1 vccd1 _1343_/X sky130_fd_sc_hd__or3_1
XFILLER_51_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1274_ peripheralBus_data[2] _1259_/X _1273_/X _1357_/A vssd1 vssd1 vccd1 vccd1 _1275_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0989_ _0991_/A _0991_/B _0999_/C _0999_/D vssd1 vssd1 vccd1 vccd1 _0990_/A sky130_fd_sc_hd__or4_1
XFILLER_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1436__68 vssd1 vssd1 vccd1 vccd1 _1436__68/HI _1550_/A sky130_fd_sc_hd__conb_1
XFILLER_6_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1133__A _1224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0912_ _0918_/A _0918_/B _0912_/C _0915_/D vssd1 vssd1 vccd1 vccd1 _0913_/A sky130_fd_sc_hd__or4_1
X_0843_ _0845_/A _0845_/B _0861_/C _0845_/D vssd1 vssd1 vccd1 vccd1 _0844_/A sky130_fd_sc_hd__or4_1
X_1450__82 vssd1 vssd1 vccd1 vccd1 _1450__82/HI _1564_/A sky130_fd_sc_hd__conb_1
X_0774_ _0774_/A vssd1 vssd1 vccd1 vccd1 _0774_/X sky130_fd_sc_hd__clkbuf_1
X_1326_ _1326_/A vssd1 vssd1 vccd1 vccd1 _1394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1188_ _1185_/X _1144_/A _1187_/X _1155_/A vssd1 vssd1 vccd1 vccd1 _1189_/B sky130_fd_sc_hd__a22o_1
XFILLER_24_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1257_ _1567_/A _1255_/X _1305_/S vssd1 vssd1 vccd1 vccd1 _1257_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0792__A _0928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1351__C1 _1147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1111_ _1117_/A _1117_/B _1113_/C _1113_/D vssd1 vssd1 vccd1 vccd1 _1112_/A sky130_fd_sc_hd__or4_1
X_1042_ _1042_/A vssd1 vssd1 vccd1 vccd1 _1042_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0852__D _0873_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0826_ _0850_/A vssd1 vssd1 vccd1 vccd1 _0845_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__1038__A _1066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0757_ _1313_/B vssd1 vssd1 vccd1 vccd1 _1202_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0877__A _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1309_ _1253_/X _1307_/X _1308_/X _1259_/X vssd1 vssd1 vccd1 vccd1 _1310_/B sky130_fd_sc_hd__a22o_1
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0762__D _0793_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1406__38 vssd1 vssd1 vccd1 vccd1 _1406__38/HI _1512_/A sky130_fd_sc_hd__conb_1
XANTENNA__1176__A2 _1144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input27_A rst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1591_ _1591_/A _0814_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[24] sky130_fd_sc_hd__ebufn_8
X_1420__52 vssd1 vssd1 vccd1 vccd1 _1420__52/HI _1526_/A sky130_fd_sc_hd__conb_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0847__D _0954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1025_ _1035_/A _1035_/B _1029_/C _1029_/D vssd1 vssd1 vccd1 vccd1 _1026_/A sky130_fd_sc_hd__or4_1
XFILLER_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0809_ _0809_/A vssd1 vssd1 vccd1 vccd1 _0809_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0948__C _0958_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0980__A _0994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1141__A _1141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1574_ _1574_/A _0930_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[7] sky130_fd_sc_hd__ebufn_8
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1368__CLK _1378_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1051__A _1065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1008_ _1065_/A vssd1 vssd1 vccd1 vccd1 _1021_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1136__A _1143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1290_ _1295_/A _1290_/B vssd1 vssd1 vccd1 vccd1 _1291_/A sky130_fd_sc_hd__and2_1
XANTENNA__1021__D _1029_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1626_ _1626_/A _0862_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[27] sky130_fd_sc_hd__ebufn_8
X_1557_ _1557_/A _1098_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[22] sky130_fd_sc_hd__ebufn_8
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0961__C _0972_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1490__122 vssd1 vssd1 vccd1 vccd1 _1490__122/HI _1620_/A sky130_fd_sc_hd__conb_1
X_0790_ _0790_/A vssd1 vssd1 vccd1 vccd1 _0790_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1273_ _1569_/A _1272_/X _1288_/S vssd1 vssd1 vccd1 vccd1 _1273_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1342_ _1340_/X _1341_/Y _1601_/A _1600_/A vssd1 vssd1 vccd1 vccd1 _1343_/C sky130_fd_sc_hd__a211o_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1313__B _1313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1279__A1 peripheralBus_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1279__B2 _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0988_ _1018_/A vssd1 vssd1 vccd1 vccd1 _0999_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__0871__C _0912_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1609_ _1609_/A _0911_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[10] sky130_fd_sc_hd__ebufn_8
XANTENNA_input1_A peripheralBus_address[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1474__106 vssd1 vssd1 vccd1 vccd1 _1474__106/HI _1596_/A sky130_fd_sc_hd__conb_1
XFILLER_6_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0842_ _0867_/A vssd1 vssd1 vccd1 vccd1 _0861_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0911_ _0911_/A vssd1 vssd1 vccd1 vccd1 _0911_/X sky130_fd_sc_hd__clkbuf_1
X_0773_ _0775_/A _0775_/B _0847_/C _0793_/D vssd1 vssd1 vccd1 vccd1 _0774_/A sky130_fd_sc_hd__or4_1
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1325_ _1325_/A _1325_/B vssd1 vssd1 vccd1 vccd1 _1326_/A sky130_fd_sc_hd__and2_1
X_1256_ _1400_/Q _1399_/Q _1602_/A vssd1 vssd1 vccd1 vccd1 _1305_/S sky130_fd_sc_hd__mux2_4
XFILLER_17_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1187_ _1510_/A _1186_/X _1193_/S vssd1 vssd1 vccd1 vccd1 _1187_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1110_ _1110_/A vssd1 vssd1 vccd1 vccd1 _1110_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1144__A _1144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1041_ _1049_/A _1049_/B _1043_/C _1043_/D vssd1 vssd1 vccd1 vccd1 _1042_/A sky130_fd_sc_hd__or4_1
X_0825_ _0849_/A vssd1 vssd1 vccd1 vccd1 _0845_/A sky130_fd_sc_hd__clkbuf_1
X_0756_ _0756_/A _0756_/B _0756_/C _0756_/D vssd1 vssd1 vccd1 vccd1 _1313_/B sky130_fd_sc_hd__or4_2
XFILLER_56_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1239_ _1539_/A vssd1 vssd1 vccd1 vccd1 _1239_/Y sky130_fd_sc_hd__clkinv_2
X_1308_ peripheralBus_data[0] peripheralBus_data[7] _1308_/S vssd1 vssd1 vccd1 vccd1
+ _1308_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1229__A _1269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1333__A0 peripheralBus_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1590_ _1590_/A _0809_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[23] sky130_fd_sc_hd__ebufn_8
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1024_ _1066_/A vssd1 vssd1 vccd1 vccd1 _1035_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1324__A0 peripheralBus_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0808_ _0808_/A _0808_/B _0808_/C _0813_/D vssd1 vssd1 vccd1 vccd1 _0809_/A sky130_fd_sc_hd__or4_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0739_ _1353_/B vssd1 vssd1 vccd1 vccd1 _1123_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1315__A0 _1145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0773__D _0793_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0948__D _0954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1141__B _1141_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1019__D _1029_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ _1573_/A _0927_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[6] sky130_fd_sc_hd__ebufn_8
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1007_ _1141_/A vssd1 vssd1 vccd1 vccd1 _1065_/A sky130_fd_sc_hd__buf_2
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1457__89 vssd1 vssd1 vccd1 vccd1 _1457__89/HI _1579_/A sky130_fd_sc_hd__conb_1
XFILLER_16_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1625_ _1625_/A _0846_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[26] sky130_fd_sc_hd__ebufn_8
X_1556_ _1556_/A _1096_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[21] sky130_fd_sc_hd__ebufn_8
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0961__D _0969_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1147__A _1147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1272_ _1570_/A _1568_/A _1308_/S vssd1 vssd1 vccd1 vccd1 _1272_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1341_ _1401_/Q _1599_/A vssd1 vssd1 vccd1 vccd1 _1341_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0987_ _1001_/A vssd1 vssd1 vccd1 vccd1 _0999_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1539_ _1539_/A _1050_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[4] sky130_fd_sc_hd__ebufn_8
X_1608_ _1608_/A _0903_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[9] sky130_fd_sc_hd__ebufn_8
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0781__D _0793_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0972__C _0972_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0841_ _0841_/A vssd1 vssd1 vccd1 vccd1 _0841_/X sky130_fd_sc_hd__clkbuf_1
X_1427__59 vssd1 vssd1 vccd1 vccd1 _1427__59/HI _1533_/A sky130_fd_sc_hd__conb_1
XFILLER_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0772_ _0772_/A vssd1 vssd1 vccd1 vccd1 _0772_/X sky130_fd_sc_hd__clkbuf_1
X_0910_ _0918_/A _0918_/B _0910_/C _1043_/C vssd1 vssd1 vccd1 vccd1 _0911_/A sky130_fd_sc_hd__or4_1
XANTENNA__1027__D _1029_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1186_ input29/X _1509_/A _1186_/S vssd1 vssd1 vccd1 vccd1 _1186_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1043__C _1043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1324_ peripheralBus_data[3] _1602_/A _1336_/S vssd1 vssd1 vccd1 vccd1 _1325_/B sky130_fd_sc_hd__mux2_1
X_1255_ _1568_/A input28/X _1298_/S vssd1 vssd1 vccd1 vccd1 _1255_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1497__129 vssd1 vssd1 vccd1 vccd1 _1497__129/HI _1627_/A sky130_fd_sc_hd__conb_1
X_1441__73 vssd1 vssd1 vccd1 vccd1 _1441__73/HI _1555_/A sky130_fd_sc_hd__conb_1
XANTENNA__1188__A1 _1185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1040_ _1040_/A vssd1 vssd1 vccd1 vccd1 _1040_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0967__C _0972_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0824_ _0824_/A vssd1 vssd1 vccd1 vccd1 _0824_/X sky130_fd_sc_hd__clkbuf_1
X_0755_ _0755_/A _0755_/B vssd1 vssd1 vccd1 vccd1 _0756_/D sky130_fd_sc_hd__or2_1
XFILLER_29_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1169_ _1508_/A _1506_/A _1186_/S vssd1 vssd1 vccd1 vccd1 _1169_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1238_ _1348_/A _1238_/B vssd1 vssd1 vccd1 vccd1 _1376_/D sky130_fd_sc_hd__nor2_1
X_1307_ _1390_/Q _1305_/X _1307_/S vssd1 vssd1 vccd1 vccd1 _1307_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1023_ _1065_/A vssd1 vssd1 vccd1 vccd1 _1035_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0994__A _0994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0807_ _0807_/A vssd1 vssd1 vccd1 vccd1 _0807_/X sky130_fd_sc_hd__clkbuf_1
X_1411__43 vssd1 vssd1 vccd1 vccd1 _1411__43/HI _1517_/A sky130_fd_sc_hd__conb_1
X_0738_ _1258_/B vssd1 vssd1 vccd1 vccd1 _1353_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__1065__A _1065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1391__CLK _1404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1572_ _1572_/A _0925_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[5] sky130_fd_sc_hd__ebufn_8
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1006_ _1006_/A vssd1 vssd1 vccd1 vccd1 _1006_/X sky130_fd_sc_hd__clkbuf_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1215__A0 peripheralBus_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1624_ _1624_/A _0844_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[25] sky130_fd_sc_hd__ebufn_8
X_1555_ _1555_/A _1092_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[20] sky130_fd_sc_hd__ebufn_8
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1253__A _1267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1340_ _1401_/Q _1599_/A vssd1 vssd1 vccd1 vccd1 _1340_/X sky130_fd_sc_hd__or2_1
XFILLER_3_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1271_ _1297_/A vssd1 vssd1 vccd1 vccd1 _1295_/A sky130_fd_sc_hd__buf_2
X_0986_ _0986_/A vssd1 vssd1 vccd1 vccd1 _0986_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1538_ _1538_/A _1048_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[3] sky130_fd_sc_hd__ebufn_8
X_1607_ _1607_/A _0901_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[8] sky130_fd_sc_hd__ebufn_8
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0840_ _0845_/A _0845_/B _0840_/C _0845_/D vssd1 vssd1 vccd1 vccd1 _0841_/A sky130_fd_sc_hd__or4_1
X_0771_ _0775_/A _0775_/B _0789_/C _0775_/D vssd1 vssd1 vccd1 vccd1 _0772_/A sky130_fd_sc_hd__or4_1
XFILLER_52_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1323_ _1323_/A vssd1 vssd1 vccd1 vccd1 _1393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1254_ _1604_/A vssd1 vssd1 vccd1 vccd1 _1298_/S sky130_fd_sc_hd__clkbuf_2
X_1185_ peripheralBus_data[7] vssd1 vssd1 vccd1 vccd1 _1185_/X sky130_fd_sc_hd__buf_2
XFILLER_32_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1188__A2 _1144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0969_ _0977_/A _0977_/B _0972_/C _0969_/D vssd1 vssd1 vccd1 vccd1 _0970_/A sky130_fd_sc_hd__or4_1
XFILLER_47_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1480__112 vssd1 vssd1 vccd1 vccd1 _1480__112/HI _1610_/A sky130_fd_sc_hd__conb_1
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0967__D _0969_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0823_ _0823_/A _0823_/B _0840_/C _0845_/D vssd1 vssd1 vccd1 vccd1 _0824_/A sky130_fd_sc_hd__or4_1
X_0754_ _0754_/A _0754_/B input3/X input2/X vssd1 vssd1 vccd1 vccd1 _0756_/C sky130_fd_sc_hd__or4_1
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1306_ _1399_/Q _1400_/Q _1602_/A vssd1 vssd1 vccd1 vccd1 _1307_/S sky130_fd_sc_hd__mux2_1
XFILLER_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1168_ _1168_/A vssd1 vssd1 vccd1 vccd1 _1362_/D sky130_fd_sc_hd__clkbuf_1
X_1099_ _1105_/A _1105_/B _1099_/C _1099_/D vssd1 vssd1 vccd1 vccd1 _1100_/A sky130_fd_sc_hd__or4_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1237_ _1236_/A _1376_/Q _1539_/A _1236_/X vssd1 vssd1 vccd1 vccd1 _1238_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1261__A _1269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1022_ _1022_/A vssd1 vssd1 vccd1 vccd1 _1022_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1260__B2 _1145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0806_ _0808_/A _0808_/B _0808_/C _0813_/D vssd1 vssd1 vccd1 vccd1 _0807_/A sky130_fd_sc_hd__or4_1
X_0737_ _0737_/A _0737_/B _0737_/C _0737_/D vssd1 vssd1 vccd1 vccd1 _1258_/B sky130_fd_sc_hd__or4_4
XFILLER_44_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input25_A peripheralBus_oe vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1571_ _1571_/A _0923_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[4] sky130_fd_sc_hd__ebufn_8
XFILLER_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1005_ _1005_/A _1005_/B _1015_/C _1015_/D vssd1 vssd1 vccd1 vccd1 _1006_/A sky130_fd_sc_hd__or4_1
XFILLER_34_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput30 _1128_/Y vssd1 vssd1 vccd1 vccd1 peripheralBus_busy sky130_fd_sc_hd__buf_2
XFILLER_48_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1623_ _1623_/A _0841_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[24] sky130_fd_sc_hd__ebufn_8
X_1554_ _1554_/A _1090_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[19] sky130_fd_sc_hd__ebufn_8
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

