magic
tech sky130A
magscale 1 2
timestamp 1653580153
<< obsli1 >>
rect 1104 2159 118864 167569
<< obsm1 >>
rect 1026 1640 119494 167816
<< metal2 >>
rect 754 169200 810 170000
rect 2318 169200 2374 170000
rect 3882 169200 3938 170000
rect 5446 169200 5502 170000
rect 7010 169200 7066 170000
rect 8574 169200 8630 170000
rect 10138 169200 10194 170000
rect 11794 169200 11850 170000
rect 13358 169200 13414 170000
rect 14922 169200 14978 170000
rect 16486 169200 16542 170000
rect 18050 169200 18106 170000
rect 19614 169200 19670 170000
rect 21270 169200 21326 170000
rect 22834 169200 22890 170000
rect 24398 169200 24454 170000
rect 25962 169200 26018 170000
rect 27526 169200 27582 170000
rect 29090 169200 29146 170000
rect 30746 169200 30802 170000
rect 32310 169200 32366 170000
rect 33874 169200 33930 170000
rect 35438 169200 35494 170000
rect 37002 169200 37058 170000
rect 38566 169200 38622 170000
rect 40130 169200 40186 170000
rect 41786 169200 41842 170000
rect 43350 169200 43406 170000
rect 44914 169200 44970 170000
rect 46478 169200 46534 170000
rect 48042 169200 48098 170000
rect 49606 169200 49662 170000
rect 51262 169200 51318 170000
rect 52826 169200 52882 170000
rect 54390 169200 54446 170000
rect 55954 169200 56010 170000
rect 57518 169200 57574 170000
rect 59082 169200 59138 170000
rect 60738 169200 60794 170000
rect 62302 169200 62358 170000
rect 63866 169200 63922 170000
rect 65430 169200 65486 170000
rect 66994 169200 67050 170000
rect 68558 169200 68614 170000
rect 70122 169200 70178 170000
rect 71778 169200 71834 170000
rect 73342 169200 73398 170000
rect 74906 169200 74962 170000
rect 76470 169200 76526 170000
rect 78034 169200 78090 170000
rect 79598 169200 79654 170000
rect 81254 169200 81310 170000
rect 82818 169200 82874 170000
rect 84382 169200 84438 170000
rect 85946 169200 86002 170000
rect 87510 169200 87566 170000
rect 89074 169200 89130 170000
rect 90730 169200 90786 170000
rect 92294 169200 92350 170000
rect 93858 169200 93914 170000
rect 95422 169200 95478 170000
rect 96986 169200 97042 170000
rect 98550 169200 98606 170000
rect 100114 169200 100170 170000
rect 101770 169200 101826 170000
rect 103334 169200 103390 170000
rect 104898 169200 104954 170000
rect 106462 169200 106518 170000
rect 108026 169200 108082 170000
rect 109590 169200 109646 170000
rect 111246 169200 111302 170000
rect 112810 169200 112866 170000
rect 114374 169200 114430 170000
rect 115938 169200 115994 170000
rect 117502 169200 117558 170000
rect 119066 169200 119122 170000
rect 1030 0 1086 800
rect 3146 0 3202 800
rect 5262 0 5318 800
rect 7378 0 7434 800
rect 9586 0 9642 800
rect 11702 0 11758 800
rect 13818 0 13874 800
rect 16026 0 16082 800
rect 18142 0 18198 800
rect 20258 0 20314 800
rect 22374 0 22430 800
rect 24582 0 24638 800
rect 26698 0 26754 800
rect 28814 0 28870 800
rect 31022 0 31078 800
rect 33138 0 33194 800
rect 35254 0 35310 800
rect 37370 0 37426 800
rect 39578 0 39634 800
rect 41694 0 41750 800
rect 43810 0 43866 800
rect 46018 0 46074 800
rect 48134 0 48190 800
rect 50250 0 50306 800
rect 52366 0 52422 800
rect 54574 0 54630 800
rect 56690 0 56746 800
rect 58806 0 58862 800
rect 61014 0 61070 800
rect 63130 0 63186 800
rect 65246 0 65302 800
rect 67362 0 67418 800
rect 69570 0 69626 800
rect 71686 0 71742 800
rect 73802 0 73858 800
rect 76010 0 76066 800
rect 78126 0 78182 800
rect 80242 0 80298 800
rect 82358 0 82414 800
rect 84566 0 84622 800
rect 86682 0 86738 800
rect 88798 0 88854 800
rect 91006 0 91062 800
rect 93122 0 93178 800
rect 95238 0 95294 800
rect 97354 0 97410 800
rect 99562 0 99618 800
rect 101678 0 101734 800
rect 103794 0 103850 800
rect 106002 0 106058 800
rect 108118 0 108174 800
rect 110234 0 110290 800
rect 112350 0 112406 800
rect 114558 0 114614 800
rect 116674 0 116730 800
rect 118790 0 118846 800
<< obsm2 >>
rect 1032 169144 2262 169266
rect 2430 169144 3826 169266
rect 3994 169144 5390 169266
rect 5558 169144 6954 169266
rect 7122 169144 8518 169266
rect 8686 169144 10082 169266
rect 10250 169144 11738 169266
rect 11906 169144 13302 169266
rect 13470 169144 14866 169266
rect 15034 169144 16430 169266
rect 16598 169144 17994 169266
rect 18162 169144 19558 169266
rect 19726 169144 21214 169266
rect 21382 169144 22778 169266
rect 22946 169144 24342 169266
rect 24510 169144 25906 169266
rect 26074 169144 27470 169266
rect 27638 169144 29034 169266
rect 29202 169144 30690 169266
rect 30858 169144 32254 169266
rect 32422 169144 33818 169266
rect 33986 169144 35382 169266
rect 35550 169144 36946 169266
rect 37114 169144 38510 169266
rect 38678 169144 40074 169266
rect 40242 169144 41730 169266
rect 41898 169144 43294 169266
rect 43462 169144 44858 169266
rect 45026 169144 46422 169266
rect 46590 169144 47986 169266
rect 48154 169144 49550 169266
rect 49718 169144 51206 169266
rect 51374 169144 52770 169266
rect 52938 169144 54334 169266
rect 54502 169144 55898 169266
rect 56066 169144 57462 169266
rect 57630 169144 59026 169266
rect 59194 169144 60682 169266
rect 60850 169144 62246 169266
rect 62414 169144 63810 169266
rect 63978 169144 65374 169266
rect 65542 169144 66938 169266
rect 67106 169144 68502 169266
rect 68670 169144 70066 169266
rect 70234 169144 71722 169266
rect 71890 169144 73286 169266
rect 73454 169144 74850 169266
rect 75018 169144 76414 169266
rect 76582 169144 77978 169266
rect 78146 169144 79542 169266
rect 79710 169144 81198 169266
rect 81366 169144 82762 169266
rect 82930 169144 84326 169266
rect 84494 169144 85890 169266
rect 86058 169144 87454 169266
rect 87622 169144 89018 169266
rect 89186 169144 90674 169266
rect 90842 169144 92238 169266
rect 92406 169144 93802 169266
rect 93970 169144 95366 169266
rect 95534 169144 96930 169266
rect 97098 169144 98494 169266
rect 98662 169144 100058 169266
rect 100226 169144 101714 169266
rect 101882 169144 103278 169266
rect 103446 169144 104842 169266
rect 105010 169144 106406 169266
rect 106574 169144 107970 169266
rect 108138 169144 109534 169266
rect 109702 169144 111190 169266
rect 111358 169144 112754 169266
rect 112922 169144 114318 169266
rect 114486 169144 115882 169266
rect 116050 169144 117446 169266
rect 117614 169144 119010 169266
rect 119178 169144 119488 169266
rect 1032 856 119488 169144
rect 1142 800 3090 856
rect 3258 800 5206 856
rect 5374 800 7322 856
rect 7490 800 9530 856
rect 9698 800 11646 856
rect 11814 800 13762 856
rect 13930 800 15970 856
rect 16138 800 18086 856
rect 18254 800 20202 856
rect 20370 800 22318 856
rect 22486 800 24526 856
rect 24694 800 26642 856
rect 26810 800 28758 856
rect 28926 800 30966 856
rect 31134 800 33082 856
rect 33250 800 35198 856
rect 35366 800 37314 856
rect 37482 800 39522 856
rect 39690 800 41638 856
rect 41806 800 43754 856
rect 43922 800 45962 856
rect 46130 800 48078 856
rect 48246 800 50194 856
rect 50362 800 52310 856
rect 52478 800 54518 856
rect 54686 800 56634 856
rect 56802 800 58750 856
rect 58918 800 60958 856
rect 61126 800 63074 856
rect 63242 800 65190 856
rect 65358 800 67306 856
rect 67474 800 69514 856
rect 69682 800 71630 856
rect 71798 800 73746 856
rect 73914 800 75954 856
rect 76122 800 78070 856
rect 78238 800 80186 856
rect 80354 800 82302 856
rect 82470 800 84510 856
rect 84678 800 86626 856
rect 86794 800 88742 856
rect 88910 800 90950 856
rect 91118 800 93066 856
rect 93234 800 95182 856
rect 95350 800 97298 856
rect 97466 800 99506 856
rect 99674 800 101622 856
rect 101790 800 103738 856
rect 103906 800 105946 856
rect 106114 800 108062 856
rect 108230 800 110178 856
rect 110346 800 112294 856
rect 112462 800 114502 856
rect 114670 800 116618 856
rect 116786 800 118734 856
rect 118902 800 119488 856
<< metal3 >>
rect 0 169056 800 169176
rect 0 167424 800 167544
rect 0 165656 800 165776
rect 0 164024 800 164144
rect 0 162256 800 162376
rect 0 160624 800 160744
rect 0 158856 800 158976
rect 0 157224 800 157344
rect 119200 155728 120000 155848
rect 0 155456 800 155576
rect 0 153824 800 153944
rect 0 152056 800 152176
rect 0 150424 800 150544
rect 0 148656 800 148776
rect 0 147024 800 147144
rect 0 145256 800 145376
rect 0 143624 800 143744
rect 0 141856 800 141976
rect 0 140224 800 140344
rect 0 138456 800 138576
rect 0 136824 800 136944
rect 0 135056 800 135176
rect 0 133424 800 133544
rect 0 131656 800 131776
rect 0 130024 800 130144
rect 0 128256 800 128376
rect 119200 127440 120000 127560
rect 0 126624 800 126744
rect 0 124856 800 124976
rect 0 123224 800 123344
rect 0 121456 800 121576
rect 0 119824 800 119944
rect 0 118056 800 118176
rect 0 116424 800 116544
rect 0 114656 800 114776
rect 0 113024 800 113144
rect 0 111256 800 111376
rect 0 109624 800 109744
rect 0 107856 800 107976
rect 0 106224 800 106344
rect 0 104456 800 104576
rect 0 102824 800 102944
rect 0 101056 800 101176
rect 0 99424 800 99544
rect 119200 99152 120000 99272
rect 0 97656 800 97776
rect 0 96024 800 96144
rect 0 94256 800 94376
rect 0 92624 800 92744
rect 0 90856 800 90976
rect 0 89224 800 89344
rect 0 87456 800 87576
rect 0 85824 800 85944
rect 0 84056 800 84176
rect 0 82424 800 82544
rect 0 80656 800 80776
rect 0 79024 800 79144
rect 0 77256 800 77376
rect 0 75624 800 75744
rect 0 73856 800 73976
rect 0 72224 800 72344
rect 119200 70728 120000 70848
rect 0 70456 800 70576
rect 0 68824 800 68944
rect 0 67056 800 67176
rect 0 65424 800 65544
rect 0 63656 800 63776
rect 0 62024 800 62144
rect 0 60256 800 60376
rect 0 58624 800 58744
rect 0 56856 800 56976
rect 0 55224 800 55344
rect 0 53456 800 53576
rect 0 51824 800 51944
rect 0 50056 800 50176
rect 0 48424 800 48544
rect 0 46656 800 46776
rect 0 45024 800 45144
rect 0 43256 800 43376
rect 119200 42440 120000 42560
rect 0 41624 800 41744
rect 0 39856 800 39976
rect 0 38224 800 38344
rect 0 36456 800 36576
rect 0 34824 800 34944
rect 0 33056 800 33176
rect 0 31424 800 31544
rect 0 29656 800 29776
rect 0 28024 800 28144
rect 0 26256 800 26376
rect 0 24624 800 24744
rect 0 22856 800 22976
rect 0 21224 800 21344
rect 0 19456 800 19576
rect 0 17824 800 17944
rect 0 16056 800 16176
rect 0 14424 800 14544
rect 119200 14152 120000 14272
rect 0 12656 800 12776
rect 0 11024 800 11144
rect 0 9256 800 9376
rect 0 7624 800 7744
rect 0 5856 800 5976
rect 0 4224 800 4344
rect 0 2456 800 2576
rect 0 824 800 944
<< obsm3 >>
rect 880 168976 119200 169149
rect 800 167624 119200 168976
rect 880 167344 119200 167624
rect 800 165856 119200 167344
rect 880 165576 119200 165856
rect 800 164224 119200 165576
rect 880 163944 119200 164224
rect 800 162456 119200 163944
rect 880 162176 119200 162456
rect 800 160824 119200 162176
rect 880 160544 119200 160824
rect 800 159056 119200 160544
rect 880 158776 119200 159056
rect 800 157424 119200 158776
rect 880 157144 119200 157424
rect 800 155928 119200 157144
rect 800 155656 119120 155928
rect 880 155648 119120 155656
rect 880 155376 119200 155648
rect 800 154024 119200 155376
rect 880 153744 119200 154024
rect 800 152256 119200 153744
rect 880 151976 119200 152256
rect 800 150624 119200 151976
rect 880 150344 119200 150624
rect 800 148856 119200 150344
rect 880 148576 119200 148856
rect 800 147224 119200 148576
rect 880 146944 119200 147224
rect 800 145456 119200 146944
rect 880 145176 119200 145456
rect 800 143824 119200 145176
rect 880 143544 119200 143824
rect 800 142056 119200 143544
rect 880 141776 119200 142056
rect 800 140424 119200 141776
rect 880 140144 119200 140424
rect 800 138656 119200 140144
rect 880 138376 119200 138656
rect 800 137024 119200 138376
rect 880 136744 119200 137024
rect 800 135256 119200 136744
rect 880 134976 119200 135256
rect 800 133624 119200 134976
rect 880 133344 119200 133624
rect 800 131856 119200 133344
rect 880 131576 119200 131856
rect 800 130224 119200 131576
rect 880 129944 119200 130224
rect 800 128456 119200 129944
rect 880 128176 119200 128456
rect 800 127640 119200 128176
rect 800 127360 119120 127640
rect 800 126824 119200 127360
rect 880 126544 119200 126824
rect 800 125056 119200 126544
rect 880 124776 119200 125056
rect 800 123424 119200 124776
rect 880 123144 119200 123424
rect 800 121656 119200 123144
rect 880 121376 119200 121656
rect 800 120024 119200 121376
rect 880 119744 119200 120024
rect 800 118256 119200 119744
rect 880 117976 119200 118256
rect 800 116624 119200 117976
rect 880 116344 119200 116624
rect 800 114856 119200 116344
rect 880 114576 119200 114856
rect 800 113224 119200 114576
rect 880 112944 119200 113224
rect 800 111456 119200 112944
rect 880 111176 119200 111456
rect 800 109824 119200 111176
rect 880 109544 119200 109824
rect 800 108056 119200 109544
rect 880 107776 119200 108056
rect 800 106424 119200 107776
rect 880 106144 119200 106424
rect 800 104656 119200 106144
rect 880 104376 119200 104656
rect 800 103024 119200 104376
rect 880 102744 119200 103024
rect 800 101256 119200 102744
rect 880 100976 119200 101256
rect 800 99624 119200 100976
rect 880 99352 119200 99624
rect 880 99344 119120 99352
rect 800 99072 119120 99344
rect 800 97856 119200 99072
rect 880 97576 119200 97856
rect 800 96224 119200 97576
rect 880 95944 119200 96224
rect 800 94456 119200 95944
rect 880 94176 119200 94456
rect 800 92824 119200 94176
rect 880 92544 119200 92824
rect 800 91056 119200 92544
rect 880 90776 119200 91056
rect 800 89424 119200 90776
rect 880 89144 119200 89424
rect 800 87656 119200 89144
rect 880 87376 119200 87656
rect 800 86024 119200 87376
rect 880 85744 119200 86024
rect 800 84256 119200 85744
rect 880 83976 119200 84256
rect 800 82624 119200 83976
rect 880 82344 119200 82624
rect 800 80856 119200 82344
rect 880 80576 119200 80856
rect 800 79224 119200 80576
rect 880 78944 119200 79224
rect 800 77456 119200 78944
rect 880 77176 119200 77456
rect 800 75824 119200 77176
rect 880 75544 119200 75824
rect 800 74056 119200 75544
rect 880 73776 119200 74056
rect 800 72424 119200 73776
rect 880 72144 119200 72424
rect 800 70928 119200 72144
rect 800 70656 119120 70928
rect 880 70648 119120 70656
rect 880 70376 119200 70648
rect 800 69024 119200 70376
rect 880 68744 119200 69024
rect 800 67256 119200 68744
rect 880 66976 119200 67256
rect 800 65624 119200 66976
rect 880 65344 119200 65624
rect 800 63856 119200 65344
rect 880 63576 119200 63856
rect 800 62224 119200 63576
rect 880 61944 119200 62224
rect 800 60456 119200 61944
rect 880 60176 119200 60456
rect 800 58824 119200 60176
rect 880 58544 119200 58824
rect 800 57056 119200 58544
rect 880 56776 119200 57056
rect 800 55424 119200 56776
rect 880 55144 119200 55424
rect 800 53656 119200 55144
rect 880 53376 119200 53656
rect 800 52024 119200 53376
rect 880 51744 119200 52024
rect 800 50256 119200 51744
rect 880 49976 119200 50256
rect 800 48624 119200 49976
rect 880 48344 119200 48624
rect 800 46856 119200 48344
rect 880 46576 119200 46856
rect 800 45224 119200 46576
rect 880 44944 119200 45224
rect 800 43456 119200 44944
rect 880 43176 119200 43456
rect 800 42640 119200 43176
rect 800 42360 119120 42640
rect 800 41824 119200 42360
rect 880 41544 119200 41824
rect 800 40056 119200 41544
rect 880 39776 119200 40056
rect 800 38424 119200 39776
rect 880 38144 119200 38424
rect 800 36656 119200 38144
rect 880 36376 119200 36656
rect 800 35024 119200 36376
rect 880 34744 119200 35024
rect 800 33256 119200 34744
rect 880 32976 119200 33256
rect 800 31624 119200 32976
rect 880 31344 119200 31624
rect 800 29856 119200 31344
rect 880 29576 119200 29856
rect 800 28224 119200 29576
rect 880 27944 119200 28224
rect 800 26456 119200 27944
rect 880 26176 119200 26456
rect 800 24824 119200 26176
rect 880 24544 119200 24824
rect 800 23056 119200 24544
rect 880 22776 119200 23056
rect 800 21424 119200 22776
rect 880 21144 119200 21424
rect 800 19656 119200 21144
rect 880 19376 119200 19656
rect 800 18024 119200 19376
rect 880 17744 119200 18024
rect 800 16256 119200 17744
rect 880 15976 119200 16256
rect 800 14624 119200 15976
rect 880 14352 119200 14624
rect 880 14344 119120 14352
rect 800 14072 119120 14344
rect 800 12856 119200 14072
rect 880 12576 119200 12856
rect 800 11224 119200 12576
rect 880 10944 119200 11224
rect 800 9456 119200 10944
rect 880 9176 119200 9456
rect 800 7824 119200 9176
rect 880 7544 119200 7824
rect 800 6056 119200 7544
rect 880 5776 119200 6056
rect 800 4424 119200 5776
rect 880 4144 119200 4424
rect 800 2656 119200 4144
rect 880 2376 119200 2656
rect 800 1024 119200 2376
rect 880 851 119200 1024
<< metal4 >>
rect 4208 2128 4528 167600
rect 19568 2128 19888 167600
rect 34928 2128 35248 167600
rect 50288 2128 50608 167600
rect 65648 2128 65968 167600
rect 81008 2128 81328 167600
rect 96368 2128 96688 167600
rect 111728 2128 112048 167600
<< obsm4 >>
rect 9259 2483 19488 167109
rect 19968 2483 34848 167109
rect 35328 2483 50208 167109
rect 50688 2483 65568 167109
rect 66048 2483 80928 167109
rect 81408 2483 96288 167109
rect 96768 2483 111648 167109
rect 112128 2483 114757 167109
<< labels >>
rlabel metal2 s 86682 0 86738 800 6 flash_csb
port 1 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 flash_io0_read
port 2 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 flash_io0_we
port 3 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 flash_io0_write
port 4 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 flash_io1_read
port 5 nsew signal output
rlabel metal2 s 97354 0 97410 800 6 flash_io1_we
port 6 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 flash_io1_write
port 7 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 flash_sck
port 8 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 internal_uart_rx
port 9 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 internal_uart_tx
port 10 nsew signal output
rlabel metal2 s 754 169200 810 170000 6 io_in[0]
port 11 nsew signal input
rlabel metal2 s 16486 169200 16542 170000 6 io_in[10]
port 12 nsew signal input
rlabel metal2 s 18050 169200 18106 170000 6 io_in[11]
port 13 nsew signal input
rlabel metal2 s 19614 169200 19670 170000 6 io_in[12]
port 14 nsew signal input
rlabel metal2 s 21270 169200 21326 170000 6 io_in[13]
port 15 nsew signal input
rlabel metal2 s 22834 169200 22890 170000 6 io_in[14]
port 16 nsew signal input
rlabel metal2 s 24398 169200 24454 170000 6 io_in[15]
port 17 nsew signal input
rlabel metal2 s 25962 169200 26018 170000 6 io_in[16]
port 18 nsew signal input
rlabel metal2 s 27526 169200 27582 170000 6 io_in[17]
port 19 nsew signal input
rlabel metal2 s 29090 169200 29146 170000 6 io_in[18]
port 20 nsew signal input
rlabel metal2 s 30746 169200 30802 170000 6 io_in[19]
port 21 nsew signal input
rlabel metal2 s 2318 169200 2374 170000 6 io_in[1]
port 22 nsew signal input
rlabel metal2 s 32310 169200 32366 170000 6 io_in[20]
port 23 nsew signal input
rlabel metal2 s 33874 169200 33930 170000 6 io_in[21]
port 24 nsew signal input
rlabel metal2 s 35438 169200 35494 170000 6 io_in[22]
port 25 nsew signal input
rlabel metal2 s 37002 169200 37058 170000 6 io_in[23]
port 26 nsew signal input
rlabel metal2 s 38566 169200 38622 170000 6 io_in[24]
port 27 nsew signal input
rlabel metal2 s 40130 169200 40186 170000 6 io_in[25]
port 28 nsew signal input
rlabel metal2 s 41786 169200 41842 170000 6 io_in[26]
port 29 nsew signal input
rlabel metal2 s 43350 169200 43406 170000 6 io_in[27]
port 30 nsew signal input
rlabel metal2 s 44914 169200 44970 170000 6 io_in[28]
port 31 nsew signal input
rlabel metal2 s 46478 169200 46534 170000 6 io_in[29]
port 32 nsew signal input
rlabel metal2 s 3882 169200 3938 170000 6 io_in[2]
port 33 nsew signal input
rlabel metal2 s 48042 169200 48098 170000 6 io_in[30]
port 34 nsew signal input
rlabel metal2 s 49606 169200 49662 170000 6 io_in[31]
port 35 nsew signal input
rlabel metal2 s 51262 169200 51318 170000 6 io_in[32]
port 36 nsew signal input
rlabel metal2 s 52826 169200 52882 170000 6 io_in[33]
port 37 nsew signal input
rlabel metal2 s 54390 169200 54446 170000 6 io_in[34]
port 38 nsew signal input
rlabel metal2 s 55954 169200 56010 170000 6 io_in[35]
port 39 nsew signal input
rlabel metal2 s 57518 169200 57574 170000 6 io_in[36]
port 40 nsew signal input
rlabel metal2 s 59082 169200 59138 170000 6 io_in[37]
port 41 nsew signal input
rlabel metal2 s 5446 169200 5502 170000 6 io_in[3]
port 42 nsew signal input
rlabel metal2 s 7010 169200 7066 170000 6 io_in[4]
port 43 nsew signal input
rlabel metal2 s 8574 169200 8630 170000 6 io_in[5]
port 44 nsew signal input
rlabel metal2 s 10138 169200 10194 170000 6 io_in[6]
port 45 nsew signal input
rlabel metal2 s 11794 169200 11850 170000 6 io_in[7]
port 46 nsew signal input
rlabel metal2 s 13358 169200 13414 170000 6 io_in[8]
port 47 nsew signal input
rlabel metal2 s 14922 169200 14978 170000 6 io_in[9]
port 48 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 io_oeb[0]
port 49 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 io_oeb[10]
port 50 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 io_oeb[11]
port 51 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 io_oeb[12]
port 52 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 io_oeb[13]
port 53 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 io_oeb[14]
port 54 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 io_oeb[15]
port 55 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 io_oeb[16]
port 56 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 io_oeb[17]
port 57 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 io_oeb[18]
port 58 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 io_oeb[19]
port 59 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 io_oeb[1]
port 60 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 io_oeb[20]
port 61 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 io_oeb[21]
port 62 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 io_oeb[22]
port 63 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 io_oeb[23]
port 64 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 io_oeb[24]
port 65 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 io_oeb[25]
port 66 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 io_oeb[26]
port 67 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 io_oeb[27]
port 68 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 io_oeb[28]
port 69 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 io_oeb[29]
port 70 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 io_oeb[2]
port 71 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 io_oeb[30]
port 72 nsew signal output
rlabel metal2 s 67362 0 67418 800 6 io_oeb[31]
port 73 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 io_oeb[32]
port 74 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 io_oeb[33]
port 75 nsew signal output
rlabel metal2 s 73802 0 73858 800 6 io_oeb[34]
port 76 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 io_oeb[35]
port 77 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 io_oeb[36]
port 78 nsew signal output
rlabel metal2 s 80242 0 80298 800 6 io_oeb[37]
port 79 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 io_oeb[3]
port 80 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 io_oeb[4]
port 81 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 io_oeb[5]
port 82 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 io_oeb[6]
port 83 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 io_oeb[7]
port 84 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 io_oeb[8]
port 85 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 io_oeb[9]
port 86 nsew signal output
rlabel metal2 s 60738 169200 60794 170000 6 io_out[0]
port 87 nsew signal output
rlabel metal2 s 76470 169200 76526 170000 6 io_out[10]
port 88 nsew signal output
rlabel metal2 s 78034 169200 78090 170000 6 io_out[11]
port 89 nsew signal output
rlabel metal2 s 79598 169200 79654 170000 6 io_out[12]
port 90 nsew signal output
rlabel metal2 s 81254 169200 81310 170000 6 io_out[13]
port 91 nsew signal output
rlabel metal2 s 82818 169200 82874 170000 6 io_out[14]
port 92 nsew signal output
rlabel metal2 s 84382 169200 84438 170000 6 io_out[15]
port 93 nsew signal output
rlabel metal2 s 85946 169200 86002 170000 6 io_out[16]
port 94 nsew signal output
rlabel metal2 s 87510 169200 87566 170000 6 io_out[17]
port 95 nsew signal output
rlabel metal2 s 89074 169200 89130 170000 6 io_out[18]
port 96 nsew signal output
rlabel metal2 s 90730 169200 90786 170000 6 io_out[19]
port 97 nsew signal output
rlabel metal2 s 62302 169200 62358 170000 6 io_out[1]
port 98 nsew signal output
rlabel metal2 s 92294 169200 92350 170000 6 io_out[20]
port 99 nsew signal output
rlabel metal2 s 93858 169200 93914 170000 6 io_out[21]
port 100 nsew signal output
rlabel metal2 s 95422 169200 95478 170000 6 io_out[22]
port 101 nsew signal output
rlabel metal2 s 96986 169200 97042 170000 6 io_out[23]
port 102 nsew signal output
rlabel metal2 s 98550 169200 98606 170000 6 io_out[24]
port 103 nsew signal output
rlabel metal2 s 100114 169200 100170 170000 6 io_out[25]
port 104 nsew signal output
rlabel metal2 s 101770 169200 101826 170000 6 io_out[26]
port 105 nsew signal output
rlabel metal2 s 103334 169200 103390 170000 6 io_out[27]
port 106 nsew signal output
rlabel metal2 s 104898 169200 104954 170000 6 io_out[28]
port 107 nsew signal output
rlabel metal2 s 106462 169200 106518 170000 6 io_out[29]
port 108 nsew signal output
rlabel metal2 s 63866 169200 63922 170000 6 io_out[2]
port 109 nsew signal output
rlabel metal2 s 108026 169200 108082 170000 6 io_out[30]
port 110 nsew signal output
rlabel metal2 s 109590 169200 109646 170000 6 io_out[31]
port 111 nsew signal output
rlabel metal2 s 111246 169200 111302 170000 6 io_out[32]
port 112 nsew signal output
rlabel metal2 s 112810 169200 112866 170000 6 io_out[33]
port 113 nsew signal output
rlabel metal2 s 114374 169200 114430 170000 6 io_out[34]
port 114 nsew signal output
rlabel metal2 s 115938 169200 115994 170000 6 io_out[35]
port 115 nsew signal output
rlabel metal2 s 117502 169200 117558 170000 6 io_out[36]
port 116 nsew signal output
rlabel metal2 s 119066 169200 119122 170000 6 io_out[37]
port 117 nsew signal output
rlabel metal2 s 65430 169200 65486 170000 6 io_out[3]
port 118 nsew signal output
rlabel metal2 s 66994 169200 67050 170000 6 io_out[4]
port 119 nsew signal output
rlabel metal2 s 68558 169200 68614 170000 6 io_out[5]
port 120 nsew signal output
rlabel metal2 s 70122 169200 70178 170000 6 io_out[6]
port 121 nsew signal output
rlabel metal2 s 71778 169200 71834 170000 6 io_out[7]
port 122 nsew signal output
rlabel metal2 s 73342 169200 73398 170000 6 io_out[8]
port 123 nsew signal output
rlabel metal2 s 74906 169200 74962 170000 6 io_out[9]
port 124 nsew signal output
rlabel metal3 s 119200 70728 120000 70848 6 jtag_tck
port 125 nsew signal output
rlabel metal3 s 119200 99152 120000 99272 6 jtag_tdi
port 126 nsew signal output
rlabel metal3 s 119200 127440 120000 127560 6 jtag_tdo
port 127 nsew signal input
rlabel metal3 s 119200 155728 120000 155848 6 jtag_tms
port 128 nsew signal output
rlabel metal3 s 119200 14152 120000 14272 6 probe_blink[0]
port 129 nsew signal output
rlabel metal3 s 119200 42440 120000 42560 6 probe_blink[1]
port 130 nsew signal output
rlabel metal4 s 4208 2128 4528 167600 6 vccd1
port 131 nsew power input
rlabel metal4 s 34928 2128 35248 167600 6 vccd1
port 131 nsew power input
rlabel metal4 s 65648 2128 65968 167600 6 vccd1
port 131 nsew power input
rlabel metal4 s 96368 2128 96688 167600 6 vccd1
port 131 nsew power input
rlabel metal2 s 108118 0 108174 800 6 vga_b[0]
port 132 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 vga_b[1]
port 133 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 vga_g[0]
port 134 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 vga_g[1]
port 135 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 vga_hsync
port 136 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 vga_r[0]
port 137 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 vga_r[1]
port 138 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 vga_vsync
port 139 nsew signal input
rlabel metal4 s 19568 2128 19888 167600 6 vssd1
port 140 nsew ground input
rlabel metal4 s 50288 2128 50608 167600 6 vssd1
port 140 nsew ground input
rlabel metal4 s 81008 2128 81328 167600 6 vssd1
port 140 nsew ground input
rlabel metal4 s 111728 2128 112048 167600 6 vssd1
port 140 nsew ground input
rlabel metal3 s 0 824 800 944 6 wb_ack_o
port 141 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 wb_adr_i[0]
port 142 nsew signal input
rlabel metal3 s 0 72224 800 72344 6 wb_adr_i[10]
port 143 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 wb_adr_i[11]
port 144 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 wb_adr_i[12]
port 145 nsew signal input
rlabel metal3 s 0 87456 800 87576 6 wb_adr_i[13]
port 146 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 wb_adr_i[14]
port 147 nsew signal input
rlabel metal3 s 0 97656 800 97776 6 wb_adr_i[15]
port 148 nsew signal input
rlabel metal3 s 0 102824 800 102944 6 wb_adr_i[16]
port 149 nsew signal input
rlabel metal3 s 0 107856 800 107976 6 wb_adr_i[17]
port 150 nsew signal input
rlabel metal3 s 0 113024 800 113144 6 wb_adr_i[18]
port 151 nsew signal input
rlabel metal3 s 0 118056 800 118176 6 wb_adr_i[19]
port 152 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 wb_adr_i[1]
port 153 nsew signal input
rlabel metal3 s 0 123224 800 123344 6 wb_adr_i[20]
port 154 nsew signal input
rlabel metal3 s 0 128256 800 128376 6 wb_adr_i[21]
port 155 nsew signal input
rlabel metal3 s 0 133424 800 133544 6 wb_adr_i[22]
port 156 nsew signal input
rlabel metal3 s 0 138456 800 138576 6 wb_adr_i[23]
port 157 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 wb_adr_i[2]
port 158 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 wb_adr_i[3]
port 159 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 wb_adr_i[4]
port 160 nsew signal input
rlabel metal3 s 0 46656 800 46776 6 wb_adr_i[5]
port 161 nsew signal input
rlabel metal3 s 0 51824 800 51944 6 wb_adr_i[6]
port 162 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 wb_adr_i[7]
port 163 nsew signal input
rlabel metal3 s 0 62024 800 62144 6 wb_adr_i[8]
port 164 nsew signal input
rlabel metal3 s 0 67056 800 67176 6 wb_adr_i[9]
port 165 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 wb_clk_i
port 166 nsew signal input
rlabel metal3 s 0 4224 800 4344 6 wb_cyc_i
port 167 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 wb_data_i[0]
port 168 nsew signal input
rlabel metal3 s 0 73856 800 73976 6 wb_data_i[10]
port 169 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 wb_data_i[11]
port 170 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 wb_data_i[12]
port 171 nsew signal input
rlabel metal3 s 0 89224 800 89344 6 wb_data_i[13]
port 172 nsew signal input
rlabel metal3 s 0 94256 800 94376 6 wb_data_i[14]
port 173 nsew signal input
rlabel metal3 s 0 99424 800 99544 6 wb_data_i[15]
port 174 nsew signal input
rlabel metal3 s 0 104456 800 104576 6 wb_data_i[16]
port 175 nsew signal input
rlabel metal3 s 0 109624 800 109744 6 wb_data_i[17]
port 176 nsew signal input
rlabel metal3 s 0 114656 800 114776 6 wb_data_i[18]
port 177 nsew signal input
rlabel metal3 s 0 119824 800 119944 6 wb_data_i[19]
port 178 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 wb_data_i[1]
port 179 nsew signal input
rlabel metal3 s 0 124856 800 124976 6 wb_data_i[20]
port 180 nsew signal input
rlabel metal3 s 0 130024 800 130144 6 wb_data_i[21]
port 181 nsew signal input
rlabel metal3 s 0 135056 800 135176 6 wb_data_i[22]
port 182 nsew signal input
rlabel metal3 s 0 140224 800 140344 6 wb_data_i[23]
port 183 nsew signal input
rlabel metal3 s 0 143624 800 143744 6 wb_data_i[24]
port 184 nsew signal input
rlabel metal3 s 0 147024 800 147144 6 wb_data_i[25]
port 185 nsew signal input
rlabel metal3 s 0 150424 800 150544 6 wb_data_i[26]
port 186 nsew signal input
rlabel metal3 s 0 153824 800 153944 6 wb_data_i[27]
port 187 nsew signal input
rlabel metal3 s 0 157224 800 157344 6 wb_data_i[28]
port 188 nsew signal input
rlabel metal3 s 0 160624 800 160744 6 wb_data_i[29]
port 189 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 wb_data_i[2]
port 190 nsew signal input
rlabel metal3 s 0 164024 800 164144 6 wb_data_i[30]
port 191 nsew signal input
rlabel metal3 s 0 167424 800 167544 6 wb_data_i[31]
port 192 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 wb_data_i[3]
port 193 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 wb_data_i[4]
port 194 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 wb_data_i[5]
port 195 nsew signal input
rlabel metal3 s 0 53456 800 53576 6 wb_data_i[6]
port 196 nsew signal input
rlabel metal3 s 0 58624 800 58744 6 wb_data_i[7]
port 197 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 wb_data_i[8]
port 198 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 wb_data_i[9]
port 199 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 wb_data_o[0]
port 200 nsew signal output
rlabel metal3 s 0 75624 800 75744 6 wb_data_o[10]
port 201 nsew signal output
rlabel metal3 s 0 80656 800 80776 6 wb_data_o[11]
port 202 nsew signal output
rlabel metal3 s 0 85824 800 85944 6 wb_data_o[12]
port 203 nsew signal output
rlabel metal3 s 0 90856 800 90976 6 wb_data_o[13]
port 204 nsew signal output
rlabel metal3 s 0 96024 800 96144 6 wb_data_o[14]
port 205 nsew signal output
rlabel metal3 s 0 101056 800 101176 6 wb_data_o[15]
port 206 nsew signal output
rlabel metal3 s 0 106224 800 106344 6 wb_data_o[16]
port 207 nsew signal output
rlabel metal3 s 0 111256 800 111376 6 wb_data_o[17]
port 208 nsew signal output
rlabel metal3 s 0 116424 800 116544 6 wb_data_o[18]
port 209 nsew signal output
rlabel metal3 s 0 121456 800 121576 6 wb_data_o[19]
port 210 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 wb_data_o[1]
port 211 nsew signal output
rlabel metal3 s 0 126624 800 126744 6 wb_data_o[20]
port 212 nsew signal output
rlabel metal3 s 0 131656 800 131776 6 wb_data_o[21]
port 213 nsew signal output
rlabel metal3 s 0 136824 800 136944 6 wb_data_o[22]
port 214 nsew signal output
rlabel metal3 s 0 141856 800 141976 6 wb_data_o[23]
port 215 nsew signal output
rlabel metal3 s 0 145256 800 145376 6 wb_data_o[24]
port 216 nsew signal output
rlabel metal3 s 0 148656 800 148776 6 wb_data_o[25]
port 217 nsew signal output
rlabel metal3 s 0 152056 800 152176 6 wb_data_o[26]
port 218 nsew signal output
rlabel metal3 s 0 155456 800 155576 6 wb_data_o[27]
port 219 nsew signal output
rlabel metal3 s 0 158856 800 158976 6 wb_data_o[28]
port 220 nsew signal output
rlabel metal3 s 0 162256 800 162376 6 wb_data_o[29]
port 221 nsew signal output
rlabel metal3 s 0 31424 800 31544 6 wb_data_o[2]
port 222 nsew signal output
rlabel metal3 s 0 165656 800 165776 6 wb_data_o[30]
port 223 nsew signal output
rlabel metal3 s 0 169056 800 169176 6 wb_data_o[31]
port 224 nsew signal output
rlabel metal3 s 0 38224 800 38344 6 wb_data_o[3]
port 225 nsew signal output
rlabel metal3 s 0 45024 800 45144 6 wb_data_o[4]
port 226 nsew signal output
rlabel metal3 s 0 50056 800 50176 6 wb_data_o[5]
port 227 nsew signal output
rlabel metal3 s 0 55224 800 55344 6 wb_data_o[6]
port 228 nsew signal output
rlabel metal3 s 0 60256 800 60376 6 wb_data_o[7]
port 229 nsew signal output
rlabel metal3 s 0 65424 800 65544 6 wb_data_o[8]
port 230 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 wb_data_o[9]
port 231 nsew signal output
rlabel metal3 s 0 5856 800 5976 6 wb_error_o
port 232 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 wb_rst_i
port 233 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 wb_sel_i[0]
port 234 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 wb_sel_i[1]
port 235 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 wb_sel_i[2]
port 236 nsew signal input
rlabel metal3 s 0 39856 800 39976 6 wb_sel_i[3]
port 237 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 wb_stall_o
port 238 nsew signal output
rlabel metal3 s 0 11024 800 11144 6 wb_stb_i
port 239 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 wb_we_i
port 240 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 170000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 54105656
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripherals_Flat/runs/Peripherals_Flat/results/finishing/Peripherals.magic.gds
string GDS_START 1109524
<< end >>

