VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Peripherals
  CLASS BLOCK ;
  FOREIGN Peripherals ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 700.000 ;
  PIN flash_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END flash_csb
  PIN flash_io0_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END flash_io0_read
  PIN flash_io0_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END flash_io0_we
  PIN flash_io0_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END flash_io0_write
  PIN flash_io1_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END flash_io1_read
  PIN flash_io1_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END flash_io1_we
  PIN flash_io1_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END flash_io1_write
  PIN flash_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END flash_sck
  PIN internal_uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END internal_uart_rx
  PIN internal_uart_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END internal_uart_tx
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 696.000 2.210 700.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 696.000 133.770 700.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 696.000 146.650 700.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 696.000 159.990 700.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 696.000 172.870 700.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 696.000 186.210 700.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 696.000 199.550 700.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 696.000 212.430 700.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 696.000 225.770 700.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 696.000 238.650 700.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 696.000 251.990 700.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 696.000 15.090 700.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 696.000 265.330 700.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 696.000 278.210 700.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 696.000 291.550 700.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 696.000 304.430 700.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 696.000 317.770 700.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 696.000 331.110 700.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 696.000 343.990 700.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 696.000 357.330 700.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 696.000 370.210 700.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 696.000 383.550 700.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 696.000 28.430 700.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 696.000 396.890 700.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 696.000 409.770 700.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 696.000 423.110 700.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 696.000 435.990 700.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 696.000 449.330 700.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 696.000 462.670 700.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 696.000 475.550 700.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 696.000 488.890 700.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 696.000 41.310 700.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 696.000 54.650 700.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 696.000 67.990 700.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 696.000 80.870 700.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 696.000 94.210 700.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 696.000 107.090 700.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 696.000 120.430 700.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 696.000 6.350 700.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 696.000 137.910 700.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 696.000 151.250 700.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 696.000 164.130 700.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 696.000 177.470 700.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 696.000 190.810 700.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 696.000 203.690 700.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 696.000 217.030 700.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 696.000 229.910 700.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 696.000 243.250 700.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 696.000 256.590 700.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 696.000 19.690 700.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 696.000 269.470 700.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 696.000 282.810 700.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 696.000 295.690 700.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 696.000 309.030 700.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 696.000 322.370 700.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 696.000 335.250 700.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 696.000 348.590 700.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 696.000 361.470 700.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 696.000 374.810 700.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 696.000 388.150 700.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 696.000 32.570 700.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 696.000 401.030 700.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 696.000 414.370 700.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 696.000 427.250 700.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 696.000 440.590 700.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 696.000 453.930 700.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 696.000 466.810 700.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 696.000 480.150 700.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 696.000 493.030 700.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 696.000 45.910 700.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 696.000 58.790 700.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 696.000 72.130 700.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 696.000 85.470 700.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 696.000 98.350 700.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 696.000 111.690 700.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 696.000 124.570 700.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 696.000 10.950 700.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 696.000 142.510 700.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 696.000 155.390 700.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 696.000 168.730 700.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 696.000 181.610 700.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 696.000 194.950 700.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 696.000 208.290 700.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 696.000 221.170 700.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 696.000 234.510 700.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 696.000 247.390 700.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 696.000 260.730 700.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 696.000 23.830 700.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 696.000 274.070 700.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 696.000 286.950 700.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 696.000 300.290 700.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 696.000 313.170 700.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 696.000 326.510 700.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 696.000 339.850 700.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 696.000 352.730 700.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 696.000 366.070 700.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 696.000 379.410 700.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 696.000 392.290 700.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 696.000 37.170 700.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 696.000 405.630 700.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 696.000 418.510 700.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 696.000 431.850 700.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 696.000 445.190 700.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 696.000 458.070 700.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 696.000 471.410 700.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 696.000 484.290 700.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 696.000 497.630 700.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 696.000 50.050 700.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 696.000 63.390 700.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 696.000 76.730 700.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 696.000 89.610 700.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 696.000 102.950 700.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 696.000 115.830 700.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 696.000 129.170 700.000 ;
    END
  END io_out[9]
  PIN irq_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END irq_en
  PIN irq_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END irq_in
  PIN jtag_tck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END jtag_tms
  PIN probe_blink[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 174.800 500.000 175.400 ;
    END
  END probe_blink[0]
  PIN probe_blink[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 524.320 500.000 524.920 ;
    END
  END probe_blink[1]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 688.400 ;
    END
  END vccd1
  PIN vga_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END vga_b[0]
  PIN vga_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END vga_b[1]
  PIN vga_g[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END vga_g[0]
  PIN vga_g[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END vga_g[1]
  PIN vga_hsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END vga_hsync
  PIN vga_r[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END vga_r[0]
  PIN vga_r[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END vga_r[1]
  PIN vga_vsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END vga_vsync
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 688.400 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.800 4.000 549.400 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END wb_cyc_i
  PIN wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END wb_data_i[0]
  PIN wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END wb_data_i[10]
  PIN wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END wb_data_i[11]
  PIN wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END wb_data_i[12]
  PIN wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END wb_data_i[13]
  PIN wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END wb_data_i[14]
  PIN wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.720 4.000 409.320 ;
    END
  END wb_data_i[15]
  PIN wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END wb_data_i[16]
  PIN wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.880 4.000 451.480 ;
    END
  END wb_data_i[17]
  PIN wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END wb_data_i[18]
  PIN wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END wb_data_i[19]
  PIN wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END wb_data_i[1]
  PIN wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END wb_data_i[20]
  PIN wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END wb_data_i[21]
  PIN wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 555.600 4.000 556.200 ;
    END
  END wb_data_i[22]
  PIN wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.680 4.000 577.280 ;
    END
  END wb_data_i[23]
  PIN wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.960 4.000 591.560 ;
    END
  END wb_data_i[24]
  PIN wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 604.560 4.000 605.160 ;
    END
  END wb_data_i[25]
  PIN wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END wb_data_i[26]
  PIN wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.120 4.000 633.720 ;
    END
  END wb_data_i[27]
  PIN wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END wb_data_i[28]
  PIN wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END wb_data_i[29]
  PIN wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END wb_data_i[2]
  PIN wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END wb_data_i[30]
  PIN wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.880 4.000 689.480 ;
    END
  END wb_data_i[31]
  PIN wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END wb_data_i[3]
  PIN wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END wb_data_i[4]
  PIN wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END wb_data_i[5]
  PIN wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END wb_data_i[6]
  PIN wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END wb_data_i[7]
  PIN wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END wb_data_i[8]
  PIN wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END wb_data_i[9]
  PIN wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END wb_data_o[0]
  PIN wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END wb_data_o[10]
  PIN wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END wb_data_o[11]
  PIN wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END wb_data_o[12]
  PIN wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END wb_data_o[13]
  PIN wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END wb_data_o[14]
  PIN wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END wb_data_o[15]
  PIN wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END wb_data_o[16]
  PIN wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END wb_data_o[17]
  PIN wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END wb_data_o[18]
  PIN wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END wb_data_o[19]
  PIN wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END wb_data_o[1]
  PIN wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END wb_data_o[20]
  PIN wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.000 4.000 542.600 ;
    END
  END wb_data_o[21]
  PIN wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END wb_data_o[22]
  PIN wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.160 4.000 584.760 ;
    END
  END wb_data_o[23]
  PIN wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.760 4.000 598.360 ;
    END
  END wb_data_o[24]
  PIN wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END wb_data_o[25]
  PIN wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END wb_data_o[26]
  PIN wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.920 4.000 640.520 ;
    END
  END wb_data_o[27]
  PIN wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 653.520 4.000 654.120 ;
    END
  END wb_data_o[28]
  PIN wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END wb_data_o[29]
  PIN wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END wb_data_o[2]
  PIN wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.080 4.000 682.680 ;
    END
  END wb_data_o[30]
  PIN wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.680 4.000 696.280 ;
    END
  END wb_data_o[31]
  PIN wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END wb_data_o[3]
  PIN wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END wb_data_o[4]
  PIN wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END wb_data_o[5]
  PIN wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END wb_data_o[6]
  PIN wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END wb_data_o[7]
  PIN wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END wb_data_o[8]
  PIN wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END wb_data_o[9]
  PIN wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END wb_error_o
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END wb_sel_i[3]
  PIN wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END wb_stall_o
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 688.245 ;
      LAYER met1 ;
        RECT 5.520 10.640 497.650 688.400 ;
      LAYER met2 ;
        RECT 6.630 695.720 10.390 696.730 ;
        RECT 11.230 695.720 14.530 696.730 ;
        RECT 15.370 695.720 19.130 696.730 ;
        RECT 19.970 695.720 23.270 696.730 ;
        RECT 24.110 695.720 27.870 696.730 ;
        RECT 28.710 695.720 32.010 696.730 ;
        RECT 32.850 695.720 36.610 696.730 ;
        RECT 37.450 695.720 40.750 696.730 ;
        RECT 41.590 695.720 45.350 696.730 ;
        RECT 46.190 695.720 49.490 696.730 ;
        RECT 50.330 695.720 54.090 696.730 ;
        RECT 54.930 695.720 58.230 696.730 ;
        RECT 59.070 695.720 62.830 696.730 ;
        RECT 63.670 695.720 67.430 696.730 ;
        RECT 68.270 695.720 71.570 696.730 ;
        RECT 72.410 695.720 76.170 696.730 ;
        RECT 77.010 695.720 80.310 696.730 ;
        RECT 81.150 695.720 84.910 696.730 ;
        RECT 85.750 695.720 89.050 696.730 ;
        RECT 89.890 695.720 93.650 696.730 ;
        RECT 94.490 695.720 97.790 696.730 ;
        RECT 98.630 695.720 102.390 696.730 ;
        RECT 103.230 695.720 106.530 696.730 ;
        RECT 107.370 695.720 111.130 696.730 ;
        RECT 111.970 695.720 115.270 696.730 ;
        RECT 116.110 695.720 119.870 696.730 ;
        RECT 120.710 695.720 124.010 696.730 ;
        RECT 124.850 695.720 128.610 696.730 ;
        RECT 129.450 695.720 133.210 696.730 ;
        RECT 134.050 695.720 137.350 696.730 ;
        RECT 138.190 695.720 141.950 696.730 ;
        RECT 142.790 695.720 146.090 696.730 ;
        RECT 146.930 695.720 150.690 696.730 ;
        RECT 151.530 695.720 154.830 696.730 ;
        RECT 155.670 695.720 159.430 696.730 ;
        RECT 160.270 695.720 163.570 696.730 ;
        RECT 164.410 695.720 168.170 696.730 ;
        RECT 169.010 695.720 172.310 696.730 ;
        RECT 173.150 695.720 176.910 696.730 ;
        RECT 177.750 695.720 181.050 696.730 ;
        RECT 181.890 695.720 185.650 696.730 ;
        RECT 186.490 695.720 190.250 696.730 ;
        RECT 191.090 695.720 194.390 696.730 ;
        RECT 195.230 695.720 198.990 696.730 ;
        RECT 199.830 695.720 203.130 696.730 ;
        RECT 203.970 695.720 207.730 696.730 ;
        RECT 208.570 695.720 211.870 696.730 ;
        RECT 212.710 695.720 216.470 696.730 ;
        RECT 217.310 695.720 220.610 696.730 ;
        RECT 221.450 695.720 225.210 696.730 ;
        RECT 226.050 695.720 229.350 696.730 ;
        RECT 230.190 695.720 233.950 696.730 ;
        RECT 234.790 695.720 238.090 696.730 ;
        RECT 238.930 695.720 242.690 696.730 ;
        RECT 243.530 695.720 246.830 696.730 ;
        RECT 247.670 695.720 251.430 696.730 ;
        RECT 252.270 695.720 256.030 696.730 ;
        RECT 256.870 695.720 260.170 696.730 ;
        RECT 261.010 695.720 264.770 696.730 ;
        RECT 265.610 695.720 268.910 696.730 ;
        RECT 269.750 695.720 273.510 696.730 ;
        RECT 274.350 695.720 277.650 696.730 ;
        RECT 278.490 695.720 282.250 696.730 ;
        RECT 283.090 695.720 286.390 696.730 ;
        RECT 287.230 695.720 290.990 696.730 ;
        RECT 291.830 695.720 295.130 696.730 ;
        RECT 295.970 695.720 299.730 696.730 ;
        RECT 300.570 695.720 303.870 696.730 ;
        RECT 304.710 695.720 308.470 696.730 ;
        RECT 309.310 695.720 312.610 696.730 ;
        RECT 313.450 695.720 317.210 696.730 ;
        RECT 318.050 695.720 321.810 696.730 ;
        RECT 322.650 695.720 325.950 696.730 ;
        RECT 326.790 695.720 330.550 696.730 ;
        RECT 331.390 695.720 334.690 696.730 ;
        RECT 335.530 695.720 339.290 696.730 ;
        RECT 340.130 695.720 343.430 696.730 ;
        RECT 344.270 695.720 348.030 696.730 ;
        RECT 348.870 695.720 352.170 696.730 ;
        RECT 353.010 695.720 356.770 696.730 ;
        RECT 357.610 695.720 360.910 696.730 ;
        RECT 361.750 695.720 365.510 696.730 ;
        RECT 366.350 695.720 369.650 696.730 ;
        RECT 370.490 695.720 374.250 696.730 ;
        RECT 375.090 695.720 378.850 696.730 ;
        RECT 379.690 695.720 382.990 696.730 ;
        RECT 383.830 695.720 387.590 696.730 ;
        RECT 388.430 695.720 391.730 696.730 ;
        RECT 392.570 695.720 396.330 696.730 ;
        RECT 397.170 695.720 400.470 696.730 ;
        RECT 401.310 695.720 405.070 696.730 ;
        RECT 405.910 695.720 409.210 696.730 ;
        RECT 410.050 695.720 413.810 696.730 ;
        RECT 414.650 695.720 417.950 696.730 ;
        RECT 418.790 695.720 422.550 696.730 ;
        RECT 423.390 695.720 426.690 696.730 ;
        RECT 427.530 695.720 431.290 696.730 ;
        RECT 432.130 695.720 435.430 696.730 ;
        RECT 436.270 695.720 440.030 696.730 ;
        RECT 440.870 695.720 444.630 696.730 ;
        RECT 445.470 695.720 448.770 696.730 ;
        RECT 449.610 695.720 453.370 696.730 ;
        RECT 454.210 695.720 457.510 696.730 ;
        RECT 458.350 695.720 462.110 696.730 ;
        RECT 462.950 695.720 466.250 696.730 ;
        RECT 467.090 695.720 470.850 696.730 ;
        RECT 471.690 695.720 474.990 696.730 ;
        RECT 475.830 695.720 479.590 696.730 ;
        RECT 480.430 695.720 483.730 696.730 ;
        RECT 484.570 695.720 488.330 696.730 ;
        RECT 489.170 695.720 492.470 696.730 ;
        RECT 493.310 695.720 497.070 696.730 ;
        RECT 6.080 4.280 497.620 695.720 ;
        RECT 6.080 3.555 9.930 4.280 ;
        RECT 10.770 3.555 30.630 4.280 ;
        RECT 31.470 3.555 51.330 4.280 ;
        RECT 52.170 3.555 72.030 4.280 ;
        RECT 72.870 3.555 93.190 4.280 ;
        RECT 94.030 3.555 113.890 4.280 ;
        RECT 114.730 3.555 134.590 4.280 ;
        RECT 135.430 3.555 155.750 4.280 ;
        RECT 156.590 3.555 176.450 4.280 ;
        RECT 177.290 3.555 197.150 4.280 ;
        RECT 197.990 3.555 217.850 4.280 ;
        RECT 218.690 3.555 239.010 4.280 ;
        RECT 239.850 3.555 259.710 4.280 ;
        RECT 260.550 3.555 280.410 4.280 ;
        RECT 281.250 3.555 301.570 4.280 ;
        RECT 302.410 3.555 322.270 4.280 ;
        RECT 323.110 3.555 342.970 4.280 ;
        RECT 343.810 3.555 363.670 4.280 ;
        RECT 364.510 3.555 384.830 4.280 ;
        RECT 385.670 3.555 405.530 4.280 ;
        RECT 406.370 3.555 426.230 4.280 ;
        RECT 427.070 3.555 447.390 4.280 ;
        RECT 448.230 3.555 468.090 4.280 ;
        RECT 468.930 3.555 488.790 4.280 ;
        RECT 489.630 3.555 497.620 4.280 ;
      LAYER met3 ;
        RECT 4.400 695.280 496.000 696.145 ;
        RECT 4.000 689.880 496.000 695.280 ;
        RECT 4.400 688.480 496.000 689.880 ;
        RECT 4.000 683.080 496.000 688.480 ;
        RECT 4.400 681.680 496.000 683.080 ;
        RECT 4.000 675.600 496.000 681.680 ;
        RECT 4.400 674.200 496.000 675.600 ;
        RECT 4.000 668.800 496.000 674.200 ;
        RECT 4.400 667.400 496.000 668.800 ;
        RECT 4.000 662.000 496.000 667.400 ;
        RECT 4.400 660.600 496.000 662.000 ;
        RECT 4.000 654.520 496.000 660.600 ;
        RECT 4.400 653.120 496.000 654.520 ;
        RECT 4.000 647.720 496.000 653.120 ;
        RECT 4.400 646.320 496.000 647.720 ;
        RECT 4.000 640.920 496.000 646.320 ;
        RECT 4.400 639.520 496.000 640.920 ;
        RECT 4.000 634.120 496.000 639.520 ;
        RECT 4.400 632.720 496.000 634.120 ;
        RECT 4.000 626.640 496.000 632.720 ;
        RECT 4.400 625.240 496.000 626.640 ;
        RECT 4.000 619.840 496.000 625.240 ;
        RECT 4.400 618.440 496.000 619.840 ;
        RECT 4.000 613.040 496.000 618.440 ;
        RECT 4.400 611.640 496.000 613.040 ;
        RECT 4.000 605.560 496.000 611.640 ;
        RECT 4.400 604.160 496.000 605.560 ;
        RECT 4.000 598.760 496.000 604.160 ;
        RECT 4.400 597.360 496.000 598.760 ;
        RECT 4.000 591.960 496.000 597.360 ;
        RECT 4.400 590.560 496.000 591.960 ;
        RECT 4.000 585.160 496.000 590.560 ;
        RECT 4.400 583.760 496.000 585.160 ;
        RECT 4.000 577.680 496.000 583.760 ;
        RECT 4.400 576.280 496.000 577.680 ;
        RECT 4.000 570.880 496.000 576.280 ;
        RECT 4.400 569.480 496.000 570.880 ;
        RECT 4.000 564.080 496.000 569.480 ;
        RECT 4.400 562.680 496.000 564.080 ;
        RECT 4.000 556.600 496.000 562.680 ;
        RECT 4.400 555.200 496.000 556.600 ;
        RECT 4.000 549.800 496.000 555.200 ;
        RECT 4.400 548.400 496.000 549.800 ;
        RECT 4.000 543.000 496.000 548.400 ;
        RECT 4.400 541.600 496.000 543.000 ;
        RECT 4.000 536.200 496.000 541.600 ;
        RECT 4.400 534.800 496.000 536.200 ;
        RECT 4.000 528.720 496.000 534.800 ;
        RECT 4.400 527.320 496.000 528.720 ;
        RECT 4.000 525.320 496.000 527.320 ;
        RECT 4.000 523.920 495.600 525.320 ;
        RECT 4.000 521.920 496.000 523.920 ;
        RECT 4.400 520.520 496.000 521.920 ;
        RECT 4.000 515.120 496.000 520.520 ;
        RECT 4.400 513.720 496.000 515.120 ;
        RECT 4.000 507.640 496.000 513.720 ;
        RECT 4.400 506.240 496.000 507.640 ;
        RECT 4.000 500.840 496.000 506.240 ;
        RECT 4.400 499.440 496.000 500.840 ;
        RECT 4.000 494.040 496.000 499.440 ;
        RECT 4.400 492.640 496.000 494.040 ;
        RECT 4.000 487.240 496.000 492.640 ;
        RECT 4.400 485.840 496.000 487.240 ;
        RECT 4.000 479.760 496.000 485.840 ;
        RECT 4.400 478.360 496.000 479.760 ;
        RECT 4.000 472.960 496.000 478.360 ;
        RECT 4.400 471.560 496.000 472.960 ;
        RECT 4.000 466.160 496.000 471.560 ;
        RECT 4.400 464.760 496.000 466.160 ;
        RECT 4.000 458.680 496.000 464.760 ;
        RECT 4.400 457.280 496.000 458.680 ;
        RECT 4.000 451.880 496.000 457.280 ;
        RECT 4.400 450.480 496.000 451.880 ;
        RECT 4.000 445.080 496.000 450.480 ;
        RECT 4.400 443.680 496.000 445.080 ;
        RECT 4.000 437.600 496.000 443.680 ;
        RECT 4.400 436.200 496.000 437.600 ;
        RECT 4.000 430.800 496.000 436.200 ;
        RECT 4.400 429.400 496.000 430.800 ;
        RECT 4.000 424.000 496.000 429.400 ;
        RECT 4.400 422.600 496.000 424.000 ;
        RECT 4.000 417.200 496.000 422.600 ;
        RECT 4.400 415.800 496.000 417.200 ;
        RECT 4.000 409.720 496.000 415.800 ;
        RECT 4.400 408.320 496.000 409.720 ;
        RECT 4.000 402.920 496.000 408.320 ;
        RECT 4.400 401.520 496.000 402.920 ;
        RECT 4.000 396.120 496.000 401.520 ;
        RECT 4.400 394.720 496.000 396.120 ;
        RECT 4.000 388.640 496.000 394.720 ;
        RECT 4.400 387.240 496.000 388.640 ;
        RECT 4.000 381.840 496.000 387.240 ;
        RECT 4.400 380.440 496.000 381.840 ;
        RECT 4.000 375.040 496.000 380.440 ;
        RECT 4.400 373.640 496.000 375.040 ;
        RECT 4.000 368.240 496.000 373.640 ;
        RECT 4.400 366.840 496.000 368.240 ;
        RECT 4.000 360.760 496.000 366.840 ;
        RECT 4.400 359.360 496.000 360.760 ;
        RECT 4.000 353.960 496.000 359.360 ;
        RECT 4.400 352.560 496.000 353.960 ;
        RECT 4.000 347.160 496.000 352.560 ;
        RECT 4.400 345.760 496.000 347.160 ;
        RECT 4.000 339.680 496.000 345.760 ;
        RECT 4.400 338.280 496.000 339.680 ;
        RECT 4.000 332.880 496.000 338.280 ;
        RECT 4.400 331.480 496.000 332.880 ;
        RECT 4.000 326.080 496.000 331.480 ;
        RECT 4.400 324.680 496.000 326.080 ;
        RECT 4.000 319.280 496.000 324.680 ;
        RECT 4.400 317.880 496.000 319.280 ;
        RECT 4.000 311.800 496.000 317.880 ;
        RECT 4.400 310.400 496.000 311.800 ;
        RECT 4.000 305.000 496.000 310.400 ;
        RECT 4.400 303.600 496.000 305.000 ;
        RECT 4.000 298.200 496.000 303.600 ;
        RECT 4.400 296.800 496.000 298.200 ;
        RECT 4.000 290.720 496.000 296.800 ;
        RECT 4.400 289.320 496.000 290.720 ;
        RECT 4.000 283.920 496.000 289.320 ;
        RECT 4.400 282.520 496.000 283.920 ;
        RECT 4.000 277.120 496.000 282.520 ;
        RECT 4.400 275.720 496.000 277.120 ;
        RECT 4.000 270.320 496.000 275.720 ;
        RECT 4.400 268.920 496.000 270.320 ;
        RECT 4.000 262.840 496.000 268.920 ;
        RECT 4.400 261.440 496.000 262.840 ;
        RECT 4.000 256.040 496.000 261.440 ;
        RECT 4.400 254.640 496.000 256.040 ;
        RECT 4.000 249.240 496.000 254.640 ;
        RECT 4.400 247.840 496.000 249.240 ;
        RECT 4.000 241.760 496.000 247.840 ;
        RECT 4.400 240.360 496.000 241.760 ;
        RECT 4.000 234.960 496.000 240.360 ;
        RECT 4.400 233.560 496.000 234.960 ;
        RECT 4.000 228.160 496.000 233.560 ;
        RECT 4.400 226.760 496.000 228.160 ;
        RECT 4.000 220.680 496.000 226.760 ;
        RECT 4.400 219.280 496.000 220.680 ;
        RECT 4.000 213.880 496.000 219.280 ;
        RECT 4.400 212.480 496.000 213.880 ;
        RECT 4.000 207.080 496.000 212.480 ;
        RECT 4.400 205.680 496.000 207.080 ;
        RECT 4.000 200.280 496.000 205.680 ;
        RECT 4.400 198.880 496.000 200.280 ;
        RECT 4.000 192.800 496.000 198.880 ;
        RECT 4.400 191.400 496.000 192.800 ;
        RECT 4.000 186.000 496.000 191.400 ;
        RECT 4.400 184.600 496.000 186.000 ;
        RECT 4.000 179.200 496.000 184.600 ;
        RECT 4.400 177.800 496.000 179.200 ;
        RECT 4.000 175.800 496.000 177.800 ;
        RECT 4.000 174.400 495.600 175.800 ;
        RECT 4.000 171.720 496.000 174.400 ;
        RECT 4.400 170.320 496.000 171.720 ;
        RECT 4.000 164.920 496.000 170.320 ;
        RECT 4.400 163.520 496.000 164.920 ;
        RECT 4.000 158.120 496.000 163.520 ;
        RECT 4.400 156.720 496.000 158.120 ;
        RECT 4.000 151.320 496.000 156.720 ;
        RECT 4.400 149.920 496.000 151.320 ;
        RECT 4.000 143.840 496.000 149.920 ;
        RECT 4.400 142.440 496.000 143.840 ;
        RECT 4.000 137.040 496.000 142.440 ;
        RECT 4.400 135.640 496.000 137.040 ;
        RECT 4.000 130.240 496.000 135.640 ;
        RECT 4.400 128.840 496.000 130.240 ;
        RECT 4.000 122.760 496.000 128.840 ;
        RECT 4.400 121.360 496.000 122.760 ;
        RECT 4.000 115.960 496.000 121.360 ;
        RECT 4.400 114.560 496.000 115.960 ;
        RECT 4.000 109.160 496.000 114.560 ;
        RECT 4.400 107.760 496.000 109.160 ;
        RECT 4.000 102.360 496.000 107.760 ;
        RECT 4.400 100.960 496.000 102.360 ;
        RECT 4.000 94.880 496.000 100.960 ;
        RECT 4.400 93.480 496.000 94.880 ;
        RECT 4.000 88.080 496.000 93.480 ;
        RECT 4.400 86.680 496.000 88.080 ;
        RECT 4.000 81.280 496.000 86.680 ;
        RECT 4.400 79.880 496.000 81.280 ;
        RECT 4.000 73.800 496.000 79.880 ;
        RECT 4.400 72.400 496.000 73.800 ;
        RECT 4.000 67.000 496.000 72.400 ;
        RECT 4.400 65.600 496.000 67.000 ;
        RECT 4.000 60.200 496.000 65.600 ;
        RECT 4.400 58.800 496.000 60.200 ;
        RECT 4.000 53.400 496.000 58.800 ;
        RECT 4.400 52.000 496.000 53.400 ;
        RECT 4.000 45.920 496.000 52.000 ;
        RECT 4.400 44.520 496.000 45.920 ;
        RECT 4.000 39.120 496.000 44.520 ;
        RECT 4.400 37.720 496.000 39.120 ;
        RECT 4.000 32.320 496.000 37.720 ;
        RECT 4.400 30.920 496.000 32.320 ;
        RECT 4.000 24.840 496.000 30.920 ;
        RECT 4.400 23.440 496.000 24.840 ;
        RECT 4.000 18.040 496.000 23.440 ;
        RECT 4.400 16.640 496.000 18.040 ;
        RECT 4.000 11.240 496.000 16.640 ;
        RECT 4.400 9.840 496.000 11.240 ;
        RECT 4.000 4.440 496.000 9.840 ;
        RECT 4.400 3.575 496.000 4.440 ;
      LAYER met4 ;
        RECT 34.335 72.935 97.440 686.625 ;
        RECT 99.840 72.935 174.240 686.625 ;
        RECT 176.640 72.935 251.040 686.625 ;
        RECT 253.440 72.935 327.840 686.625 ;
        RECT 330.240 72.935 404.640 686.625 ;
        RECT 407.040 72.935 409.105 686.625 ;
  END
END Peripherals
END LIBRARY

