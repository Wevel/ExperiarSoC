* NGSPICE file created from ExperiarCore.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

.subckt ExperiarCore addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6]
+ addr0[7] addr0[8] addr1[0] addr1[1] addr1[2] addr1[3] addr1[4] addr1[5] addr1[6]
+ addr1[7] addr1[8] clk0 clk1 coreIndex[0] coreIndex[1] coreIndex[2] coreIndex[3]
+ coreIndex[4] coreIndex[5] coreIndex[6] coreIndex[7] core_wb_ack_i core_wb_adr_o[0]
+ core_wb_adr_o[10] core_wb_adr_o[11] core_wb_adr_o[12] core_wb_adr_o[13] core_wb_adr_o[14]
+ core_wb_adr_o[15] core_wb_adr_o[16] core_wb_adr_o[17] core_wb_adr_o[18] core_wb_adr_o[19]
+ core_wb_adr_o[1] core_wb_adr_o[20] core_wb_adr_o[21] core_wb_adr_o[22] core_wb_adr_o[23]
+ core_wb_adr_o[24] core_wb_adr_o[25] core_wb_adr_o[26] core_wb_adr_o[27] core_wb_adr_o[2]
+ core_wb_adr_o[3] core_wb_adr_o[4] core_wb_adr_o[5] core_wb_adr_o[6] core_wb_adr_o[7]
+ core_wb_adr_o[8] core_wb_adr_o[9] core_wb_cyc_o core_wb_data_i[0] core_wb_data_i[10]
+ core_wb_data_i[11] core_wb_data_i[12] core_wb_data_i[13] core_wb_data_i[14] core_wb_data_i[15]
+ core_wb_data_i[16] core_wb_data_i[17] core_wb_data_i[18] core_wb_data_i[19] core_wb_data_i[1]
+ core_wb_data_i[20] core_wb_data_i[21] core_wb_data_i[22] core_wb_data_i[23] core_wb_data_i[24]
+ core_wb_data_i[25] core_wb_data_i[26] core_wb_data_i[27] core_wb_data_i[28] core_wb_data_i[29]
+ core_wb_data_i[2] core_wb_data_i[30] core_wb_data_i[31] core_wb_data_i[3] core_wb_data_i[4]
+ core_wb_data_i[5] core_wb_data_i[6] core_wb_data_i[7] core_wb_data_i[8] core_wb_data_i[9]
+ core_wb_data_o[0] core_wb_data_o[10] core_wb_data_o[11] core_wb_data_o[12] core_wb_data_o[13]
+ core_wb_data_o[14] core_wb_data_o[15] core_wb_data_o[16] core_wb_data_o[17] core_wb_data_o[18]
+ core_wb_data_o[19] core_wb_data_o[1] core_wb_data_o[20] core_wb_data_o[21] core_wb_data_o[22]
+ core_wb_data_o[23] core_wb_data_o[24] core_wb_data_o[25] core_wb_data_o[26] core_wb_data_o[27]
+ core_wb_data_o[28] core_wb_data_o[29] core_wb_data_o[2] core_wb_data_o[30] core_wb_data_o[31]
+ core_wb_data_o[3] core_wb_data_o[4] core_wb_data_o[5] core_wb_data_o[6] core_wb_data_o[7]
+ core_wb_data_o[8] core_wb_data_o[9] core_wb_error_i core_wb_sel_o[0] core_wb_sel_o[1]
+ core_wb_sel_o[2] core_wb_sel_o[3] core_wb_stall_i core_wb_stb_o core_wb_we_o csb0[0]
+ csb0[1] csb1[0] csb1[1] din0[0] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15]
+ din0[16] din0[17] din0[18] din0[19] din0[1] din0[20] din0[21] din0[22] din0[23]
+ din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[2] din0[30] din0[31]
+ din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] dout0[0] dout0[10] dout0[11]
+ dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19]
+ dout0[1] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27]
+ dout0[28] dout0[29] dout0[2] dout0[30] dout0[31] dout0[32] dout0[33] dout0[34] dout0[35]
+ dout0[36] dout0[37] dout0[38] dout0[39] dout0[3] dout0[40] dout0[41] dout0[42] dout0[43]
+ dout0[44] dout0[45] dout0[46] dout0[47] dout0[48] dout0[49] dout0[4] dout0[50] dout0[51]
+ dout0[52] dout0[53] dout0[54] dout0[55] dout0[56] dout0[57] dout0[58] dout0[59]
+ dout0[5] dout0[60] dout0[61] dout0[62] dout0[63] dout0[6] dout0[7] dout0[8] dout0[9]
+ dout1[0] dout1[10] dout1[11] dout1[12] dout1[13] dout1[14] dout1[15] dout1[16] dout1[17]
+ dout1[18] dout1[19] dout1[1] dout1[20] dout1[21] dout1[22] dout1[23] dout1[24] dout1[25]
+ dout1[26] dout1[27] dout1[28] dout1[29] dout1[2] dout1[30] dout1[31] dout1[32] dout1[33]
+ dout1[34] dout1[35] dout1[36] dout1[37] dout1[38] dout1[39] dout1[3] dout1[40] dout1[41]
+ dout1[42] dout1[43] dout1[44] dout1[45] dout1[46] dout1[47] dout1[48] dout1[49]
+ dout1[4] dout1[50] dout1[51] dout1[52] dout1[53] dout1[54] dout1[55] dout1[56] dout1[57]
+ dout1[58] dout1[59] dout1[5] dout1[60] dout1[61] dout1[62] dout1[63] dout1[6] dout1[7]
+ dout1[8] dout1[9] irq[0] irq[10] irq[11] irq[12] irq[13] irq[14] irq[15] irq[1]
+ irq[2] irq[3] irq[4] irq[5] irq[6] irq[7] irq[8] irq[9] jtag_tck jtag_tdi jtag_tdo
+ jtag_tms localMemory_wb_ack_o localMemory_wb_adr_i[0] localMemory_wb_adr_i[10] localMemory_wb_adr_i[11]
+ localMemory_wb_adr_i[12] localMemory_wb_adr_i[13] localMemory_wb_adr_i[14] localMemory_wb_adr_i[15]
+ localMemory_wb_adr_i[16] localMemory_wb_adr_i[17] localMemory_wb_adr_i[18] localMemory_wb_adr_i[19]
+ localMemory_wb_adr_i[1] localMemory_wb_adr_i[20] localMemory_wb_adr_i[21] localMemory_wb_adr_i[22]
+ localMemory_wb_adr_i[23] localMemory_wb_adr_i[2] localMemory_wb_adr_i[3] localMemory_wb_adr_i[4]
+ localMemory_wb_adr_i[5] localMemory_wb_adr_i[6] localMemory_wb_adr_i[7] localMemory_wb_adr_i[8]
+ localMemory_wb_adr_i[9] localMemory_wb_cyc_i localMemory_wb_data_i[0] localMemory_wb_data_i[10]
+ localMemory_wb_data_i[11] localMemory_wb_data_i[12] localMemory_wb_data_i[13] localMemory_wb_data_i[14]
+ localMemory_wb_data_i[15] localMemory_wb_data_i[16] localMemory_wb_data_i[17] localMemory_wb_data_i[18]
+ localMemory_wb_data_i[19] localMemory_wb_data_i[1] localMemory_wb_data_i[20] localMemory_wb_data_i[21]
+ localMemory_wb_data_i[22] localMemory_wb_data_i[23] localMemory_wb_data_i[24] localMemory_wb_data_i[25]
+ localMemory_wb_data_i[26] localMemory_wb_data_i[27] localMemory_wb_data_i[28] localMemory_wb_data_i[29]
+ localMemory_wb_data_i[2] localMemory_wb_data_i[30] localMemory_wb_data_i[31] localMemory_wb_data_i[3]
+ localMemory_wb_data_i[4] localMemory_wb_data_i[5] localMemory_wb_data_i[6] localMemory_wb_data_i[7]
+ localMemory_wb_data_i[8] localMemory_wb_data_i[9] localMemory_wb_data_o[0] localMemory_wb_data_o[10]
+ localMemory_wb_data_o[11] localMemory_wb_data_o[12] localMemory_wb_data_o[13] localMemory_wb_data_o[14]
+ localMemory_wb_data_o[15] localMemory_wb_data_o[16] localMemory_wb_data_o[17] localMemory_wb_data_o[18]
+ localMemory_wb_data_o[19] localMemory_wb_data_o[1] localMemory_wb_data_o[20] localMemory_wb_data_o[21]
+ localMemory_wb_data_o[22] localMemory_wb_data_o[23] localMemory_wb_data_o[24] localMemory_wb_data_o[25]
+ localMemory_wb_data_o[26] localMemory_wb_data_o[27] localMemory_wb_data_o[28] localMemory_wb_data_o[29]
+ localMemory_wb_data_o[2] localMemory_wb_data_o[30] localMemory_wb_data_o[31] localMemory_wb_data_o[3]
+ localMemory_wb_data_o[4] localMemory_wb_data_o[5] localMemory_wb_data_o[6] localMemory_wb_data_o[7]
+ localMemory_wb_data_o[8] localMemory_wb_data_o[9] localMemory_wb_error_o localMemory_wb_sel_i[0]
+ localMemory_wb_sel_i[1] localMemory_wb_sel_i[2] localMemory_wb_sel_i[3] localMemory_wb_stall_o
+ localMemory_wb_stb_i localMemory_wb_we_i manufacturerID[0] manufacturerID[10] manufacturerID[1]
+ manufacturerID[2] manufacturerID[3] manufacturerID[4] manufacturerID[5] manufacturerID[6]
+ manufacturerID[7] manufacturerID[8] manufacturerID[9] partID[0] partID[10] partID[11]
+ partID[12] partID[13] partID[14] partID[15] partID[1] partID[2] partID[3] partID[4]
+ partID[5] partID[6] partID[7] partID[8] partID[9] probe_env[0] probe_env[1] probe_jtagInstruction[0]
+ probe_jtagInstruction[1] probe_jtagInstruction[2] probe_jtagInstruction[3] probe_jtagInstruction[4]
+ probe_programCounter[0] probe_programCounter[10] probe_programCounter[11] probe_programCounter[12]
+ probe_programCounter[13] probe_programCounter[14] probe_programCounter[15] probe_programCounter[16]
+ probe_programCounter[17] probe_programCounter[18] probe_programCounter[19] probe_programCounter[1]
+ probe_programCounter[20] probe_programCounter[21] probe_programCounter[22] probe_programCounter[23]
+ probe_programCounter[24] probe_programCounter[25] probe_programCounter[26] probe_programCounter[27]
+ probe_programCounter[28] probe_programCounter[29] probe_programCounter[2] probe_programCounter[30]
+ probe_programCounter[31] probe_programCounter[3] probe_programCounter[4] probe_programCounter[5]
+ probe_programCounter[6] probe_programCounter[7] probe_programCounter[8] probe_programCounter[9]
+ probe_state vccd1 versionID[0] versionID[1] versionID[2] versionID[3] vssd1 wb_clk_i
+ wb_rst_i web0 wmask0[0] wmask0[1] wmask0[2] wmask0[3]
XFILLER_228_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18869_ _27115_/Q _18748_/X _18867_/X _18868_/X vssd1 vssd1 vccd1 vccd1 _18869_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20900_ _23715_/A vssd1 vssd1 vccd1 vccd1 _20900_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_255_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21880_ _24455_/A vssd1 vssd1 vccd1 vccd1 _24473_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20831_ _20831_/A vssd1 vssd1 vccd1 vccd1 _25811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_254_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23550_ _26696_/Q _23549_/X _23556_/S vssd1 vssd1 vccd1 vccd1 _23551_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20762_ _20762_/A vssd1 vssd1 vccd1 vccd1 _25777_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_260 _20707_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_271 _18404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_282 _25815_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22501_ _22501_/A vssd1 vssd1 vccd1 vccd1 _26275_/D sky130_fd_sc_hd__clkbuf_1
X_23481_ _23481_/A vssd1 vssd1 vccd1 vccd1 _26671_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_293 _25823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20693_ _26287_/Q _20686_/X _20692_/Y _20684_/X vssd1 vssd1 vccd1 vccd1 _25750_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22432_ _22459_/A vssd1 vssd1 vccd1 vccd1 _22432_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25220_ _24988_/X _19624_/X _24771_/X _24725_/B _25219_/X vssd1 vssd1 vccd1 vccd1
+ _25220_/X sky130_fd_sc_hd__a221o_1
XFILLER_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22363_ _22388_/A _22362_/Y _22337_/A vssd1 vssd1 vccd1 vccd1 _22376_/S sky130_fd_sc_hd__o21a_2
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25151_ _25151_/A _25151_/B vssd1 vssd1 vccd1 vccd1 _25151_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24102_ _24102_/A vssd1 vssd1 vccd1 vccd1 _26918_/D sky130_fd_sc_hd__clkbuf_1
X_21314_ _20637_/A _21278_/X _21279_/X _21313_/X vssd1 vssd1 vccd1 vccd1 _21314_/X
+ sky130_fd_sc_hd__o211a_1
X_25082_ _25109_/A vssd1 vssd1 vccd1 vccd1 _25082_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22294_ _22310_/A vssd1 vssd1 vccd1 vccd1 _22294_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24033_ _26888_/Q _23549_/X _24037_/S vssd1 vssd1 vccd1 vccd1 _24034_/A sky130_fd_sc_hd__mux2_1
X_21245_ _21275_/A vssd1 vssd1 vccd1 vccd1 _21544_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21176_ _21188_/A _21176_/B vssd1 vssd1 vccd1 vccd1 _21177_/A sky130_fd_sc_hd__or2_1
XFILLER_278_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20127_ _20127_/A _20204_/B vssd1 vssd1 vccd1 vccd1 _20127_/X sky130_fd_sc_hd__xor2_1
XFILLER_131_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25984_ _25985_/CLK _25984_/D vssd1 vssd1 vccd1 vccd1 _25984_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_246_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24935_ _19930_/A _24927_/X _24934_/Y vssd1 vssd1 vccd1 vccd1 _27143_/D sky130_fd_sc_hd__o21a_1
X_20058_ _19881_/A _20056_/X _19771_/X _20664_/A vssd1 vssd1 vccd1 vccd1 _20084_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_58_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ _25482_/Q _12878_/B _12860_/B vssd1 vssd1 vccd1 vccd1 _13916_/C sky130_fd_sc_hd__o21ai_2
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24866_ _27123_/Q _24873_/B vssd1 vssd1 vccd1 vccd1 _24866_/Y sky130_fd_sc_hd__nand2_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26605_ _27330_/A _26605_/D vssd1 vssd1 vccd1 vccd1 _26605_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23817_ _23725_/X _26792_/Q _23821_/S vssd1 vssd1 vccd1 vccd1 _23818_/A sky130_fd_sc_hd__mux2_1
XFILLER_233_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24797_ _24794_/Y _24795_/X _24796_/X vssd1 vssd1 vccd1 vccd1 _27104_/D sky130_fd_sc_hd__a21oi_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _26064_/Q _25869_/Q _14551_/S vssd1 vssd1 vccd1 vccd1 _14550_/X sky130_fd_sc_hd__mux2_1
XFILLER_214_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26536_ _26673_/CLK _26536_/D vssd1 vssd1 vccd1 vccd1 _26536_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23748_ _23747_/X _26767_/Q _23748_/S vssd1 vssd1 vccd1 vccd1 _23749_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13472_/X _26886_/Q _26758_/Q _15496_/S _13494_/X vssd1 vssd1 vccd1 vccd1
+ _13501_/X sky130_fd_sc_hd__a221o_1
XFILLER_202_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26467_ _26467_/CLK _26467_/D vssd1 vssd1 vccd1 vccd1 _26467_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_198_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _25725_/Q _14481_/B vssd1 vssd1 vccd1 vccd1 _14481_/X sky130_fd_sc_hd__or2_1
XFILLER_202_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23679_ _23679_/A vssd1 vssd1 vccd1 vccd1 _26745_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16220_ _16218_/X _16219_/X _16224_/S vssd1 vssd1 vccd1 vccd1 _16220_/X sky130_fd_sc_hd__mux2_1
X_25418_ _23718_/X _27305_/Q _25426_/S vssd1 vssd1 vccd1 vccd1 _25419_/A sky130_fd_sc_hd__mux2_1
X_13432_ _12770_/A _26598_/Q _15471_/S _26338_/Q _13431_/X vssd1 vssd1 vccd1 vccd1
+ _13432_/X sky130_fd_sc_hd__o221a_1
X_26398_ _26462_/CLK _26398_/D vssd1 vssd1 vccd1 vccd1 _26398_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16151_ _26641_/Q _26737_/Q _16151_/S vssd1 vssd1 vccd1 vccd1 _16151_/X sky130_fd_sc_hd__mux2_1
X_25349_ _25349_/A vssd1 vssd1 vccd1 vccd1 _27274_/D sky130_fd_sc_hd__clkbuf_1
X_13363_ _13363_/A vssd1 vssd1 vccd1 vccd1 _15317_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_167_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15102_ _14793_/A _15095_/X _15101_/X _14808_/A vssd1 vssd1 vccd1 vccd1 _15102_/X
+ sky130_fd_sc_hd__o211a_1
X_16082_ _16065_/X _16081_/X _14591_/A vssd1 vssd1 vccd1 vccd1 _16082_/X sky130_fd_sc_hd__a21o_2
X_13294_ _15331_/A vssd1 vssd1 vccd1 vccd1 _15321_/A sky130_fd_sc_hd__buf_4
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27019_ _27022_/CLK _27019_/D vssd1 vssd1 vccd1 vccd1 _27019_/Q sky130_fd_sc_hd__dfxtp_1
X_19910_ _19910_/A vssd1 vssd1 vccd1 vccd1 _20194_/B sky130_fd_sc_hd__clkbuf_2
X_15033_ _15029_/X _15030_/X _16241_/S vssd1 vssd1 vccd1 vccd1 _15033_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19841_ _19841_/A _19841_/B vssd1 vssd1 vccd1 vccd1 _19841_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_150_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19772_ _19772_/A vssd1 vssd1 vccd1 vccd1 _20637_/A sky130_fd_sc_hd__buf_6
X_16984_ _16883_/X _16954_/A _16956_/A _16882_/X _16983_/X vssd1 vssd1 vccd1 vccd1
+ _16984_/X sky130_fd_sc_hd__a221o_1
XFILLER_283_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15935_ _13472_/X _26889_/Q _26761_/Q _15197_/A _13359_/A vssd1 vssd1 vccd1 vccd1
+ _15935_/X sky130_fd_sc_hd__a221o_1
X_18723_ _19087_/A vssd1 vssd1 vccd1 vccd1 _18723_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_60_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26468_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18654_ _27079_/Q _18508_/X _18509_/X _27177_/Q _18510_/X vssd1 vssd1 vccd1 vccd1
+ _18654_/X sky130_fd_sc_hd__a221o_1
XFILLER_236_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ _13638_/X _15849_/Y _15865_/Y _14827_/A vssd1 vssd1 vccd1 vccd1 _15866_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_252_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17605_ _25920_/Q _17554_/A _13389_/Y _17577_/X vssd1 vssd1 vccd1 vccd1 _17605_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14817_ _14817_/A vssd1 vssd1 vccd1 vccd1 _14818_/A sky130_fd_sc_hd__buf_4
XFILLER_236_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18585_ _13798_/X _18285_/X _18584_/X _18409_/X _25606_/Q vssd1 vssd1 vccd1 vccd1
+ _18586_/B sky130_fd_sc_hd__a32o_1
XFILLER_251_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15797_ _26922_/Q _15797_/B vssd1 vssd1 vccd1 vccd1 _15797_/X sky130_fd_sc_hd__or2_1
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17536_ _17554_/A vssd1 vssd1 vccd1 vccd1 _17536_/X sky130_fd_sc_hd__buf_2
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14748_ _14891_/A vssd1 vssd1 vccd1 vccd1 _14991_/S sky130_fd_sc_hd__buf_4
XFILLER_225_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17467_ _26250_/Q _17454_/A _17460_/A _25978_/Q vssd1 vssd1 vccd1 vccd1 _17694_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_178_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14679_ _14679_/A vssd1 vssd1 vccd1 vccd1 _14679_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19206_ _25524_/Q _18559_/X _19203_/X _19205_/X _18574_/X vssd1 vssd1 vccd1 vccd1
+ _19206_/X sky130_fd_sc_hd__o221a_1
X_16418_ _27290_/Q _26483_/Q _16422_/S vssd1 vssd1 vccd1 vccd1 _16418_/X sky130_fd_sc_hd__mux2_1
X_17398_ _17395_/X _17399_/C _25551_/Q vssd1 vssd1 vccd1 vccd1 _17400_/B sky130_fd_sc_hd__a21oi_1
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19137_ _25554_/Q _18568_/X _19136_/X _19069_/X _18572_/X vssd1 vssd1 vccd1 vccd1
+ _19137_/X sky130_fd_sc_hd__a221o_1
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16349_ _16339_/X _16342_/X _16345_/X _16348_/X _14758_/A _14778_/A vssd1 vssd1 vccd1
+ vccd1 _16350_/B sky130_fd_sc_hd__mux4_1
XFILLER_146_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19068_ _26960_/Q _18569_/X _18570_/X _26992_/Q vssd1 vssd1 vccd1 vccd1 _19068_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput401 _17009_/X vssd1 vssd1 vccd1 vccd1 din0[3] sky130_fd_sc_hd__buf_2
Xoutput412 _25947_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[11] sky130_fd_sc_hd__buf_2
XFILLER_161_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18019_ _20141_/B vssd1 vssd1 vccd1 vccd1 _18019_/X sky130_fd_sc_hd__buf_2
Xoutput423 _25957_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[21] sky130_fd_sc_hd__buf_2
Xoutput434 _25967_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[31] sky130_fd_sc_hd__buf_2
Xoutput445 _26232_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[0] sky130_fd_sc_hd__buf_2
XFILLER_99_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21030_ _21030_/A vssd1 vssd1 vccd1 vccd1 _25884_/D sky130_fd_sc_hd__clkbuf_1
Xoutput456 _25739_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[15] sky130_fd_sc_hd__buf_2
Xoutput467 _25749_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[25] sky130_fd_sc_hd__buf_2
XFILLER_99_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput478 _25730_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[6] sky130_fd_sc_hd__buf_2
XFILLER_102_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22981_ _22981_/A vssd1 vssd1 vccd1 vccd1 _26463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_274_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24720_ _24720_/A vssd1 vssd1 vccd1 vccd1 _24720_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_256_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21932_ _21932_/A vssd1 vssd1 vccd1 vccd1 _26082_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24651_ _27071_/Q _24636_/X _24650_/X vssd1 vssd1 vccd1 vccd1 _27071_/D sky130_fd_sc_hd__o21ba_1
XFILLER_282_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21863_ _21863_/A vssd1 vssd1 vccd1 vccd1 _26059_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23602_ _23602_/A vssd1 vssd1 vccd1 vccd1 _26712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_271_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20814_ _25803_/Q vssd1 vssd1 vccd1 vccd1 _20815_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_179_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24582_ _24582_/A _24582_/B vssd1 vssd1 vccd1 vccd1 _24582_/Y sky130_fd_sc_hd__nand2_1
X_21794_ _22962_/A _23788_/A vssd1 vssd1 vccd1 vccd1 _21851_/A sky130_fd_sc_hd__nor2_8
XFILLER_196_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26321_ _26326_/CLK _26321_/D vssd1 vssd1 vccd1 vccd1 _26321_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_169_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23533_ _23533_/A vssd1 vssd1 vccd1 vccd1 _23533_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20745_ _20745_/A vssd1 vssd1 vccd1 vccd1 _25769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26252_ _26307_/CLK _26252_/D vssd1 vssd1 vccd1 vccd1 _26252_/Q sky130_fd_sc_hd__dfxtp_1
X_23464_ _23464_/A vssd1 vssd1 vccd1 vccd1 _26663_/D sky130_fd_sc_hd__clkbuf_1
X_20676_ _26280_/Q _20673_/X _20675_/X _20671_/X vssd1 vssd1 vccd1 vccd1 _25743_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25203_ _24703_/B _25198_/X _25196_/X _27213_/Q _25199_/X vssd1 vssd1 vccd1 vccd1
+ _27213_/D sky130_fd_sc_hd__o221a_1
X_22415_ _22415_/A vssd1 vssd1 vccd1 vccd1 _22554_/A sky130_fd_sc_hd__clkbuf_2
X_26183_ _26319_/CLK _26183_/D vssd1 vssd1 vccd1 vccd1 _26183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23395_ _26633_/Q _23079_/X _23397_/S vssd1 vssd1 vccd1 vccd1 _23396_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25134_ _19246_/A _25113_/X _25133_/X vssd1 vssd1 vccd1 vccd1 _25134_/Y sky130_fd_sc_hd__o21ai_1
X_22346_ _26235_/Q _26227_/Q _22350_/S vssd1 vssd1 vccd1 vccd1 _22346_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22277_ _26204_/Q _22264_/X _22270_/X _26305_/Q _22271_/X vssd1 vssd1 vccd1 vccd1
+ _22277_/X sky130_fd_sc_hd__a221o_1
XFILLER_163_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25065_ _25065_/A vssd1 vssd1 vccd1 vccd1 _25065_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_275_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24016_ _24016_/A vssd1 vssd1 vccd1 vccd1 _26880_/D sky130_fd_sc_hd__clkbuf_1
X_21228_ _21244_/A _22536_/B _21227_/X vssd1 vssd1 vccd1 vccd1 _21228_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_151_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21159_ _21159_/A vssd1 vssd1 vccd1 vccd1 _25924_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25967_ _27049_/CLK _25967_/D vssd1 vssd1 vccd1 vccd1 _25967_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_58_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13981_ _13180_/A _19800_/A _13980_/X vssd1 vssd1 vccd1 vccd1 _14022_/A sky130_fd_sc_hd__o21a_2
XFILLER_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15720_ _15716_/X _15719_/X _15720_/S vssd1 vssd1 vccd1 vccd1 _15720_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12932_ _13397_/B vssd1 vssd1 vccd1 vccd1 _14025_/B sky130_fd_sc_hd__clkbuf_1
X_24918_ _24559_/A _24917_/X _24909_/X vssd1 vssd1 vccd1 vccd1 _24918_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_86_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25898_ _27292_/CLK _25898_/D vssd1 vssd1 vccd1 vccd1 _25898_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_74_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _15645_/S _15650_/X _13703_/A vssd1 vssd1 vccd1 vccd1 _15651_/X sky130_fd_sc_hd__a21o_1
XFILLER_233_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12863_ _13569_/A _15704_/A _12873_/A vssd1 vssd1 vccd1 vccd1 _12863_/X sky130_fd_sc_hd__a21o_1
XFILLER_160_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24849_ _24874_/A vssd1 vssd1 vccd1 vccd1 _24849_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14602_ _14602_/A vssd1 vssd1 vccd1 vccd1 _14603_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18370_ _18734_/A vssd1 vssd1 vccd1 vccd1 _18371_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15582_/A vssd1 vssd1 vccd1 vccd1 _16176_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_15_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _25578_/Q _17162_/A vssd1 vssd1 vccd1 vccd1 _18194_/B sky130_fd_sc_hd__nor2_2
XFILLER_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _17317_/X _17322_/C _25527_/Q vssd1 vssd1 vccd1 vccd1 _17323_/B sky130_fd_sc_hd__a21oi_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _14453_/X _26684_/Q _26812_/Q _16021_/S _13943_/A vssd1 vssd1 vccd1 vccd1
+ _14533_/X sky130_fd_sc_hd__a221o_1
XFILLER_42_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26519_ _26939_/CLK _26519_/D vssd1 vssd1 vccd1 vccd1 _26519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17252_ _17252_/A _17252_/B vssd1 vssd1 vccd1 vccd1 _25505_/D sky130_fd_sc_hd__nor2_1
X_14464_ _26781_/Q _26425_/Q _14539_/S vssd1 vssd1 vccd1 vccd1 _14464_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16203_ _19141_/A vssd1 vssd1 vccd1 vccd1 _20227_/A sky130_fd_sc_hd__inv_2
X_13415_ _14713_/B _13406_/X _13414_/X _15538_/A vssd1 vssd1 vccd1 vccd1 _13415_/X
+ sky130_fd_sc_hd__a211o_1
X_17183_ _25488_/Q _17185_/B vssd1 vssd1 vccd1 vccd1 _17183_/X sky130_fd_sc_hd__or2_1
X_14395_ _14077_/A _14387_/X _14394_/X _13508_/A vssd1 vssd1 vccd1 vccd1 _14395_/X
+ sky130_fd_sc_hd__a31o_1
X_16134_ _27316_/Q _26573_/Q _16134_/S vssd1 vssd1 vccd1 vccd1 _16134_/X sky130_fd_sc_hd__mux2_1
X_13346_ _13346_/A vssd1 vssd1 vccd1 vccd1 _13347_/A sky130_fd_sc_hd__buf_8
XFILLER_183_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16065_ _14621_/A _16052_/X _16056_/X _16064_/X _14681_/A vssd1 vssd1 vccd1 vccd1
+ _16065_/X sky130_fd_sc_hd__a311o_1
X_13277_ _13277_/A vssd1 vssd1 vccd1 vccd1 _13278_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15016_ _16396_/S vssd1 vssd1 vccd1 vccd1 _16385_/S sky130_fd_sc_hd__buf_2
XFILLER_190_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19824_ _19824_/A _19824_/B vssd1 vssd1 vccd1 vccd1 _19824_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19755_ _20186_/A vssd1 vssd1 vccd1 vccd1 _19755_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16967_ _14977_/X _16952_/X _16887_/X vssd1 vssd1 vccd1 vccd1 _16970_/B sky130_fd_sc_hd__o21ai_2
XFILLER_111_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18706_ _18474_/A _18703_/Y _18705_/X vssd1 vssd1 vccd1 vccd1 _18706_/X sky130_fd_sc_hd__o21ba_1
X_15918_ _13254_/A _25842_/Q _26042_/Q _15496_/S _15932_/A vssd1 vssd1 vccd1 vccd1
+ _15918_/X sky130_fd_sc_hd__a221o_1
XFILLER_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16898_ _16887_/X _16896_/X _16897_/X vssd1 vssd1 vccd1 vccd1 _16899_/B sky130_fd_sc_hd__a21boi_4
X_19686_ _19686_/A _19686_/B vssd1 vssd1 vccd1 vccd1 _19687_/B sky130_fd_sc_hd__and2_1
XFILLER_64_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15849_ _15837_/X _15840_/X _15848_/X vssd1 vssd1 vccd1 vccd1 _15849_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_37_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18637_ _19046_/B _19574_/A _18636_/X vssd1 vssd1 vccd1 vccd1 _18637_/X sky130_fd_sc_hd__o21a_1
XFILLER_280_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18568_ _18568_/A vssd1 vssd1 vccd1 vccd1 _18568_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17519_ _25902_/Q _17517_/X _14489_/Y _17518_/X vssd1 vssd1 vccd1 vccd1 _17519_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_177_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18499_ _18366_/X _18498_/X _13909_/B vssd1 vssd1 vccd1 vccd1 _18499_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20530_ _20529_/X _25701_/Q _20530_/S vssd1 vssd1 vccd1 vccd1 _20531_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20461_ _27163_/Q _20460_/Y _20461_/S vssd1 vssd1 vccd1 vccd1 _20461_/X sky130_fd_sc_hd__mux2_2
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22200_ _22200_/A vssd1 vssd1 vccd1 vccd1 _22200_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_23180_ _23180_/A vssd1 vssd1 vccd1 vccd1 _26537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20392_ _27160_/Q _20391_/Y _20461_/S vssd1 vssd1 vccd1 vccd1 _20392_/X sky130_fd_sc_hd__mux2_2
XFILLER_106_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22131_ _24441_/A vssd1 vssd1 vccd1 vccd1 _22195_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_173_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22062_ _26140_/Q _20910_/X _22066_/S vssd1 vssd1 vccd1 vccd1 _22063_/A sky130_fd_sc_hd__mux2_1
X_21013_ _25877_/Q _20897_/X _21015_/S vssd1 vssd1 vccd1 vccd1 _21014_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput286 _17064_/X vssd1 vssd1 vccd1 vccd1 addr0[1] sky130_fd_sc_hd__buf_2
Xoutput297 _16994_/X vssd1 vssd1 vccd1 vccd1 addr1[3] sky130_fd_sc_hd__buf_2
XFILLER_114_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26870_ _27257_/CLK _26870_/D vssd1 vssd1 vccd1 vccd1 _26870_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_4 _22368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_25821_ _27314_/CLK _25821_/D vssd1 vssd1 vccd1 vccd1 _25821_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25752_ _26292_/CLK _25752_/D vssd1 vssd1 vccd1 vccd1 _25752_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22964_ _23032_/S vssd1 vssd1 vccd1 vccd1 _22973_/S sky130_fd_sc_hd__buf_2
XFILLER_229_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24703_ _24703_/A _24703_/B vssd1 vssd1 vccd1 vccd1 _24703_/Y sky130_fd_sc_hd__nand2_2
X_21915_ _21915_/A vssd1 vssd1 vccd1 vccd1 _26074_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25683_ _26286_/CLK _25683_/D vssd1 vssd1 vccd1 vccd1 _25683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22895_ _26425_/Q _22647_/X _22901_/S vssd1 vssd1 vccd1 vccd1 _22896_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24634_ _24749_/A _24740_/A vssd1 vssd1 vccd1 vccd1 _24635_/A sky130_fd_sc_hd__nand2_1
X_21846_ _21846_/A vssd1 vssd1 vccd1 vccd1 _26051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24565_ _24923_/A _24569_/B vssd1 vssd1 vccd1 vccd1 _24565_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21777_ _21777_/A vssd1 vssd1 vccd1 vccd1 _26021_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26304_ _26327_/CLK _26304_/D vssd1 vssd1 vccd1 vccd1 _26304_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_169_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23516_ _23516_/A vssd1 vssd1 vccd1 vccd1 _26685_/D sky130_fd_sc_hd__clkbuf_1
X_20728_ _20508_/X _25762_/Q _20728_/S vssd1 vssd1 vccd1 vccd1 _20729_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27284_ _27284_/CLK _27284_/D vssd1 vssd1 vccd1 vccd1 _27284_/Q sky130_fd_sc_hd__dfxtp_1
X_24496_ _24472_/X _25621_/Q _24495_/X vssd1 vssd1 vccd1 vccd1 _24739_/B sky130_fd_sc_hd__o21a_4
XFILLER_11_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26235_ _26520_/CLK _26235_/D vssd1 vssd1 vccd1 vccd1 _26235_/Q sky130_fd_sc_hd__dfxtp_4
X_23447_ _26656_/Q _23050_/X _23447_/S vssd1 vssd1 vccd1 vccd1 _23448_/A sky130_fd_sc_hd__mux2_1
X_20659_ _26274_/Q _20646_/X _20656_/X _20658_/X vssd1 vssd1 vccd1 vccd1 _25737_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ _20868_/B vssd1 vssd1 vccd1 vccd1 _21793_/A sky130_fd_sc_hd__inv_2
X_26166_ _27264_/CLK _26166_/D vssd1 vssd1 vccd1 vccd1 _26166_/Q sky130_fd_sc_hd__dfxtp_1
X_14180_ _12767_/A _26592_/Q _14169_/B _26332_/Q _13062_/A vssd1 vssd1 vccd1 vccd1
+ _14180_/X sky130_fd_sc_hd__o221a_1
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23378_ _26625_/Q _23053_/X _23386_/S vssd1 vssd1 vccd1 vccd1 _23379_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _14352_/S vssd1 vssd1 vccd1 vccd1 _14515_/S sky130_fd_sc_hd__buf_2
X_25117_ _24729_/Y _25097_/X _25116_/Y _25109_/X vssd1 vssd1 vccd1 vccd1 _25117_/X
+ sky130_fd_sc_hd__a31o_1
X_22329_ _26222_/Q _22154_/A _22270_/A _26323_/Q _22271_/A vssd1 vssd1 vccd1 vccd1
+ _22329_/X sky130_fd_sc_hd__a221o_1
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26097_ _26240_/CLK _26097_/D vssd1 vssd1 vccd1 vccd1 _26097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13062_ _13062_/A vssd1 vssd1 vccd1 vccd1 _14264_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_155_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25048_ _25668_/Q _25038_/X _25033_/X _18541_/A _25024_/X vssd1 vssd1 vccd1 vccd1
+ _25048_/X sky130_fd_sc_hd__a221o_1
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17870_ _14570_/B _17780_/B _17909_/S vssd1 vssd1 vccd1 vccd1 _17870_/X sky130_fd_sc_hd__mux2_1
XFILLER_215_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16821_ _16828_/A _16824_/B _16862_/B vssd1 vssd1 vccd1 vccd1 _16822_/A sky130_fd_sc_hd__and3_4
XFILLER_238_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26999_ _27000_/CLK _26999_/D vssd1 vssd1 vccd1 vccd1 _26999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19540_ _25650_/Q _19549_/B vssd1 vssd1 vccd1 vccd1 _19540_/X sky130_fd_sc_hd__or2_1
X_16752_ _22505_/A _16742_/X _16743_/X _18968_/B vssd1 vssd1 vccd1 vccd1 _16752_/X
+ sky130_fd_sc_hd__a22o_1
X_13964_ _13239_/A _13962_/X _13963_/X _13278_/A vssd1 vssd1 vccd1 vccd1 _13964_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_93_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15703_ _18938_/S _15703_/B vssd1 vssd1 vccd1 vccd1 _16625_/A sky130_fd_sc_hd__nand2_2
XFILLER_46_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12915_ _12915_/A vssd1 vssd1 vccd1 vccd1 _13922_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_74_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19471_ _18742_/X _19461_/X _19470_/X vssd1 vssd1 vccd1 vccd1 _19471_/X sky130_fd_sc_hd__a21o_4
X_16683_ _16678_/Y _16679_/X _16681_/Y vssd1 vssd1 vccd1 vccd1 _16683_/X sky130_fd_sc_hd__a21bo_1
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13895_ _15982_/S _13894_/X _14089_/S vssd1 vssd1 vccd1 vccd1 _13895_/X sky130_fd_sc_hd__a21o_1
XFILLER_46_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15634_ _27279_/Q _26472_/Q _15634_/S vssd1 vssd1 vccd1 vccd1 _15634_/X sky130_fd_sc_hd__mux2_1
X_18422_ _16717_/A _18328_/A _17803_/B vssd1 vssd1 vccd1 vccd1 _18423_/B sky130_fd_sc_hd__a21o_1
X_12846_ _14403_/A _12846_/B vssd1 vssd1 vccd1 vccd1 _12846_/X sky130_fd_sc_hd__or2_1
XFILLER_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _18942_/B vssd1 vssd1 vccd1 vccd1 _19046_/B sky130_fd_sc_hd__buf_2
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15565_ _26537_/Q _26145_/Q _15566_/S vssd1 vssd1 vccd1 vccd1 _15565_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _12777_/A vssd1 vssd1 vccd1 vccd1 _17712_/B sky130_fd_sc_hd__buf_6
XFILLER_199_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _17332_/A _17304_/B _17305_/B vssd1 vssd1 vccd1 vccd1 _25521_/D sky130_fd_sc_hd__nor3_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _13029_/A _14512_/Y _14515_/X _13124_/A vssd1 vssd1 vccd1 vccd1 _14516_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18284_ _18284_/A vssd1 vssd1 vccd1 vccd1 _25601_/D sky130_fd_sc_hd__clkbuf_1
X_15496_ _26082_/Q _25887_/Q _15496_/S vssd1 vssd1 vccd1 vccd1 _15496_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17235_ _17414_/A vssd1 vssd1 vccd1 vccd1 _17235_/X sky130_fd_sc_hd__buf_12
XFILLER_202_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14447_ _14447_/A _14447_/B vssd1 vssd1 vccd1 vccd1 _23514_/A sky130_fd_sc_hd__and2_4
XFILLER_266_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17166_ _17992_/B vssd1 vssd1 vccd1 vccd1 _18077_/A sky130_fd_sc_hd__clkbuf_2
X_14378_ _13540_/A _14374_/X _14377_/X _13210_/A vssd1 vssd1 vccd1 vccd1 _14378_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16117_ _16117_/A _16117_/B vssd1 vssd1 vccd1 vccd1 _16117_/Y sky130_fd_sc_hd__nor2_1
X_13329_ _15769_/A vssd1 vssd1 vccd1 vccd1 _13330_/A sky130_fd_sc_hd__clkbuf_4
X_17097_ _22387_/B _22406_/B vssd1 vssd1 vccd1 vccd1 _22230_/C sky130_fd_sc_hd__nor2_1
XFILLER_143_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16048_ _25617_/Q _14596_/A _16047_/X _14617_/A vssd1 vssd1 vccd1 vccd1 _23571_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_9_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19807_ _19808_/A _19808_/B vssd1 vssd1 vccd1 vccd1 _19809_/A sky130_fd_sc_hd__or2_1
XFILLER_69_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17999_ _16801_/A _16788_/A _18366_/A _16800_/B _17998_/Y vssd1 vssd1 vccd1 vccd1
+ _17999_/X sky130_fd_sc_hd__o221a_1
XFILLER_284_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19738_ _19926_/A vssd1 vssd1 vccd1 vccd1 _19738_/X sky130_fd_sc_hd__buf_2
XFILLER_244_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19669_ _19661_/X _19666_/X _19708_/A _19709_/A vssd1 vssd1 vccd1 vccd1 _19673_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_241_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21700_ _21700_/A vssd1 vssd1 vccd1 vccd1 _25988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22680_ _26339_/Q _22679_/X _22689_/S vssd1 vssd1 vccd1 vccd1 _22681_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21631_ _21586_/X _19441_/X _21587_/X _25827_/Q _21346_/X vssd1 vssd1 vccd1 vccd1
+ _21631_/X sky130_fd_sc_hd__a221o_1
XFILLER_178_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24350_ _25490_/Q _21208_/D _24350_/S vssd1 vssd1 vccd1 vccd1 _24989_/A sky130_fd_sc_hd__mux2_1
X_21562_ _26587_/Q _21562_/B _21562_/C _21562_/D vssd1 vssd1 vccd1 vccd1 _21563_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_20_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23301_ _23301_/A vssd1 vssd1 vccd1 vccd1 _26591_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20513_ _20622_/S vssd1 vssd1 vccd1 vccd1 _20530_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_220_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24281_ _26984_/Q _24284_/C _24271_/X vssd1 vssd1 vccd1 vccd1 _24281_/Y sky130_fd_sc_hd__a21oi_1
X_21493_ _21487_/Y _21491_/X _21492_/X vssd1 vssd1 vccd1 vccd1 _21493_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_176_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26020_ _27329_/A _26020_/D vssd1 vssd1 vccd1 vccd1 _26020_/Q sky130_fd_sc_hd__dfxtp_1
X_23232_ _23232_/A vssd1 vssd1 vccd1 vccd1 _26560_/D sky130_fd_sc_hd__clkbuf_1
X_20444_ _20405_/B _20426_/B _20470_/A vssd1 vssd1 vccd1 vccd1 _20450_/B sky130_fd_sc_hd__o21ai_1
XFILLER_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23163_ _23209_/S vssd1 vssd1 vccd1 vccd1 _23172_/S sky130_fd_sc_hd__buf_6
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20375_ _25751_/Q vssd1 vssd1 vccd1 vccd1 _20694_/A sky130_fd_sc_hd__buf_6
XFILLER_279_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22114_ _22121_/A _22170_/A vssd1 vssd1 vccd1 vccd1 _22206_/A sky130_fd_sc_hd__nor2_1
X_23094_ _23094_/A vssd1 vssd1 vccd1 vccd1 _26505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22045_ _22045_/A vssd1 vssd1 vccd1 vccd1 _26132_/D sky130_fd_sc_hd__clkbuf_1
X_26922_ _27278_/CLK _26922_/D vssd1 vssd1 vccd1 vccd1 _26922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26853_ _26916_/CLK _26853_/D vssd1 vssd1 vccd1 vccd1 _26853_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_134_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25804_ _27295_/CLK _25804_/D vssd1 vssd1 vccd1 vccd1 _25804_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_188_wb_clk_i _26681_/CLK vssd1 vssd1 vccd1 vccd1 _27292_/CLK sky130_fd_sc_hd__clkbuf_16
X_26784_ _27299_/CLK _26784_/D vssd1 vssd1 vccd1 vccd1 _26784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23996_ _26872_/Q _23600_/X _23998_/S vssd1 vssd1 vccd1 vccd1 _23997_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_117_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26995_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_25735_ _26271_/CLK _25735_/D vssd1 vssd1 vccd1 vccd1 _25735_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22947_ _22947_/A vssd1 vssd1 vccd1 vccd1 _22956_/S sky130_fd_sc_hd__buf_6
XFILLER_16_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12700_ _12700_/A vssd1 vssd1 vccd1 vccd1 _14362_/A sky130_fd_sc_hd__buf_12
XFILLER_245_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13680_ _13791_/A _13675_/X _13679_/X _13479_/A vssd1 vssd1 vccd1 vccd1 _13680_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25666_ _27132_/CLK _25666_/D vssd1 vssd1 vccd1 vccd1 _25666_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_70_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22878_ _26418_/Q _22727_/X _22884_/S vssd1 vssd1 vccd1 vccd1 _22879_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24617_ _27062_/Q _24615_/X _24616_/Y _24606_/X vssd1 vssd1 vccd1 vccd1 _27062_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21829_ _21851_/A vssd1 vssd1 vccd1 vccd1 _21838_/S sky130_fd_sc_hd__buf_4
XPHY_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25597_ _25599_/CLK _25597_/D vssd1 vssd1 vccd1 vccd1 _25597_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15350_ _27315_/Q _26572_/Q _16395_/S vssd1 vssd1 vccd1 vccd1 _15350_/X sky130_fd_sc_hd__mux2_1
XPHY_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24548_ _24548_/A _24553_/B vssd1 vssd1 vccd1 vccd1 _24548_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14301_ _26911_/Q _26395_/Q _14308_/S vssd1 vssd1 vccd1 vccd1 _14301_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27267_ _27267_/CLK _27267_/D vssd1 vssd1 vccd1 vccd1 _27267_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_196_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15281_ _15279_/X _15280_/X _16324_/S vssd1 vssd1 vccd1 vccd1 _15281_/X sky130_fd_sc_hd__mux2_1
X_24479_ _27024_/Q _24448_/X _24478_/Y _24470_/X vssd1 vssd1 vccd1 vccd1 _27024_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_200_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17020_ _17020_/A vssd1 vssd1 vccd1 vccd1 _17063_/A sky130_fd_sc_hd__clkbuf_2
X_26218_ _26319_/CLK _26218_/D vssd1 vssd1 vccd1 vccd1 _26218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14232_ _25728_/Q _16031_/S vssd1 vssd1 vccd1 vccd1 _14232_/X sky130_fd_sc_hd__or2_2
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27198_ _27198_/CLK _27198_/D vssd1 vssd1 vccd1 vccd1 _27198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14163_ _14153_/X _26688_/Q _26816_/Q _14009_/S _13611_/A vssd1 vssd1 vccd1 vccd1
+ _14163_/X sky130_fd_sc_hd__a221o_1
XFILLER_171_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26149_ _27284_/CLK _26149_/D vssd1 vssd1 vccd1 vccd1 _26149_/Q sky130_fd_sc_hd__dfxtp_1
X_13114_ _13114_/A vssd1 vssd1 vccd1 vccd1 _14621_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_152_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14094_ _14268_/S vssd1 vssd1 vccd1 vccd1 _14165_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18971_ _19287_/B vssd1 vssd1 vccd1 vccd1 _18971_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13045_ _26631_/Q _26727_/Q _15566_/S vssd1 vssd1 vccd1 vccd1 _13045_/X sky130_fd_sc_hd__mux2_1
X_17922_ _14562_/B _17852_/B _18681_/A vssd1 vssd1 vccd1 vccd1 _17922_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17853_ _19389_/B _17849_/Y _19389_/C _17852_/Y _16462_/A vssd1 vssd1 vccd1 vccd1
+ _17853_/X sky130_fd_sc_hd__a311o_1
XFILLER_94_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16804_ _16952_/A _16842_/A _16697_/D _16803_/X vssd1 vssd1 vccd1 vccd1 _16804_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17784_ _17784_/A _17784_/B vssd1 vssd1 vccd1 vccd1 _17784_/Y sky130_fd_sc_hd__nand2_1
X_14996_ _26936_/Q _26420_/Q _14996_/S vssd1 vssd1 vccd1 vccd1 _14996_/X sky130_fd_sc_hd__mux2_1
XFILLER_219_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19523_ _25644_/Q _19523_/B vssd1 vssd1 vccd1 vccd1 _19523_/X sky130_fd_sc_hd__or2_1
X_13947_ _14535_/A _13947_/B _13947_/C vssd1 vssd1 vccd1 vccd1 _13947_/X sky130_fd_sc_hd__or3_1
XFILLER_35_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16735_ _16735_/A _16735_/B vssd1 vssd1 vccd1 vccd1 _16735_/X sky130_fd_sc_hd__xor2_4
XFILLER_35_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16666_ _25996_/Q vssd1 vssd1 vccd1 vccd1 _20977_/A sky130_fd_sc_hd__clkbuf_4
X_19454_ _19454_/A _19454_/B vssd1 vssd1 vccd1 vccd1 _19454_/X sky130_fd_sc_hd__or2_1
X_13878_ _25836_/Q _26036_/Q _14008_/S vssd1 vssd1 vccd1 vccd1 _13878_/X sky130_fd_sc_hd__mux2_1
XFILLER_234_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15617_ _17838_/A _16043_/B vssd1 vssd1 vccd1 vccd1 _16621_/B sky130_fd_sc_hd__nor2_2
X_18405_ _18435_/A _18404_/X _18386_/B vssd1 vssd1 vccd1 vccd1 _18405_/X sky130_fd_sc_hd__a21o_1
XFILLER_201_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12829_ _12975_/A _12975_/B _25470_/Q vssd1 vssd1 vccd1 vccd1 _12981_/A sky130_fd_sc_hd__or3b_4
X_19385_ _19449_/A _19385_/B vssd1 vssd1 vccd1 vccd1 _19385_/Y sky130_fd_sc_hd__nand2_1
X_16597_ _16597_/A _16890_/A vssd1 vssd1 vccd1 vccd1 _16597_/X sky130_fd_sc_hd__or2_1
XFILLER_203_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15548_ _27280_/Q _26473_/Q _15548_/S vssd1 vssd1 vccd1 vccd1 _15548_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18336_ _18336_/A _18336_/B vssd1 vssd1 vccd1 vccd1 _18337_/A sky130_fd_sc_hd__and2_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18267_ _18263_/X _18266_/X _18487_/A vssd1 vssd1 vccd1 vccd1 _18267_/X sky130_fd_sc_hd__mux2_1
X_15479_ _13114_/A _15466_/X _15470_/X _15478_/X _13168_/A vssd1 vssd1 vccd1 vccd1
+ _15479_/X sky130_fd_sc_hd__a311o_1
XFILLER_129_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17218_ _17218_/A vssd1 vssd1 vccd1 vccd1 _17219_/A sky130_fd_sc_hd__buf_2
X_18198_ _18202_/A vssd1 vssd1 vccd1 vccd1 _18348_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_128_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17149_ _17149_/A vssd1 vssd1 vccd1 vccd1 _25477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20160_ _20160_/A _20160_/B vssd1 vssd1 vccd1 vccd1 _20160_/X sky130_fd_sc_hd__xor2_1
XFILLER_157_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20091_ _20091_/A vssd1 vssd1 vccd1 vccd1 _20355_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_257_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_257_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23850_ _23773_/X _26807_/Q _23854_/S vssd1 vssd1 vccd1 vccd1 _23851_/A sky130_fd_sc_hd__mux2_1
XFILLER_273_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22801_ _22801_/A vssd1 vssd1 vccd1 vccd1 _26384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23781_ _23781_/A vssd1 vssd1 vccd1 vccd1 _26777_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20993_ _23211_/A _25321_/B vssd1 vssd1 vccd1 vccd1 _21050_/A sky130_fd_sc_hd__nor2_8
XFILLER_214_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25520_ _27022_/CLK _25520_/D vssd1 vssd1 vccd1 vccd1 _25520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22732_ _22732_/A vssd1 vssd1 vccd1 vccd1 _26355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_281_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_53_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25451_ _23766_/X _27320_/Q _25459_/S vssd1 vssd1 vccd1 vccd1 _25452_/A sky130_fd_sc_hd__mux2_1
X_22663_ _23706_/A vssd1 vssd1 vccd1 vccd1 _22663_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24402_ _24408_/A _24923_/A vssd1 vssd1 vccd1 vccd1 _24402_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21614_ _21276_/A _21613_/X _21603_/X vssd1 vssd1 vccd1 vccd1 _21614_/Y sky130_fd_sc_hd__o21ai_1
X_25382_ _25382_/A vssd1 vssd1 vccd1 vccd1 _27289_/D sky130_fd_sc_hd__clkbuf_1
X_22594_ _22607_/A vssd1 vssd1 vccd1 vccd1 _22604_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_205_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27121_ _27122_/CLK _27121_/D vssd1 vssd1 vccd1 vccd1 _27121_/Q sky130_fd_sc_hd__dfxtp_4
X_24333_ _27002_/Q _24329_/B _24332_/Y vssd1 vssd1 vccd1 vccd1 _27002_/D sky130_fd_sc_hd__o21a_1
X_21545_ _21545_/A vssd1 vssd1 vccd1 vccd1 _21545_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27052_ _27062_/CLK _27052_/D vssd1 vssd1 vccd1 vccd1 _27052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24264_ _26978_/Q _24266_/C _24263_/Y vssd1 vssd1 vccd1 vccd1 _26978_/D sky130_fd_sc_hd__o21a_1
X_21476_ _21476_/A vssd1 vssd1 vccd1 vccd1 _21476_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26003_ _27269_/CLK _26003_/D vssd1 vssd1 vccd1 vccd1 _26003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23215_ _23215_/A vssd1 vssd1 vccd1 vccd1 _26552_/D sky130_fd_sc_hd__clkbuf_1
X_20427_ _20427_/A _20427_/B vssd1 vssd1 vccd1 vccd1 _20427_/X sky130_fd_sc_hd__xor2_1
X_24195_ _24216_/A _24195_/B vssd1 vssd1 vccd1 vccd1 _24195_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23146_ _26522_/Q _23044_/X _23150_/S vssd1 vssd1 vccd1 vccd1 _23147_/A sky130_fd_sc_hd__mux2_1
X_20358_ _19315_/A _20355_/X _20356_/Y _20357_/X vssd1 vssd1 vccd1 vccd1 _20399_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_161_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23077_ _26500_/Q _23076_/X _23083_/S vssd1 vssd1 vccd1 vccd1 _23078_/A sky130_fd_sc_hd__mux2_1
X_20289_ _20289_/A _20289_/B vssd1 vssd1 vccd1 vccd1 _20289_/Y sky130_fd_sc_hd__nand2_1
XTAP_5501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22028_ _22028_/A vssd1 vssd1 vccd1 vccd1 _26125_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26905_ _26905_/CLK _26905_/D vssd1 vssd1 vccd1 vccd1 _26905_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14850_ _27260_/Q _15026_/B vssd1 vssd1 vccd1 vccd1 _14850_/X sky130_fd_sc_hd__or2_1
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26836_ _26900_/CLK _26836_/D vssd1 vssd1 vccd1 vccd1 _26836_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _16728_/B vssd1 vssd1 vccd1 vccd1 _13801_/Y sky130_fd_sc_hd__inv_2
XFILLER_264_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14781_ _14747_/A _26906_/Q _26778_/Q _14767_/S _14773_/A vssd1 vssd1 vccd1 vccd1
+ _14781_/X sky130_fd_sc_hd__a221o_1
X_26767_ _27314_/CLK _26767_/D vssd1 vssd1 vccd1 vccd1 _26767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_251_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23979_ _26864_/Q _23574_/X _23987_/S vssd1 vssd1 vccd1 vccd1 _23980_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16520_ _16517_/X _16518_/X _16519_/X _14760_/X vssd1 vssd1 vccd1 vccd1 _16521_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_217_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13732_ _14713_/B _13730_/X _13731_/X _13144_/A vssd1 vssd1 vccd1 vccd1 _13732_/X
+ sky130_fd_sc_hd__a211o_1
X_25718_ _27321_/CLK _25718_/D vssd1 vssd1 vccd1 vccd1 _25718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26698_ _27278_/CLK _26698_/D vssd1 vssd1 vccd1 vccd1 _26698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16451_ _25751_/Q _16450_/Y _16451_/S vssd1 vssd1 vccd1 vccd1 _17780_/B sky130_fd_sc_hd__mux2_2
X_25649_ _25661_/CLK _25649_/D vssd1 vssd1 vccd1 vccd1 _25649_/Q sky130_fd_sc_hd__dfxtp_1
X_13663_ _26789_/Q _26433_/Q _15292_/A vssd1 vssd1 vccd1 vccd1 _13663_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15402_ _16104_/A vssd1 vssd1 vccd1 vccd1 _15417_/A sky130_fd_sc_hd__clkbuf_2
X_19170_ _25555_/Q _18825_/X _19169_/X _18829_/X _18830_/X vssd1 vssd1 vccd1 vccd1
+ _19170_/X sky130_fd_sc_hd__a221o_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16382_ _14859_/X _16379_/X _16381_/X _14649_/A vssd1 vssd1 vccd1 vccd1 _16382_/X
+ sky130_fd_sc_hd__a211o_1
X_13594_ _26073_/Q _15796_/S _15806_/S _13593_/X vssd1 vssd1 vccd1 vccd1 _13594_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_85_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26908_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18121_ _18121_/A _18121_/B vssd1 vssd1 vccd1 vccd1 _18823_/A sky130_fd_sc_hd__and2_2
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27319_ _27319_/CLK _27319_/D vssd1 vssd1 vccd1 vccd1 _27319_/Q sky130_fd_sc_hd__dfxtp_1
X_15333_ _15333_/A vssd1 vssd1 vccd1 vccd1 _15333_/X sky130_fd_sc_hd__clkbuf_4
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26796_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18052_ _17910_/X _17906_/X _18062_/S vssd1 vssd1 vccd1 vccd1 _18052_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15264_ _27285_/Q _26478_/Q _16325_/S vssd1 vssd1 vccd1 vccd1 _15264_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17003_ _17016_/A vssd1 vssd1 vccd1 vccd1 _17003_/X sky130_fd_sc_hd__buf_2
X_14215_ _26912_/Q _26396_/Q _14289_/S vssd1 vssd1 vccd1 vccd1 _14215_/X sky130_fd_sc_hd__mux2_1
X_15195_ _26676_/Q _25716_/Q _16428_/S vssd1 vssd1 vccd1 vccd1 _15195_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14146_ _25634_/Q _15443_/B _13578_/A _25602_/Q vssd1 vssd1 vccd1 vccd1 _14147_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_263_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14077_ _14077_/A _14077_/B _14077_/C vssd1 vssd1 vccd1 vccd1 _14077_/X sky130_fd_sc_hd__and3_1
X_18954_ _27053_/Q _19055_/A _18951_/X _18953_/X _19066_/A vssd1 vssd1 vccd1 vccd1
+ _18954_/X sky130_fd_sc_hd__o221a_1
XFILLER_267_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13028_ _13028_/A vssd1 vssd1 vccd1 vccd1 _15388_/A sky130_fd_sc_hd__buf_4
X_17905_ _17900_/X _17904_/X _18050_/S vssd1 vssd1 vccd1 vccd1 _17905_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18885_ _18723_/X _18882_/X _18883_/Y _18884_/X vssd1 vssd1 vccd1 vccd1 _18886_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17836_ _18941_/A _18941_/B _17836_/C vssd1 vssd1 vccd1 vccd1 _19109_/B sky130_fd_sc_hd__or3_1
XFILLER_67_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17767_ _14559_/X _13641_/B _19140_/A vssd1 vssd1 vccd1 vccd1 _17767_/X sky130_fd_sc_hd__mux2_1
XFILLER_207_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14979_ _19847_/A _15012_/S _14978_/Y vssd1 vssd1 vccd1 vccd1 _17851_/A sky130_fd_sc_hd__o21ai_2
XFILLER_207_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19506_ _25637_/Q _19510_/B vssd1 vssd1 vccd1 vccd1 _19506_/X sky130_fd_sc_hd__or2_1
XFILLER_208_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16718_ _22480_/A _16703_/X _16705_/X _18357_/A vssd1 vssd1 vccd1 vccd1 _16718_/X
+ sky130_fd_sc_hd__a22o_2
X_17698_ _17697_/A _21208_/B _17697_/Y vssd1 vssd1 vccd1 vccd1 _17745_/A sky130_fd_sc_hd__o21ai_2
XINSDIODE2_420 _17099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_431 _26236_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19437_ _27067_/Q _18747_/X _19434_/X _19436_/X _18761_/X vssd1 vssd1 vccd1 vccd1
+ _19437_/X sky130_fd_sc_hd__o221a_2
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_442 _25730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_453 _17059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16649_ _26940_/Q vssd1 vssd1 vccd1 vccd1 _24986_/A sky130_fd_sc_hd__clkbuf_8
XINSDIODE2_464 _19246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_475 _17653_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_486 _14886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19368_ _27033_/Q _18514_/A _19367_/X _18455_/A vssd1 vssd1 vccd1 vccd1 _19368_/X
+ sky130_fd_sc_hd__a22o_1
XINSDIODE2_497 _18483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18319_ _18270_/X _18318_/X _18349_/S vssd1 vssd1 vccd1 vccd1 _18683_/B sky130_fd_sc_hd__mux2_1
XFILLER_175_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19299_ _27225_/Q _19299_/B vssd1 vssd1 vccd1 vccd1 _19299_/X sky130_fd_sc_hd__and2_1
XFILLER_175_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21330_ _24871_/A vssd1 vssd1 vccd1 vccd1 _21330_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21261_ _21273_/A _21261_/B vssd1 vssd1 vccd1 vccd1 _21261_/Y sky130_fd_sc_hd__nor2_2
XFILLER_237_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23000_ _26472_/Q _22695_/X _23006_/S vssd1 vssd1 vccd1 vccd1 _23001_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20212_ _20206_/X _20208_/Y _20211_/X vssd1 vssd1 vccd1 vccd1 _20212_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_opt_5_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_21192_ input9/X _21070_/A _21065_/Y _21195_/A vssd1 vssd1 vccd1 vccd1 _21192_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_132_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20143_ _25742_/Q _20091_/A _20142_/Y _20115_/A vssd1 vssd1 vccd1 vccd1 _20144_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_131_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24951_ hold3/X _24951_/B vssd1 vssd1 vccd1 vccd1 _24951_/Y sky130_fd_sc_hd__nand2_1
X_20074_ _19649_/A _20071_/Y _20072_/X _20073_/X vssd1 vssd1 vccd1 vccd1 _20074_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_170_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23902_ _23744_/X _26830_/Q _23904_/S vssd1 vssd1 vccd1 vccd1 _23903_/A sky130_fd_sc_hd__mux2_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24882_ _20692_/A _19724_/X _25147_/A _24896_/B vssd1 vssd1 vccd1 vccd1 _24882_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_57_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26621_ _26813_/CLK _26621_/D vssd1 vssd1 vccd1 vccd1 _26621_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23833_ _23833_/A vssd1 vssd1 vccd1 vccd1 _26799_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26552_ _27295_/CLK _26552_/D vssd1 vssd1 vccd1 vccd1 _26552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23764_ _23763_/X _26772_/Q _23764_/S vssd1 vssd1 vccd1 vccd1 _23765_/A sky130_fd_sc_hd__mux2_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20976_ _21349_/B vssd1 vssd1 vccd1 vccd1 _20986_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_213_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25503_ _27014_/CLK _25503_/D vssd1 vssd1 vccd1 vccd1 _25503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22715_ _26350_/Q _22714_/X _22721_/S vssd1 vssd1 vccd1 vccd1 _22716_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26483_ _26483_/CLK _26483_/D vssd1 vssd1 vccd1 vccd1 _26483_/Q sky130_fd_sc_hd__dfxtp_1
X_23695_ _23695_/A vssd1 vssd1 vccd1 vccd1 _26750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25434_ _25434_/A vssd1 vssd1 vccd1 vccd1 _27312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22646_ _22646_/A vssd1 vssd1 vccd1 vccd1 _26328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25365_ _27282_/Q _23747_/A _25365_/S vssd1 vssd1 vccd1 vccd1 _25366_/A sky130_fd_sc_hd__mux2_1
X_22577_ _22567_/X _22576_/Y _22574_/X vssd1 vssd1 vccd1 vccd1 _26306_/D sky130_fd_sc_hd__a21oi_1
XFILLER_22_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27104_ _27110_/CLK _27104_/D vssd1 vssd1 vccd1 vccd1 _27104_/Q sky130_fd_sc_hd__dfxtp_2
X_24316_ _26996_/Q _24318_/C _24315_/Y vssd1 vssd1 vccd1 vccd1 _26996_/D sky130_fd_sc_hd__o21a_1
XFILLER_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21528_ _21528_/A vssd1 vssd1 vccd1 vccd1 _21528_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25296_ _23750_/X _27251_/Q _25304_/S vssd1 vssd1 vccd1 vccd1 _25297_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27035_ _27133_/CLK _27035_/D vssd1 vssd1 vccd1 vccd1 _27035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24247_ _26972_/Q _24250_/C _24246_/Y vssd1 vssd1 vccd1 vccd1 _26972_/D sky130_fd_sc_hd__o21a_1
XFILLER_147_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21459_ _21459_/A vssd1 vssd1 vccd1 vccd1 _21459_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14000_ _27301_/Q _26558_/Q _14004_/S vssd1 vssd1 vccd1 vccd1 _14000_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24178_ _26950_/Q _26949_/Q _24178_/C vssd1 vssd1 vccd1 vccd1 _24184_/C sky130_fd_sc_hd__and3_1
XFILLER_269_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23129_ _23129_/A vssd1 vssd1 vccd1 vccd1 _26516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_132_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27160_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_150_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15951_ _16631_/A vssd1 vssd1 vccd1 vccd1 _17816_/C sky130_fd_sc_hd__inv_2
XTAP_5331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput120 dout1[21] vssd1 vssd1 vccd1 vccd1 input120/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput131 dout1[31] vssd1 vssd1 vccd1 vccd1 input131/X sky130_fd_sc_hd__clkbuf_1
XFILLER_209_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput142 dout1[41] vssd1 vssd1 vccd1 vccd1 input142/X sky130_fd_sc_hd__clkbuf_2
X_14902_ _14890_/X _26713_/Q _26841_/Q _14984_/S _14773_/A vssd1 vssd1 vccd1 vccd1
+ _14902_/X sky130_fd_sc_hd__a221o_1
Xinput153 dout1[51] vssd1 vssd1 vccd1 vccd1 input153/X sky130_fd_sc_hd__buf_2
XTAP_5364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15882_ _26665_/Q _25705_/Q _15888_/S vssd1 vssd1 vccd1 vccd1 _15882_/X sky130_fd_sc_hd__mux2_1
X_18670_ _19253_/A vssd1 vssd1 vccd1 vccd1 _18973_/A sky130_fd_sc_hd__buf_2
XFILLER_102_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput164 dout1[61] vssd1 vssd1 vccd1 vccd1 input164/X sky130_fd_sc_hd__clkbuf_2
XTAP_5375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput175 irq[13] vssd1 vssd1 vccd1 vccd1 input175/X sky130_fd_sc_hd__buf_6
XTAP_5397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput186 irq[9] vssd1 vssd1 vccd1 vccd1 _19612_/C sky130_fd_sc_hd__buf_4
XFILLER_264_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _14706_/X _17612_/X _17608_/X _17620_/X vssd1 vssd1 vccd1 vccd1 _17622_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput197 localMemory_wb_adr_i[16] vssd1 vssd1 vccd1 vccd1 input197/X sky130_fd_sc_hd__clkbuf_1
X_26819_ _27304_/CLK _26819_/D vssd1 vssd1 vccd1 vccd1 _26819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14833_ _14833_/A vssd1 vssd1 vccd1 vccd1 _18785_/A sky130_fd_sc_hd__buf_2
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14764_ _14764_/A vssd1 vssd1 vccd1 vccd1 _14765_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17552_ _19650_/A vssd1 vssd1 vccd1 vccd1 _17608_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13715_ _13086_/X _26884_/Q _26756_/Q _16078_/S _13051_/A vssd1 vssd1 vccd1 vccd1
+ _13715_/X sky130_fd_sc_hd__a221o_1
XFILLER_32_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16503_ _16480_/S _16500_/X _16502_/X _14662_/X vssd1 vssd1 vccd1 vccd1 _16503_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_205_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17483_ _17682_/B vssd1 vssd1 vccd1 vccd1 _17483_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14695_ _16398_/S vssd1 vssd1 vccd1 vccd1 _16221_/S sky130_fd_sc_hd__buf_4
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19222_ _27093_/Q _18508_/A _18509_/A _27191_/Q _18510_/A vssd1 vssd1 vccd1 vccd1
+ _19222_/X sky130_fd_sc_hd__a221o_1
XFILLER_232_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13646_ _13779_/A _13639_/X _13645_/X _15932_/A vssd1 vssd1 vccd1 vccd1 _13646_/X
+ sky130_fd_sc_hd__a211o_1
X_16434_ _15406_/X _26711_/Q _26839_/Q _16443_/S _15210_/X vssd1 vssd1 vccd1 vccd1
+ _16434_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16365_ _14808_/A _16353_/X _16357_/X _16364_/X _16280_/S vssd1 vssd1 vccd1 vccd1
+ _16365_/X sky130_fd_sc_hd__a311o_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19153_ _19287_/B vssd1 vssd1 vccd1 vccd1 _19153_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_201_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ _13577_/A vssd1 vssd1 vccd1 vccd1 _13578_/A sky130_fd_sc_hd__clkbuf_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18104_ _18811_/A vssd1 vssd1 vccd1 vccd1 _19055_/A sky130_fd_sc_hd__buf_2
XFILLER_157_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15316_ _15111_/A _25780_/Q _16443_/S _26866_/Q _14729_/A vssd1 vssd1 vccd1 vccd1
+ _15316_/X sky130_fd_sc_hd__o221a_1
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19084_ _19448_/A _19045_/Y _19083_/X vssd1 vssd1 vccd1 vccd1 _19084_/Y sky130_fd_sc_hd__o21ai_4
X_16296_ _23590_/A vssd1 vssd1 vccd1 vccd1 _16296_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15247_ _25652_/Q _16212_/B vssd1 vssd1 vccd1 vccd1 _15247_/X sky130_fd_sc_hd__and2_1
X_18035_ _18035_/A _19290_/A vssd1 vssd1 vccd1 vccd1 _18035_/X sky130_fd_sc_hd__or2_1
XFILLER_274_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15178_ _16060_/S vssd1 vssd1 vccd1 vccd1 _16143_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_153_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14129_ _17800_/A vssd1 vssd1 vccd1 vccd1 _16717_/A sky130_fd_sc_hd__clkbuf_4
X_19986_ _22496_/A _20017_/C vssd1 vssd1 vccd1 vccd1 _19986_/Y sky130_fd_sc_hd__nor2_1
XFILLER_259_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18937_ _17967_/X _17918_/X _18364_/X _18269_/A vssd1 vssd1 vccd1 vccd1 _18940_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_228_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18868_ _27083_/Q _18751_/X _18752_/X _27181_/Q _18753_/X vssd1 vssd1 vccd1 vccd1
+ _18868_/X sky130_fd_sc_hd__a221o_1
XFILLER_255_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17819_ _13689_/A _17819_/B vssd1 vssd1 vccd1 vccd1 _18634_/A sky130_fd_sc_hd__and2b_1
XFILLER_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18799_ _18799_/A _18799_/B vssd1 vssd1 vccd1 vccd1 _18799_/Y sky130_fd_sc_hd__nand2_1
XFILLER_227_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20830_ _25811_/Q vssd1 vssd1 vccd1 vccd1 _20831_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20761_ _20571_/X _25777_/Q _20761_/S vssd1 vssd1 vccd1 vccd1 _20762_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_250 _16804_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_261 _25466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22500_ _22500_/A _22502_/B vssd1 vssd1 vccd1 vccd1 _22501_/A sky130_fd_sc_hd__and2_1
XFILLER_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_272 _18524_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_283 _25815_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23480_ _26671_/Q _23098_/X _23480_/S vssd1 vssd1 vccd1 vccd1 _23481_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_294 _25824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20692_ _20692_/A _20703_/B vssd1 vssd1 vccd1 vccd1 _20692_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22431_ _26197_/Q _22418_/X _22430_/X _22428_/X vssd1 vssd1 vccd1 vccd1 _26245_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25150_ _20694_/A _25138_/X _25149_/X vssd1 vssd1 vccd1 vccd1 _25150_/X sky130_fd_sc_hd__o21a_1
XFILLER_109_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22362_ _22387_/B _22362_/B vssd1 vssd1 vccd1 vccd1 _22362_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24101_ _26918_/Q _23542_/X _24109_/S vssd1 vssd1 vccd1 vccd1 _24102_/A sky130_fd_sc_hd__mux2_1
X_21313_ _21311_/X _21312_/X _21290_/X vssd1 vssd1 vccd1 vccd1 _21313_/X sky130_fd_sc_hd__a21o_1
XFILLER_248_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25081_ _20662_/A _25059_/X _25080_/X vssd1 vssd1 vccd1 vccd1 _25081_/Y sky130_fd_sc_hd__o21ai_1
X_22293_ _26210_/Q _22284_/X _22292_/X _22288_/X vssd1 vssd1 vccd1 vccd1 _26210_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24032_ _24032_/A vssd1 vssd1 vccd1 vccd1 _26887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21244_ _21244_/A _21244_/B vssd1 vssd1 vccd1 vccd1 _21275_/A sky130_fd_sc_hd__or2_1
XFILLER_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21175_ _25929_/Q _21166_/X _21167_/X input29/X vssd1 vssd1 vccd1 vccd1 _21176_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_104_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20126_ _20126_/A _20126_/B vssd1 vssd1 vccd1 vccd1 _20204_/B sky130_fd_sc_hd__nand2_1
X_25983_ _25985_/CLK _25983_/D vssd1 vssd1 vccd1 vccd1 _25983_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24934_ _24577_/A _24917_/X _24909_/X vssd1 vssd1 vccd1 vccd1 _24934_/Y sky130_fd_sc_hd__a21oi_1
X_20057_ _25739_/Q vssd1 vssd1 vccd1 vccd1 _20664_/A sky130_fd_sc_hd__buf_8
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_274_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24865_ _24863_/Y _24864_/X _24854_/X vssd1 vssd1 vccd1 vccd1 _27122_/D sky130_fd_sc_hd__a21oi_1
XFILLER_100_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23816_ _23816_/A vssd1 vssd1 vccd1 vccd1 _26791_/D sky130_fd_sc_hd__clkbuf_1
X_26604_ _26604_/CLK _26604_/D vssd1 vssd1 vccd1 vccd1 _26604_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24796_ _24835_/A vssd1 vssd1 vccd1 vccd1 _24796_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26535_ _27313_/CLK _26535_/D vssd1 vssd1 vccd1 vccd1 _26535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23747_ _23747_/A vssd1 vssd1 vccd1 vccd1 _23747_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_214_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20959_ _25856_/Q _20958_/X _20965_/S vssd1 vssd1 vccd1 vccd1 _20960_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13500_ _26662_/Q _25702_/Q _15408_/A vssd1 vssd1 vccd1 vccd1 _13500_/X sky130_fd_sc_hd__mux2_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26466_ _27277_/CLK _26466_/D vssd1 vssd1 vccd1 vccd1 _26466_/Q sky130_fd_sc_hd__dfxtp_1
X_14480_ _13464_/A _23514_/A _14479_/X _13212_/A vssd1 vssd1 vccd1 vccd1 _14480_/X
+ sky130_fd_sc_hd__o211a_4
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23678_ _26745_/Q _23603_/X _23678_/S vssd1 vssd1 vccd1 vccd1 _23679_/A sky130_fd_sc_hd__mux2_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13431_ _13431_/A vssd1 vssd1 vccd1 vccd1 _13431_/X sky130_fd_sc_hd__buf_2
X_25417_ _25463_/S vssd1 vssd1 vccd1 vccd1 _25426_/S sky130_fd_sc_hd__buf_6
XFILLER_13_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22629_ _22629_/A _26326_/Q vssd1 vssd1 vccd1 vccd1 _22638_/D sky130_fd_sc_hd__and2_1
XFILLER_201_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26397_ _27267_/CLK _26397_/D vssd1 vssd1 vccd1 vccd1 _26397_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_173_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16150_ _14622_/A _16137_/X _16141_/X _16149_/X _14682_/A vssd1 vssd1 vccd1 vccd1
+ _16150_/X sky130_fd_sc_hd__a311o_1
X_25348_ _27274_/Q _23722_/A _25354_/S vssd1 vssd1 vccd1 vccd1 _25349_/A sky130_fd_sc_hd__mux2_1
X_13362_ _15776_/A vssd1 vssd1 vccd1 vccd1 _13363_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15101_ _15085_/X _15096_/X _15100_/X _14803_/A vssd1 vssd1 vccd1 vccd1 _15101_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_166_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16081_ _14706_/A _16072_/X _16080_/X _14708_/A vssd1 vssd1 vccd1 vccd1 _16081_/X
+ sky130_fd_sc_hd__a211o_1
X_25279_ _25279_/A vssd1 vssd1 vccd1 vccd1 _27243_/D sky130_fd_sc_hd__clkbuf_1
X_13293_ _16261_/S vssd1 vssd1 vccd1 vccd1 _16342_/S sky130_fd_sc_hd__buf_4
XFILLER_182_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27018_ _27022_/CLK _27018_/D vssd1 vssd1 vccd1 vccd1 _27018_/Q sky130_fd_sc_hd__dfxtp_1
X_15032_ _16308_/S vssd1 vssd1 vccd1 vccd1 _16241_/S sky130_fd_sc_hd__buf_4
XFILLER_6_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19840_ _19814_/Y _19819_/B _19816_/B vssd1 vssd1 vccd1 vccd1 _19841_/B sky130_fd_sc_hd__o21ai_1
XFILLER_218_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19771_ _19771_/A vssd1 vssd1 vccd1 vccd1 _19771_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16983_ _16983_/A _16983_/B _16983_/C vssd1 vssd1 vccd1 vccd1 _16983_/X sky130_fd_sc_hd__and3_1
XFILLER_256_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18722_ _19252_/A vssd1 vssd1 vccd1 vccd1 _18967_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15934_ _13351_/A _26697_/Q _26825_/Q _15197_/A _13363_/A vssd1 vssd1 vccd1 vccd1
+ _15934_/X sky130_fd_sc_hd__a221o_1
XTAP_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18653_ _27209_/Q _19258_/B vssd1 vssd1 vccd1 vccd1 _18653_/X sky130_fd_sc_hd__and2_1
XFILLER_64_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15865_ _15853_/X _15856_/X _15864_/Y vssd1 vssd1 vccd1 vccd1 _15865_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_225_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17604_ _19636_/A vssd1 vssd1 vccd1 vccd1 _17604_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_280_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14816_ _14816_/A vssd1 vssd1 vccd1 vccd1 _14817_/A sky130_fd_sc_hd__buf_6
X_18584_ _18340_/A _18541_/A _18553_/X _18583_/X vssd1 vssd1 vccd1 vccd1 _18584_/X
+ sky130_fd_sc_hd__a211o_1
X_15796_ _27309_/Q _26566_/Q _15796_/S vssd1 vssd1 vccd1 vccd1 _15796_/X sky130_fd_sc_hd__mux2_1
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17535_ _17597_/A vssd1 vssd1 vccd1 vccd1 _17554_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_233_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14747_ _14747_/A vssd1 vssd1 vccd1 vccd1 _16513_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17466_ _26252_/Q _17453_/A _17460_/A _25980_/Q vssd1 vssd1 vccd1 vccd1 _17701_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_177_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14678_ _14678_/A vssd1 vssd1 vccd1 vccd1 _14679_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_220_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19205_ _25556_/Q _18568_/X _19204_/X _19069_/X _18572_/X vssd1 vssd1 vccd1 vccd1
+ _19205_/X sky130_fd_sc_hd__a221o_1
X_13629_ _15818_/S _13627_/X _13628_/X _13614_/A vssd1 vssd1 vccd1 vccd1 _13629_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16417_ _17780_/A vssd1 vssd1 vccd1 vccd1 _16453_/A sky130_fd_sc_hd__inv_2
XFILLER_158_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17397_ _17395_/X _17399_/C _17396_/Y vssd1 vssd1 vccd1 vccd1 _25550_/D sky130_fd_sc_hd__o21a_1
XFILLER_220_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19136_ _26962_/Q _18569_/X _18570_/X _26994_/Q vssd1 vssd1 vccd1 vccd1 _19136_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16348_ _16346_/X _16347_/X _16348_/S vssd1 vssd1 vccd1 vccd1 _16348_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19067_ _27056_/Q _19055_/X _19062_/X _19065_/X _19066_/X vssd1 vssd1 vccd1 vccd1
+ _19067_/X sky130_fd_sc_hd__o221a_2
X_16279_ _16269_/X _16272_/X _16275_/X _16278_/X _14758_/A _14778_/A vssd1 vssd1 vccd1
+ vccd1 _16279_/X sky130_fd_sc_hd__mux4_2
XFILLER_218_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput402 _17010_/X vssd1 vssd1 vccd1 vccd1 din0[4] sky130_fd_sc_hd__buf_2
XFILLER_172_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18018_ _19910_/A vssd1 vssd1 vccd1 vccd1 _20141_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput413 _25948_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[12] sky130_fd_sc_hd__buf_2
Xoutput424 _25958_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[22] sky130_fd_sc_hd__buf_2
Xoutput435 _25939_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[3] sky130_fd_sc_hd__buf_2
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput446 _26233_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[1] sky130_fd_sc_hd__buf_2
XFILLER_126_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput457 _25740_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[16] sky130_fd_sc_hd__buf_2
XFILLER_259_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput468 _25750_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[26] sky130_fd_sc_hd__buf_2
Xoutput479 _25731_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[7] sky130_fd_sc_hd__buf_2
XFILLER_271_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19969_ _17992_/A _19914_/X _19774_/B _20089_/A vssd1 vssd1 vccd1 vccd1 _20006_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22980_ _26463_/Q _22666_/X _22984_/S vssd1 vssd1 vccd1 vccd1 _22981_/A sky130_fd_sc_hd__mux2_1
XFILLER_255_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21931_ _20567_/X _26082_/Q _21933_/S vssd1 vssd1 vccd1 vccd1 _21932_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24650_ _19634_/C _24636_/A _24649_/Y _21597_/A vssd1 vssd1 vccd1 vccd1 _24650_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21862_ _26059_/Q _20967_/X _21864_/S vssd1 vssd1 vccd1 vccd1 _21863_/A sky130_fd_sc_hd__mux2_1
XFILLER_270_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23601_ _26712_/Q _23600_/X _23604_/S vssd1 vssd1 vccd1 vccd1 _23602_/A sky130_fd_sc_hd__mux2_1
X_20813_ _20813_/A vssd1 vssd1 vccd1 vccd1 _25802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24581_ _27048_/Q _24576_/X _24579_/Y _24580_/X vssd1 vssd1 vccd1 vccd1 _27048_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_270_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21793_ _21793_/A _21793_/B vssd1 vssd1 vccd1 vccd1 _22962_/A sky130_fd_sc_hd__nand2_8
XFILLER_23_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26320_ _26326_/CLK _26320_/D vssd1 vssd1 vccd1 vccd1 _26320_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23532_ _23532_/A vssd1 vssd1 vccd1 vccd1 _26690_/D sky130_fd_sc_hd__clkbuf_1
X_20744_ _20538_/X _25769_/Q _20750_/S vssd1 vssd1 vccd1 vccd1 _20745_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26251_ _26307_/CLK _26251_/D vssd1 vssd1 vccd1 vccd1 _26251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23463_ _26663_/Q _23073_/X _23469_/S vssd1 vssd1 vccd1 vccd1 _23464_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20675_ _20675_/A _20683_/B vssd1 vssd1 vccd1 vccd1 _20675_/X sky130_fd_sc_hd__or2_1
XFILLER_177_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25202_ _24696_/B _25198_/X _25196_/X _27212_/Q _25199_/X vssd1 vssd1 vccd1 vccd1
+ _27212_/D sky130_fd_sc_hd__o221a_1
X_22414_ _26325_/Q vssd1 vssd1 vccd1 vccd1 _22638_/A sky130_fd_sc_hd__clkbuf_2
X_26182_ _26319_/CLK _26182_/D vssd1 vssd1 vccd1 vccd1 _26182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23394_ _23394_/A vssd1 vssd1 vccd1 vccd1 _26632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25133_ _22522_/A _25119_/X _25114_/X _19252_/B _25024_/A vssd1 vssd1 vccd1 vccd1
+ _25133_/X sky130_fd_sc_hd__a221o_1
X_22345_ _22335_/Y _22343_/X _22344_/X _22330_/X vssd1 vssd1 vccd1 vccd1 _26227_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25064_ _27177_/Q _25058_/X _25063_/X vssd1 vssd1 vccd1 vccd1 _27177_/D sky130_fd_sc_hd__o21ba_1
XFILLER_124_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22276_ _26204_/Q _22269_/X _22275_/X _22273_/X vssd1 vssd1 vccd1 vccd1 _26204_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24015_ _26880_/Q _23523_/X _24015_/S vssd1 vssd1 vccd1 vccd1 _24016_/A sky130_fd_sc_hd__mux2_1
X_21227_ _21407_/A vssd1 vssd1 vccd1 vccd1 _21227_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21158_ _21172_/A _21158_/B vssd1 vssd1 vccd1 vccd1 _21159_/A sky130_fd_sc_hd__or2_1
XFILLER_78_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20109_ _19993_/X _20106_/X _20131_/B _20108_/Y vssd1 vssd1 vccd1 vccd1 _20109_/X
+ sky130_fd_sc_hd__o31a_2
X_13980_ _25730_/Q _14317_/B vssd1 vssd1 vccd1 vccd1 _13980_/X sky130_fd_sc_hd__or2_1
XFILLER_77_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25966_ _27000_/CLK _25966_/D vssd1 vssd1 vccd1 vccd1 _25966_/Q sky130_fd_sc_hd__dfxtp_1
X_21089_ _21100_/A _21089_/B vssd1 vssd1 vccd1 vccd1 _21090_/A sky130_fd_sc_hd__or2_1
XFILLER_247_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12931_ _15791_/A _16409_/A _14604_/B _12930_/X vssd1 vssd1 vccd1 vccd1 _12931_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24917_ _24954_/A vssd1 vssd1 vccd1 vccd1 _24917_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25897_ _27292_/CLK _25897_/D vssd1 vssd1 vccd1 vccd1 _25897_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12862_ _12862_/A vssd1 vssd1 vccd1 vccd1 _13569_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _12772_/A _26892_/Q _26764_/Q _15540_/S vssd1 vssd1 vccd1 vccd1 _15650_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24848_ _24848_/A vssd1 vssd1 vccd1 vccd1 _24848_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _14601_/A vssd1 vssd1 vccd1 vccd1 _14601_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15581_ _15581_/A _15581_/B vssd1 vssd1 vccd1 vccd1 _15581_/Y sky130_fd_sc_hd__nor2_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24779_ _24779_/A vssd1 vssd1 vccd1 vccd1 _24798_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _13269_/A _25577_/Q vssd1 vssd1 vccd1 vccd1 _17162_/A sky130_fd_sc_hd__nand2_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _17317_/X _17322_/C _17319_/Y vssd1 vssd1 vccd1 vccd1 _25526_/D sky130_fd_sc_hd__o21a_1
X_14532_ _26620_/Q _26716_/Q _14539_/S vssd1 vssd1 vccd1 vccd1 _14532_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26518_ _27293_/CLK _26518_/D vssd1 vssd1 vccd1 vccd1 _26518_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _13311_/A _14451_/X _14455_/X _14462_/X vssd1 vssd1 vccd1 vccd1 _14463_/X
+ sky130_fd_sc_hd__a31o_1
X_17251_ _25505_/Q _17253_/C _20973_/A vssd1 vssd1 vccd1 vccd1 _17252_/B sky130_fd_sc_hd__o21ai_1
X_26449_ _27259_/CLK _26449_/D vssd1 vssd1 vccd1 vccd1 _26449_/Q sky130_fd_sc_hd__dfxtp_1
X_13414_ _12771_/A _26402_/Q _13410_/X _13413_/X vssd1 vssd1 vccd1 vccd1 _13414_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16202_ _14723_/A _16133_/Y _16201_/Y _14827_/A vssd1 vssd1 vccd1 vccd1 _19141_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17182_ _25487_/Q _17159_/X _17181_/Y _17175_/X vssd1 vssd1 vccd1 vccd1 _25487_/D
+ sky130_fd_sc_hd__o211a_1
X_14394_ _13939_/A _14390_/X _14393_/X _14542_/A vssd1 vssd1 vccd1 vccd1 _14394_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_168_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16133_ _23578_/A vssd1 vssd1 vccd1 vccd1 _16133_/Y sky130_fd_sc_hd__inv_2
X_13345_ _13512_/A vssd1 vssd1 vccd1 vccd1 _13346_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16064_ _15538_/X _16059_/X _16063_/X _14677_/A vssd1 vssd1 vccd1 vccd1 _16064_/X
+ sky130_fd_sc_hd__o211a_1
X_13276_ _13276_/A _13276_/B vssd1 vssd1 vccd1 vccd1 _13276_/Y sky130_fd_sc_hd__nor2_1
X_15015_ _16320_/S vssd1 vssd1 vccd1 vccd1 _15060_/S sky130_fd_sc_hd__buf_2
XFILLER_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19823_ _19823_/A _19803_/B vssd1 vssd1 vccd1 vccd1 _19830_/A sky130_fd_sc_hd__or2b_1
XFILLER_64_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_12_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25501_/CLK
+ sky130_fd_sc_hd__clkbuf_4
X_19754_ _19753_/Y _27137_/Q _19820_/S vssd1 vssd1 vccd1 vccd1 _19754_/X sky130_fd_sc_hd__mux2_2
XFILLER_231_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16966_ _16966_/A vssd1 vssd1 vccd1 vccd1 _16966_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_204_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18705_ _18705_/A vssd1 vssd1 vccd1 vccd1 _18705_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_238_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15917_ _13335_/A _15914_/X _15916_/X _13762_/X vssd1 vssd1 vccd1 vccd1 _15921_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_253_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19685_ _19686_/A _19686_/B vssd1 vssd1 vccd1 vccd1 _19687_/A sky130_fd_sc_hd__nor2_1
XFILLER_209_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16897_ _16955_/B _16848_/B _16847_/Y _16868_/A _16939_/B vssd1 vssd1 vccd1 vccd1
+ _16897_/X sky130_fd_sc_hd__o221a_1
XFILLER_225_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18636_ _18636_/A vssd1 vssd1 vccd1 vccd1 _18636_/X sky130_fd_sc_hd__buf_2
XFILLER_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15848_ _15844_/X _15847_/X _14816_/A vssd1 vssd1 vccd1 vccd1 _15848_/X sky130_fd_sc_hd__o21a_1
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18567_ _27045_/Q _18503_/X _18562_/X _18566_/X _18519_/X vssd1 vssd1 vccd1 vccd1
+ _18567_/X sky130_fd_sc_hd__o221a_1
XFILLER_91_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15779_ _13488_/A _26859_/Q _25773_/Q _15485_/S _15776_/A vssd1 vssd1 vccd1 vccd1
+ _15779_/X sky130_fd_sc_hd__a221o_1
XFILLER_52_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17518_ _25794_/Q vssd1 vssd1 vccd1 vccd1 _17518_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18498_ _18368_/X _18371_/X _18498_/S vssd1 vssd1 vccd1 vccd1 _18498_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17449_ _26327_/Q _26326_/Q vssd1 vssd1 vccd1 vccd1 _22415_/A sky130_fd_sc_hd__or2_2
XFILLER_32_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20460_ _20460_/A _20460_/B vssd1 vssd1 vccd1 vccd1 _20460_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_174_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19119_ _17444_/C _18890_/X _19117_/Y _19118_/X _18933_/X vssd1 vssd1 vccd1 vccd1
+ _19119_/X sky130_fd_sc_hd__a221o_4
XFILLER_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20391_ _20391_/A _20391_/B vssd1 vssd1 vccd1 vccd1 _20391_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_118_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22130_ _22130_/A vssd1 vssd1 vccd1 vccd1 _24441_/A sky130_fd_sc_hd__buf_4
XFILLER_118_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22061_ _22061_/A vssd1 vssd1 vccd1 vccd1 _26139_/D sky130_fd_sc_hd__clkbuf_1
X_21012_ _21012_/A vssd1 vssd1 vccd1 vccd1 _25876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput287 _17065_/X vssd1 vssd1 vccd1 vccd1 addr0[2] sky130_fd_sc_hd__buf_2
XFILLER_87_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput298 _16995_/X vssd1 vssd1 vccd1 vccd1 addr1[4] sky130_fd_sc_hd__buf_2
XFILLER_99_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_5 _22368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25820_ _26715_/CLK _25820_/D vssd1 vssd1 vccd1 vccd1 _25820_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_275_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25751_ _26292_/CLK _25751_/D vssd1 vssd1 vccd1 vccd1 _25751_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22963_ _23019_/A vssd1 vssd1 vccd1 vccd1 _23032_/S sky130_fd_sc_hd__buf_6
XFILLER_55_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_261_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21914_ _20533_/X _26074_/Q _21922_/S vssd1 vssd1 vccd1 vccd1 _21915_/A sky130_fd_sc_hd__mux2_1
X_24702_ _24944_/A vssd1 vssd1 vccd1 vccd1 _24703_/B sky130_fd_sc_hd__clkinv_2
X_25682_ _26286_/CLK _25682_/D vssd1 vssd1 vccd1 vccd1 _25682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22894_ _22894_/A vssd1 vssd1 vccd1 vccd1 _26424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24633_ _24900_/C _25206_/C _24633_/C _24341_/A vssd1 vssd1 vccd1 vccd1 _24740_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_55_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21845_ _26051_/Q _20942_/X _21849_/S vssd1 vssd1 vccd1 vccd1 _21846_/A sky130_fd_sc_hd__mux2_1
XFILLER_254_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24564_ _27042_/Q _24562_/X _24563_/Y _24551_/X vssd1 vssd1 vccd1 vccd1 _27042_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21776_ _20592_/X _26021_/Q _21776_/S vssd1 vssd1 vccd1 vccd1 _21777_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26303_ _26307_/CLK _26303_/D vssd1 vssd1 vccd1 vccd1 _26303_/Q sky130_fd_sc_hd__dfxtp_2
X_23515_ _26685_/Q _23514_/X _23524_/S vssd1 vssd1 vccd1 vccd1 _23516_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20727_ _20727_/A vssd1 vssd1 vccd1 vccd1 _25761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27283_ _27283_/CLK _27283_/D vssd1 vssd1 vccd1 vccd1 _27283_/Q sky130_fd_sc_hd__dfxtp_1
X_24495_ _26316_/Q _24473_/X _24474_/X input230/X _24384_/X vssd1 vssd1 vccd1 vccd1
+ _24495_/X sky130_fd_sc_hd__a221o_2
XFILLER_157_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26234_ _26297_/CLK _26234_/D vssd1 vssd1 vccd1 vccd1 _26234_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_196_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23446_ _23446_/A vssd1 vssd1 vccd1 vccd1 _26655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20658_ _21878_/A vssd1 vssd1 vccd1 vccd1 _20658_/X sky130_fd_sc_hd__buf_2
X_26165_ _27264_/CLK _26165_/D vssd1 vssd1 vccd1 vccd1 _26165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23377_ _23434_/S vssd1 vssd1 vccd1 vccd1 _23386_/S sky130_fd_sc_hd__buf_2
XFILLER_164_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20589_ _20588_/X _25715_/Q _20593_/S vssd1 vssd1 vccd1 vccd1 _20590_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13130_ _26855_/Q _25769_/Q _15540_/S vssd1 vssd1 vccd1 vccd1 _13130_/X sky130_fd_sc_hd__mux2_1
X_25116_ _20677_/A _25113_/X _25115_/X vssd1 vssd1 vccd1 vccd1 _25116_/Y sky130_fd_sc_hd__o21ai_1
X_22328_ _26222_/Q _22315_/X _22327_/X _22319_/X vssd1 vssd1 vccd1 vccd1 _26222_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26096_ _27264_/CLK _26096_/D vssd1 vssd1 vccd1 vccd1 _26096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13061_ _25840_/Q _26040_/Q _15557_/S vssd1 vssd1 vccd1 vccd1 _13061_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25047_ _27174_/Q _25030_/X _25046_/X vssd1 vssd1 vccd1 vccd1 _27174_/D sky130_fd_sc_hd__o21ba_1
X_22259_ _26198_/Q _22254_/X _22257_/X _22258_/X vssd1 vssd1 vccd1 vccd1 _26198_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_39_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27308_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_78_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16820_ _16838_/A _16820_/B vssd1 vssd1 vccd1 vccd1 _16862_/B sky130_fd_sc_hd__nor2_4
XFILLER_94_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26998_ _27001_/CLK _26998_/D vssd1 vssd1 vccd1 vccd1 _26998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16751_ _16751_/A vssd1 vssd1 vccd1 vccd1 _18968_/B sky130_fd_sc_hd__clkbuf_4
X_13963_ _13521_/A _25764_/Q _14365_/S _26850_/Q _13244_/A vssd1 vssd1 vccd1 vccd1
+ _13963_/X sky130_fd_sc_hd__o221a_1
X_25949_ _25985_/CLK _25949_/D vssd1 vssd1 vccd1 vccd1 _25949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15702_ _15702_/A vssd1 vssd1 vccd1 vccd1 _15703_/B sky130_fd_sc_hd__inv_2
X_19470_ _17336_/X _18746_/X _19467_/X _19469_/X _18770_/X vssd1 vssd1 vccd1 vccd1
+ _19470_/X sky130_fd_sc_hd__o221a_1
X_12914_ _13916_/A _13923_/B _13397_/B vssd1 vssd1 vccd1 vccd1 _15345_/A sky130_fd_sc_hd__or3_1
XFILLER_47_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13894_ _13890_/X _26883_/Q _26755_/Q _15980_/S vssd1 vssd1 vccd1 vccd1 _13894_/X
+ sky130_fd_sc_hd__a22o_1
X_16682_ _16678_/Y _16679_/X _16681_/Y vssd1 vssd1 vccd1 vccd1 _16682_/X sky130_fd_sc_hd__a21o_1
XFILLER_262_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18421_ _18495_/A _18421_/B vssd1 vssd1 vccd1 vccd1 _18421_/Y sky130_fd_sc_hd__nor2_1
XFILLER_222_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12845_ input168/X input139/X _25868_/Q vssd1 vssd1 vccd1 vccd1 _12846_/B sky130_fd_sc_hd__mux2_8
X_15633_ _15631_/X _15632_/X _15633_/S vssd1 vssd1 vccd1 vccd1 _15633_/X sky130_fd_sc_hd__mux2_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _18495_/A _18352_/B vssd1 vssd1 vccd1 vccd1 _18352_/Y sky130_fd_sc_hd__nor2_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _16071_/S _15563_/X _13071_/A vssd1 vssd1 vccd1 vccd1 _15564_/X sky130_fd_sc_hd__a21o_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _12776_/A vssd1 vssd1 vccd1 vccd1 _12777_/A sky130_fd_sc_hd__buf_2
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _25520_/Q _25521_/Q _17303_/C vssd1 vssd1 vccd1 vccd1 _17305_/B sky130_fd_sc_hd__and3_1
XFILLER_14_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ _14513_/X _14514_/X _14515_/S vssd1 vssd1 vccd1 vccd1 _14515_/X sky130_fd_sc_hd__mux2_1
X_15495_ _15495_/A _15495_/B vssd1 vssd1 vccd1 vccd1 _15495_/Y sky130_fd_sc_hd__nor2_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18283_ _18336_/A _18283_/B vssd1 vssd1 vccd1 vccd1 _18284_/A sky130_fd_sc_hd__and2_1
XFILLER_159_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17234_ _24208_/A vssd1 vssd1 vccd1 vccd1 _17414_/A sky130_fd_sc_hd__buf_2
X_14446_ _15376_/S _14362_/B _14444_/X _14445_/X vssd1 vssd1 vccd1 vccd1 _18059_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_266_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14377_ _13644_/A _14375_/X _14376_/X _13277_/A vssd1 vssd1 vccd1 vccd1 _14377_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_155_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17165_ _25481_/Q _17159_/X _17164_/X _17134_/X vssd1 vssd1 vccd1 vccd1 _25481_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13328_ _13358_/A vssd1 vssd1 vccd1 vccd1 _15769_/A sky130_fd_sc_hd__buf_2
XFILLER_115_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16116_ _15301_/S _16114_/X _16115_/X _13367_/X vssd1 vssd1 vccd1 vccd1 _16117_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_127_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17096_ _26240_/Q _26239_/Q vssd1 vssd1 vccd1 vccd1 _22406_/B sky130_fd_sc_hd__or2b_1
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13259_ _14308_/S vssd1 vssd1 vccd1 vccd1 _15938_/S sky130_fd_sc_hd__clkbuf_4
X_16047_ _14600_/A _16045_/Y _16046_/X _15135_/A vssd1 vssd1 vccd1 vccd1 _16047_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_143_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19806_ _19777_/A _19777_/B _19804_/X _19805_/X vssd1 vssd1 vccd1 vccd1 _19808_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_269_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17998_ _17998_/A _19393_/B vssd1 vssd1 vccd1 vccd1 _17998_/Y sky130_fd_sc_hd__nand2_1
XFILLER_215_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19737_ _19737_/A _19777_/B vssd1 vssd1 vccd1 vccd1 _19737_/X sky130_fd_sc_hd__or2_1
XFILLER_284_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16949_ _16986_/A _16949_/B vssd1 vssd1 vccd1 vccd1 _16950_/A sky130_fd_sc_hd__and2_1
XFILLER_272_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19668_ _19727_/A vssd1 vssd1 vccd1 vccd1 _19708_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_225_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18619_ _26950_/Q _18461_/A _18463_/A _26982_/Q vssd1 vssd1 vccd1 vccd1 _18619_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_253_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19599_ _14480_/X _18032_/Y _20227_/B vssd1 vssd1 vccd1 vccd1 _19658_/A sky130_fd_sc_hd__mux2_2
XFILLER_253_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21630_ _21630_/A _21641_/B vssd1 vssd1 vccd1 vccd1 _21630_/Y sky130_fd_sc_hd__nand2_1
XFILLER_212_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21561_ _21559_/X _21560_/X _21290_/A vssd1 vssd1 vccd1 vccd1 _21561_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23300_ _20504_/X _26591_/Q _23302_/S vssd1 vssd1 vccd1 vccd1 _23301_/A sky130_fd_sc_hd__mux2_1
X_20512_ _23702_/A vssd1 vssd1 vccd1 vccd1 _20512_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_24280_ _26983_/Q _24278_/B _24279_/Y vssd1 vssd1 vccd1 vccd1 _26983_/D sky130_fd_sc_hd__o21a_1
X_21492_ _21556_/A vssd1 vssd1 vccd1 vccd1 _21492_/X sky130_fd_sc_hd__buf_4
XFILLER_147_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23231_ _26560_/Q _23063_/X _23233_/S vssd1 vssd1 vccd1 vccd1 _23232_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20443_ _20427_/B _20443_/B _20443_/C vssd1 vssd1 vccd1 vccd1 _20450_/A sky130_fd_sc_hd__nand3b_1
XFILLER_119_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23162_ _23162_/A vssd1 vssd1 vccd1 vccd1 _26529_/D sky130_fd_sc_hd__clkbuf_1
X_20374_ _20470_/A _20399_/A _20362_/A vssd1 vssd1 vccd1 vccd1 _20380_/A sky130_fd_sc_hd__a21bo_1
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22113_ _22310_/A vssd1 vssd1 vccd1 vccd1 _22113_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23093_ _26505_/Q _23092_/X _23099_/S vssd1 vssd1 vccd1 vccd1 _23094_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22044_ _26132_/Q _20884_/X _22044_/S vssd1 vssd1 vccd1 vccd1 _22045_/A sky130_fd_sc_hd__mux2_1
X_26921_ _27308_/CLK _26921_/D vssd1 vssd1 vccd1 vccd1 _26921_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26852_ _26916_/CLK _26852_/D vssd1 vssd1 vccd1 vccd1 _26852_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25803_ _26520_/CLK _25803_/D vssd1 vssd1 vccd1 vccd1 _25803_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_229_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26783_ _27298_/CLK _26783_/D vssd1 vssd1 vccd1 vccd1 _26783_/Q sky130_fd_sc_hd__dfxtp_1
X_23995_ _23995_/A vssd1 vssd1 vccd1 vccd1 _26871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22946_ _22946_/A vssd1 vssd1 vccd1 vccd1 _26448_/D sky130_fd_sc_hd__clkbuf_1
X_25734_ _26271_/CLK _25734_/D vssd1 vssd1 vccd1 vccd1 _25734_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25665_ _26264_/CLK _25665_/D vssd1 vssd1 vccd1 vccd1 _25665_/Q sky130_fd_sc_hd__dfxtp_1
X_22877_ _22877_/A vssd1 vssd1 vccd1 vccd1 _26417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21828_ _21828_/A vssd1 vssd1 vccd1 vccd1 _26043_/D sky130_fd_sc_hd__clkbuf_1
X_24616_ _24972_/A _24621_/B vssd1 vssd1 vccd1 vccd1 _24616_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_157_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27198_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25596_ _25596_/CLK _25596_/D vssd1 vssd1 vccd1 vccd1 _25596_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24547_ _24561_/A vssd1 vssd1 vccd1 vccd1 _24553_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_54_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21759_ _20559_/X _26013_/Q _21765_/S vssd1 vssd1 vccd1 vccd1 _21760_/A sky130_fd_sc_hd__mux2_1
XPHY_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14300_ _27298_/Q _26555_/Q _14308_/S vssd1 vssd1 vccd1 vccd1 _14300_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15280_ _25851_/Q _26051_/Q _16315_/S vssd1 vssd1 vccd1 vccd1 _15280_/X sky130_fd_sc_hd__mux2_1
X_27266_ _27266_/CLK _27266_/D vssd1 vssd1 vccd1 vccd1 _27266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24478_ _24492_/A _24600_/A vssd1 vssd1 vccd1 vccd1 _24478_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14231_ _13638_/X _23523_/A _14230_/X _13683_/X vssd1 vssd1 vccd1 vccd1 _19728_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_156_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26217_ _26319_/CLK _26217_/D vssd1 vssd1 vccd1 vccd1 _26217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23429_ _23429_/A vssd1 vssd1 vccd1 vccd1 _26648_/D sky130_fd_sc_hd__clkbuf_1
X_27197_ _27198_/CLK _27197_/D vssd1 vssd1 vccd1 vccd1 _27197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14162_ _26624_/Q _26720_/Q _15904_/S vssd1 vssd1 vccd1 vccd1 _14162_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26148_ _26610_/CLK _26148_/D vssd1 vssd1 vccd1 vccd1 _26148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13113_ _14713_/A vssd1 vssd1 vccd1 vccd1 _13114_/A sky130_fd_sc_hd__clkbuf_4
X_26079_ _27278_/CLK _26079_/D vssd1 vssd1 vccd1 vccd1 _26079_/Q sky130_fd_sc_hd__dfxtp_1
X_14093_ _14268_/S _14093_/B vssd1 vssd1 vccd1 vccd1 _14093_/X sky130_fd_sc_hd__or2_1
X_18970_ _25614_/Q _18719_/X _18969_/X _18790_/X vssd1 vssd1 vccd1 vccd1 _25614_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_180_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13044_ _15459_/S vssd1 vssd1 vccd1 vccd1 _15566_/S sky130_fd_sc_hd__buf_2
X_17921_ _17950_/S vssd1 vssd1 vccd1 vccd1 _18681_/A sky130_fd_sc_hd__buf_2
XFILLER_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17852_ _17852_/A _17852_/B vssd1 vssd1 vccd1 vccd1 _17852_/Y sky130_fd_sc_hd__nor2_1
XFILLER_182_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16803_ _16838_/A _16910_/A _16589_/B _16597_/A vssd1 vssd1 vccd1 vccd1 _16803_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17783_ _17783_/A vssd1 vssd1 vccd1 vccd1 _17784_/B sky130_fd_sc_hd__inv_2
XFILLER_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14995_ _27323_/Q _26580_/Q _14996_/S vssd1 vssd1 vccd1 vccd1 _14995_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19522_ _19512_/X _18834_/X _19521_/X _19515_/X vssd1 vssd1 vccd1 vccd1 _25643_/D
+ sky130_fd_sc_hd__o211a_1
X_16734_ _25670_/Q vssd1 vssd1 vccd1 vccd1 _22491_/A sky130_fd_sc_hd__buf_4
X_13946_ _13941_/X _13942_/X _13944_/X _13945_/X vssd1 vssd1 vccd1 vccd1 _13947_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19453_ _19582_/B _25166_/A _19453_/S vssd1 vssd1 vccd1 vccd1 _19453_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16665_ _25981_/Q _16662_/X _21562_/B vssd1 vssd1 vccd1 vccd1 _16673_/A sky130_fd_sc_hd__o21a_1
XFILLER_207_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13877_ _14713_/A _13858_/X _13864_/X _13875_/X _13876_/X vssd1 vssd1 vccd1 vccd1
+ _13877_/X sky130_fd_sc_hd__a311o_1
XFILLER_222_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18404_ _18555_/A _18387_/X _18403_/X vssd1 vssd1 vccd1 vccd1 _18404_/X sky130_fd_sc_hd__a21o_4
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15616_ _16620_/B vssd1 vssd1 vccd1 vccd1 _16043_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12828_ _12822_/A _25469_/Q _25468_/Q vssd1 vssd1 vccd1 vccd1 _12975_/B sky130_fd_sc_hd__nand3b_2
X_19384_ _19448_/A _19384_/B vssd1 vssd1 vccd1 vccd1 _19384_/Y sky130_fd_sc_hd__nand2_1
XFILLER_222_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16596_ _19571_/A _19571_/B vssd1 vssd1 vccd1 vccd1 _16890_/A sky130_fd_sc_hd__nand2_1
X_18335_ _14232_/X _18285_/X _18334_/Y _18022_/X _25602_/Q vssd1 vssd1 vccd1 vccd1
+ _18336_/B sky130_fd_sc_hd__a32o_1
X_15547_ _15547_/A vssd1 vssd1 vccd1 vccd1 _16079_/S sky130_fd_sc_hd__clkbuf_4
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _26940_/Q vssd1 vssd1 vccd1 vccd1 _20487_/A sky130_fd_sc_hd__clkinv_4
XFILLER_175_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18266_ _18264_/X _18265_/X _18416_/S vssd1 vssd1 vccd1 vccd1 _18266_/X sky130_fd_sc_hd__mux2_1
X_15478_ _15538_/A _15473_/X _15477_/X _13164_/A vssd1 vssd1 vccd1 vccd1 _15478_/X
+ sky130_fd_sc_hd__o211a_1
X_17217_ _17217_/A vssd1 vssd1 vccd1 vccd1 _25497_/D sky130_fd_sc_hd__clkbuf_1
X_14429_ _13082_/A _26877_/Q _26749_/Q _14095_/A _13029_/A vssd1 vssd1 vccd1 vccd1
+ _14431_/B sky130_fd_sc_hd__a221o_1
X_18197_ _17904_/X _17955_/X _18197_/S vssd1 vssd1 vccd1 vccd1 _18197_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17148_ _17200_/A _17148_/B vssd1 vssd1 vccd1 vccd1 _17149_/A sky130_fd_sc_hd__and2_1
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17079_ _26236_/Q vssd1 vssd1 vccd1 vccd1 _17087_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20090_ _16517_/X _18016_/A _20125_/A _20125_/B vssd1 vssd1 vccd1 vccd1 _20095_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_276_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22800_ _26384_/Q _22720_/X _22800_/S vssd1 vssd1 vccd1 vccd1 _22801_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23780_ _23779_/X _26777_/Q _23780_/S vssd1 vssd1 vccd1 vccd1 _23781_/A sky130_fd_sc_hd__mux2_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20992_ _22641_/B _25249_/B vssd1 vssd1 vccd1 vccd1 _25321_/B sky130_fd_sc_hd__or2_4
XFILLER_214_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22731_ _26355_/Q _22730_/X _22737_/S vssd1 vssd1 vccd1 vccd1 _22732_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25450_ _25450_/A vssd1 vssd1 vccd1 vccd1 _25459_/S sky130_fd_sc_hd__buf_4
XFILLER_280_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22662_ _22662_/A vssd1 vssd1 vccd1 vccd1 _26333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24401_ _24392_/X _25604_/Q _24400_/X vssd1 vssd1 vccd1 vccd1 _24923_/A sky130_fd_sc_hd__o21ai_4
X_21613_ _19381_/A _21278_/A _21563_/X _21612_/X vssd1 vssd1 vccd1 vccd1 _21613_/X
+ sky130_fd_sc_hd__o211a_2
X_25381_ _27289_/Q _23770_/A _25387_/S vssd1 vssd1 vccd1 vccd1 _25382_/A sky130_fd_sc_hd__mux2_1
X_22593_ _22606_/A vssd1 vssd1 vccd1 vccd1 _22593_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_179_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24332_ _24335_/A _24334_/B vssd1 vssd1 vccd1 vccd1 _24332_/Y sky130_fd_sc_hd__nor2_1
X_27120_ _27122_/CLK _27120_/D vssd1 vssd1 vccd1 vccd1 _27120_/Q sky130_fd_sc_hd__dfxtp_4
X_21544_ _21544_/A vssd1 vssd1 vccd1 vccd1 _21544_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27051_ _27062_/CLK _27051_/D vssd1 vssd1 vccd1 vccd1 _27051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24263_ _26978_/Q _24266_/C _24209_/X vssd1 vssd1 vccd1 vccd1 _24263_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_194_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21475_ input51/X input86/X _21489_/S vssd1 vssd1 vccd1 vccd1 _21476_/A sky130_fd_sc_hd__mux2_8
XFILLER_101_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26002_ _26593_/CLK _26002_/D vssd1 vssd1 vccd1 vccd1 _26002_/Q sky130_fd_sc_hd__dfxtp_2
X_23214_ _26552_/Q _23034_/X _23222_/S vssd1 vssd1 vccd1 vccd1 _23215_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20426_ _20426_/A _20426_/B vssd1 vssd1 vccd1 vccd1 _20427_/B sky130_fd_sc_hd__xnor2_1
X_24194_ _26955_/Q _24197_/C vssd1 vssd1 vccd1 vccd1 _24195_/B sky130_fd_sc_hd__and2_1
XFILLER_101_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23145_ _23145_/A vssd1 vssd1 vccd1 vccd1 _26521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20357_ _20357_/A vssd1 vssd1 vccd1 vccd1 _20357_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23076_ _23549_/A vssd1 vssd1 vccd1 vccd1 _23076_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20288_ _19833_/X _20334_/C _20287_/Y _20100_/X vssd1 vssd1 vccd1 vccd1 _20289_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_5502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22027_ _26125_/Q _20964_/X _22027_/S vssd1 vssd1 vccd1 vccd1 _22028_/A sky130_fd_sc_hd__mux2_1
X_26904_ _26904_/CLK _26904_/D vssd1 vssd1 vccd1 vccd1 _26904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26835_ _26931_/CLK _26835_/D vssd1 vssd1 vccd1 vccd1 _26835_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13800_ _14575_/A _17818_/B vssd1 vssd1 vccd1 vccd1 _16728_/B sky130_fd_sc_hd__nor2_1
XFILLER_63_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26766_ _26827_/CLK _26766_/D vssd1 vssd1 vccd1 vccd1 _26766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14780_ _26682_/Q _25722_/Q _16510_/A vssd1 vssd1 vccd1 vccd1 _14780_/X sky130_fd_sc_hd__mux2_1
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23978_ _23989_/A vssd1 vssd1 vccd1 vccd1 _23987_/S sky130_fd_sc_hd__buf_4
XFILLER_84_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13731_ _13694_/A _25766_/Q _13719_/A _26852_/Q _13410_/X vssd1 vssd1 vccd1 vccd1
+ _13731_/X sky130_fd_sc_hd__o221a_1
XFILLER_72_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25717_ _27324_/CLK _25717_/D vssd1 vssd1 vccd1 vccd1 _25717_/Q sky130_fd_sc_hd__dfxtp_1
X_22929_ _22929_/A vssd1 vssd1 vccd1 vccd1 _26440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26697_ _26889_/CLK _26697_/D vssd1 vssd1 vccd1 vccd1 _26697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16450_ _19341_/A vssd1 vssd1 vccd1 vccd1 _16450_/Y sky130_fd_sc_hd__clkinv_2
X_25648_ _27295_/CLK _25648_/D vssd1 vssd1 vccd1 vccd1 _25648_/Q sky130_fd_sc_hd__dfxtp_1
X_13662_ _13313_/A _13646_/X _13650_/X _13661_/X vssd1 vssd1 vccd1 vccd1 _13662_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_72_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15401_ _15401_/A vssd1 vssd1 vccd1 vccd1 _16104_/A sky130_fd_sc_hd__clkbuf_8
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _25878_/Q _15820_/B vssd1 vssd1 vccd1 vccd1 _13593_/X sky130_fd_sc_hd__or2_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16381_ _15065_/X _26419_/Q _15142_/X _16380_/X vssd1 vssd1 vccd1 vccd1 _16381_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25579_ _26683_/CLK _25579_/D vssd1 vssd1 vccd1 vccd1 _25579_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18120_ _18234_/A _18120_/B _18120_/C _18120_/D vssd1 vssd1 vccd1 vccd1 _18121_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_40_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27318_ _27319_/CLK _27318_/D vssd1 vssd1 vccd1 vccd1 _27318_/Q sky130_fd_sc_hd__dfxtp_1
X_15332_ _15406_/A _26610_/Q _16189_/S _26350_/Q _16195_/S vssd1 vssd1 vccd1 vccd1
+ _15332_/X sky130_fd_sc_hd__o221a_1
XFILLER_196_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18051_ _17907_/X _17875_/X _18062_/S vssd1 vssd1 vccd1 vccd1 _18051_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27249_ _27249_/CLK _27249_/D vssd1 vssd1 vccd1 vccd1 _27249_/Q sky130_fd_sc_hd__dfxtp_1
X_15263_ _15261_/X _15262_/X _15263_/S vssd1 vssd1 vccd1 vccd1 _15263_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17002_ _16676_/A _16676_/B _20978_/B _16679_/B vssd1 vssd1 vccd1 vccd1 _17016_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14214_ _27299_/Q _26556_/Q _14289_/S vssd1 vssd1 vccd1 vccd1 _14214_/X sky130_fd_sc_hd__mux2_1
X_15194_ _25748_/Q vssd1 vssd1 vccd1 vccd1 _20687_/A sky130_fd_sc_hd__clkinv_4
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27309_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14145_ _14135_/X _14138_/Y _14141_/Y _14144_/Y _14610_/A vssd1 vssd1 vccd1 vccd1
+ _14147_/A sky130_fd_sc_hd__a311o_1
XFILLER_153_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14076_ _14076_/A _14076_/B _14076_/C vssd1 vssd1 vccd1 vccd1 _14077_/C sky130_fd_sc_hd__or3_1
X_18953_ _27021_/Q _19063_/A _18952_/X _18565_/A vssd1 vssd1 vccd1 vccd1 _18953_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_140_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13027_ _13027_/A vssd1 vssd1 vccd1 vccd1 _13028_/A sky130_fd_sc_hd__clkbuf_2
X_17904_ _17902_/X _17903_/X _17958_/S vssd1 vssd1 vccd1 vccd1 _17904_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18884_ _18891_/A vssd1 vssd1 vccd1 vccd1 _18884_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17835_ _19011_/A _19045_/B _17835_/C vssd1 vssd1 vccd1 vccd1 _17836_/C sky130_fd_sc_hd__or3_1
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17766_ _18303_/S vssd1 vssd1 vccd1 vccd1 _19140_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_212_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14978_ _16250_/A _14977_/X _14718_/X vssd1 vssd1 vccd1 vccd1 _14978_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_35_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19505_ _19499_/X _18471_/X _19504_/X _19502_/X vssd1 vssd1 vccd1 vccd1 _25636_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16717_ _16717_/A _16717_/B vssd1 vssd1 vccd1 vccd1 _18357_/A sky130_fd_sc_hd__xor2_4
X_13929_ _25916_/Q _12902_/X _15874_/A _13928_/Y vssd1 vssd1 vccd1 vccd1 _13929_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_228_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17697_ _17697_/A _17697_/B vssd1 vssd1 vccd1 vccd1 _17697_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_410 _17046_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_421 _12781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19436_ _27035_/Q _18756_/X _19435_/X _18759_/X vssd1 vssd1 vccd1 vccd1 _19436_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_432 _26236_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_443 _25731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16648_ _16657_/A _17533_/A vssd1 vssd1 vccd1 vccd1 _16648_/X sky130_fd_sc_hd__or2_1
XFILLER_35_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_454 hold1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_465 _20683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_476 _23546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19367_ _27161_/Q _19367_/B vssd1 vssd1 vccd1 vccd1 _19367_/X sky130_fd_sc_hd__or2_1
XINSDIODE2_487 _20692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_498 _19118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16579_ _17856_/A _19639_/A vssd1 vssd1 vccd1 vccd1 _16932_/B sky130_fd_sc_hd__or2_1
XFILLER_188_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18318_ _17913_/X _17880_/X _18318_/S vssd1 vssd1 vccd1 vccd1 _18318_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19298_ _25527_/Q _18807_/X _18808_/X _17427_/A vssd1 vssd1 vccd1 vccd1 _19298_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18249_ _18910_/A _18247_/X _18705_/A vssd1 vssd1 vccd1 vccd1 _18250_/C sky130_fd_sc_hd__o21ba_1
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21260_ _21407_/A _21256_/X _21258_/Y _21259_/X vssd1 vssd1 vccd1 vccd1 _21261_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20211_ _19926_/X _20209_/Y _20210_/X _24986_/B vssd1 vssd1 vccd1 vccd1 _20211_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_274_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21191_ _21195_/B _21195_/C _21195_/A vssd1 vssd1 vccd1 vccd1 _21191_/X sky130_fd_sc_hd__o21ba_1
XFILLER_116_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20142_ _20141_/B _19039_/X _19911_/X _20141_/Y vssd1 vssd1 vccd1 vccd1 _20142_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_131_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24950_ _27149_/Q _24930_/X _24948_/Y _24949_/X vssd1 vssd1 vccd1 vccd1 _27149_/D
+ sky130_fd_sc_hd__o211a_1
X_20073_ _27148_/Q _20295_/B vssd1 vssd1 vccd1 vccd1 _20073_/X sky130_fd_sc_hd__and2_1
XFILLER_258_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_257_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23901_ _23901_/A vssd1 vssd1 vccd1 vccd1 _26829_/D sky130_fd_sc_hd__clkbuf_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24881_ _27127_/Q _24890_/B vssd1 vssd1 vccd1 vccd1 _24881_/Y sky130_fd_sc_hd__nand2_1
XFILLER_245_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26620_ _26813_/CLK _26620_/D vssd1 vssd1 vccd1 vccd1 _26620_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23832_ _23747_/X _26799_/Q _23832_/S vssd1 vssd1 vccd1 vccd1 _23833_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23763_ _23763_/A vssd1 vssd1 vccd1 vccd1 _23763_/X sky130_fd_sc_hd__buf_2
X_26551_ _26939_/CLK _26551_/D vssd1 vssd1 vccd1 vccd1 _26551_/Q sky130_fd_sc_hd__dfxtp_1
X_20975_ _21562_/B vssd1 vssd1 vccd1 vccd1 _21349_/B sky130_fd_sc_hd__buf_2
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25502_ _27014_/CLK _25502_/D vssd1 vssd1 vccd1 vccd1 _25502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22714_ _23757_/A vssd1 vssd1 vccd1 vccd1 _22714_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_23694_ _23693_/X _26750_/Q _23700_/S vssd1 vssd1 vccd1 vccd1 _23695_/A sky130_fd_sc_hd__mux2_1
X_26482_ _27292_/CLK _26482_/D vssd1 vssd1 vccd1 vccd1 _26482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22645_ _26328_/Q _22640_/X _22657_/S vssd1 vssd1 vccd1 vccd1 _22646_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25433_ _23741_/X _27312_/Q _25437_/S vssd1 vssd1 vccd1 vccd1 _25434_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25364_ _25364_/A vssd1 vssd1 vccd1 vccd1 _27281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22576_ _26306_/Q _22578_/B vssd1 vssd1 vccd1 vccd1 _22576_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27103_ _27173_/CLK _27103_/D vssd1 vssd1 vccd1 vccd1 _27103_/Q sky130_fd_sc_hd__dfxtp_2
X_24315_ _26996_/Q _24318_/C _24314_/X vssd1 vssd1 vccd1 vccd1 _24315_/Y sky130_fd_sc_hd__a21oi_1
X_21527_ input56/X input91/X _21553_/S vssd1 vssd1 vccd1 vccd1 _21528_/A sky130_fd_sc_hd__mux2_8
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25295_ _25306_/A vssd1 vssd1 vccd1 vccd1 _25304_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_194_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24246_ _26972_/Q _24250_/C _24209_/X vssd1 vssd1 vccd1 vccd1 _24246_/Y sky130_fd_sc_hd__a21oi_1
X_27034_ _27164_/CLK _27034_/D vssd1 vssd1 vccd1 vccd1 _27034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21458_ _26586_/Q _21562_/B _21562_/C _21562_/D vssd1 vssd1 vccd1 vccd1 _21459_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20409_ _20396_/X _20397_/Y _19941_/X _20408_/X vssd1 vssd1 vccd1 vccd1 _20409_/Y
+ sky130_fd_sc_hd__o211ai_1
X_24177_ _26949_/Q _24178_/C _24176_/Y vssd1 vssd1 vccd1 vccd1 _26949_/D sky130_fd_sc_hd__o21a_1
XFILLER_181_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21389_ _25946_/Q _21378_/X _21388_/Y _21330_/X vssd1 vssd1 vccd1 vccd1 _25946_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23128_ _26516_/Q _23127_/X _23131_/S vssd1 vssd1 vccd1 vccd1 _23129_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23059_ _23059_/A vssd1 vssd1 vccd1 vccd1 _26494_/D sky130_fd_sc_hd__clkbuf_1
X_15950_ _17829_/A _16037_/A vssd1 vssd1 vccd1 vccd1 _16631_/A sky130_fd_sc_hd__xnor2_4
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput110 dout1[12] vssd1 vssd1 vccd1 vccd1 input110/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput121 dout1[22] vssd1 vssd1 vccd1 vccd1 input121/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput132 dout1[32] vssd1 vssd1 vccd1 vccd1 input132/X sky130_fd_sc_hd__clkbuf_2
X_14901_ _26649_/Q _26745_/Q _14981_/S vssd1 vssd1 vccd1 vccd1 _14901_/X sky130_fd_sc_hd__mux2_1
XTAP_5354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput143 dout1[42] vssd1 vssd1 vccd1 vccd1 input143/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput154 dout1[52] vssd1 vssd1 vccd1 vccd1 input154/X sky130_fd_sc_hd__clkbuf_2
XTAP_5365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15881_ _15982_/S _15879_/X _15880_/X _13998_/S vssd1 vssd1 vccd1 vccd1 _15885_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput165 dout1[62] vssd1 vssd1 vccd1 vccd1 input165/X sky130_fd_sc_hd__clkbuf_2
XTAP_5387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ _25924_/Q _17517_/X _13921_/Y _17518_/X vssd1 vssd1 vccd1 vccd1 _17620_/X
+ sky130_fd_sc_hd__a2bb2o_1
Xinput176 irq[14] vssd1 vssd1 vccd1 vccd1 _19616_/C sky130_fd_sc_hd__buf_6
XFILLER_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26818_ _27301_/CLK _26818_/D vssd1 vssd1 vccd1 vccd1 _26818_/Q sky130_fd_sc_hd__dfxtp_1
Xinput187 jtag_tck vssd1 vssd1 vccd1 vccd1 _22356_/A sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_172_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26271_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14832_ _19427_/S _14832_/B vssd1 vssd1 vccd1 vccd1 _16462_/A sky130_fd_sc_hd__nor2_4
Xinput198 localMemory_wb_adr_i[17] vssd1 vssd1 vccd1 vccd1 input198/X sky130_fd_sc_hd__clkbuf_1
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_101_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26222_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17551_ _17612_/A vssd1 vssd1 vccd1 vccd1 _17551_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_205_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26749_ _26813_/CLK _26749_/D vssd1 vssd1 vccd1 vccd1 _26749_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14763_ _14763_/A vssd1 vssd1 vccd1 vccd1 _14764_/A sky130_fd_sc_hd__buf_2
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _26095_/Q _16490_/B _16499_/S _16501_/X vssd1 vssd1 vccd1 vccd1 _16502_/X
+ sky130_fd_sc_hd__o211a_1
X_13714_ _15453_/A vssd1 vssd1 vccd1 vccd1 _16078_/S sky130_fd_sc_hd__buf_4
XFILLER_17_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17482_ _17482_/A _17482_/B vssd1 vssd1 vccd1 vccd1 _17682_/B sky130_fd_sc_hd__nor2_1
XFILLER_189_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14694_ _14694_/A vssd1 vssd1 vccd1 vccd1 _16398_/S sky130_fd_sc_hd__buf_4
XFILLER_205_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19221_ _27223_/Q _19364_/B vssd1 vssd1 vccd1 vccd1 _19221_/X sky130_fd_sc_hd__and2_1
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16433_ _26647_/Q _26743_/Q _16433_/S vssd1 vssd1 vccd1 vccd1 _16433_/X sky130_fd_sc_hd__mux2_1
X_13645_ _26073_/Q _13829_/S _13643_/X _13644_/X vssd1 vssd1 vccd1 vccd1 _13645_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19152_ _25619_/Q _18971_/X _19151_/X _19007_/X vssd1 vssd1 vccd1 vccd1 _25619_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16364_ _14802_/A _16360_/X _16363_/X _13314_/X vssd1 vssd1 vccd1 vccd1 _16364_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13576_ _12871_/A _13564_/Y _13568_/Y _13574_/X _13575_/X vssd1 vssd1 vccd1 vccd1
+ _13576_/X sky130_fd_sc_hd__o32a_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _18103_/A vssd1 vssd1 vccd1 vccd1 _18811_/A sky130_fd_sc_hd__clkbuf_2
X_15315_ _16267_/S vssd1 vssd1 vccd1 vccd1 _16443_/S sky130_fd_sc_hd__buf_4
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19083_ _18976_/X _19079_/X _19082_/X _19003_/X vssd1 vssd1 vccd1 vccd1 _19083_/X
+ sky130_fd_sc_hd__a22o_1
X_16295_ _25623_/Q _14597_/A _16294_/X _14618_/A vssd1 vssd1 vccd1 vccd1 _23590_/A
+ sky130_fd_sc_hd__o22a_4
X_18034_ _18356_/A vssd1 vssd1 vccd1 vccd1 _19290_/A sky130_fd_sc_hd__clkbuf_2
X_15246_ _15245_/X _13925_/B _14604_/A vssd1 vssd1 vccd1 vccd1 _15246_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15177_ _15171_/X _15176_/X _16398_/S vssd1 vssd1 vccd1 vccd1 _15177_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14128_ _18372_/S _14128_/B vssd1 vssd1 vccd1 vccd1 _17800_/A sky130_fd_sc_hd__or2_1
XFILLER_113_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19985_ _25672_/Q _25671_/Q _19985_/C vssd1 vssd1 vccd1 vccd1 _19985_/X sky130_fd_sc_hd__and3_1
XFILLER_113_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14059_ _13311_/A _14045_/X _14049_/X _14058_/X vssd1 vssd1 vccd1 vccd1 _14059_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_140_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18936_ _18936_/A _18936_/B _18936_/C vssd1 vssd1 vccd1 vccd1 _18936_/X sky130_fd_sc_hd__or3_1
XFILLER_268_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18867_ _27213_/Q _19299_/B vssd1 vssd1 vccd1 vccd1 _18867_/X sky130_fd_sc_hd__and2_1
XFILLER_39_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17818_ _14575_/A _17818_/B vssd1 vssd1 vccd1 vccd1 _18593_/C sky130_fd_sc_hd__and2b_2
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18798_ _18347_/X _18345_/X _18858_/S vssd1 vssd1 vccd1 vccd1 _18798_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17749_ _18116_/A _17749_/B vssd1 vssd1 vccd1 vccd1 _18111_/C sky130_fd_sc_hd__or2_1
XFILLER_282_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20760_ _20760_/A vssd1 vssd1 vccd1 vccd1 _25776_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_240 _16636_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_251 _16811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_262 _22535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19419_ _25627_/Q _18719_/A _19418_/X _19352_/X vssd1 vssd1 vccd1 vccd1 _25627_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_251_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_273 INSDIODE2_273/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20691_ _26286_/Q _20686_/X _20690_/Y _20684_/X vssd1 vssd1 vccd1 vccd1 _25749_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_284 _25816_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_295 _25826_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22430_ _26245_/Q _22430_/B vssd1 vssd1 vccd1 vccd1 _22430_/X sky130_fd_sc_hd__or2_1
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22361_ _22361_/A _22361_/B vssd1 vssd1 vccd1 vccd1 _22362_/B sky130_fd_sc_hd__or2_1
XFILLER_248_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24100_ _24146_/S vssd1 vssd1 vccd1 vccd1 _24109_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_136_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21312_ _21284_/X _18404_/X _21286_/X _25802_/Q _21641_/B vssd1 vssd1 vccd1 vccd1
+ _21312_/X sky130_fd_sc_hd__a221o_1
XFILLER_175_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25080_ _22500_/A _25065_/X _25060_/X _16636_/C _25079_/X vssd1 vssd1 vccd1 vccd1
+ _25080_/X sky130_fd_sc_hd__a221o_1
X_22292_ _26209_/Q _22279_/X _22285_/X _26310_/Q _22286_/X vssd1 vssd1 vccd1 vccd1
+ _22292_/X sky130_fd_sc_hd__a221o_1
XFILLER_191_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24031_ _26887_/Q _23546_/X _24037_/S vssd1 vssd1 vccd1 vccd1 _24032_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21243_ _25936_/Q _21202_/X _21240_/Y _21242_/X vssd1 vssd1 vccd1 vccd1 _25936_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_117_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21174_ _21174_/A vssd1 vssd1 vccd1 vccd1 _21188_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20125_ _20125_/A _20125_/B _20125_/C _20125_/D vssd1 vssd1 vccd1 vccd1 _20126_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_259_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25982_ _25985_/CLK _25982_/D vssd1 vssd1 vccd1 vccd1 _25982_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_58_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24933_ _19896_/A _24930_/X _24932_/Y _24921_/X vssd1 vssd1 vccd1 vccd1 _27142_/D
+ sky130_fd_sc_hd__o211a_1
X_20056_ _19824_/B _18894_/X _19663_/X _20055_/X vssd1 vssd1 vccd1 vccd1 _20056_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24864_ _20679_/A _24848_/X _24732_/Y _24849_/X vssd1 vssd1 vccd1 vccd1 _24864_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_73_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26603_ _27278_/CLK _26603_/D vssd1 vssd1 vccd1 vccd1 _26603_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23815_ _23722_/X _26791_/Q _23821_/S vssd1 vssd1 vccd1 vccd1 _23816_/A sky130_fd_sc_hd__mux2_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24795_ _20630_/A _24789_/X _24654_/A _24791_/X vssd1 vssd1 vccd1 vccd1 _24795_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26534_ _27309_/CLK _26534_/D vssd1 vssd1 vccd1 vccd1 _26534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23746_ _23746_/A vssd1 vssd1 vccd1 vccd1 _26766_/D sky130_fd_sc_hd__clkbuf_1
X_20958_ _23773_/A vssd1 vssd1 vccd1 vccd1 _20958_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26465_ _26465_/CLK _26465_/D vssd1 vssd1 vccd1 vccd1 _26465_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20889_ _25834_/Q _20887_/X _20901_/S vssd1 vssd1 vccd1 vccd1 _20890_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23677_ _23677_/A vssd1 vssd1 vccd1 vccd1 _26744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13430_ _26498_/Q _26370_/Q _15800_/S vssd1 vssd1 vccd1 vccd1 _13430_/X sky130_fd_sc_hd__mux2_1
X_25416_ _25416_/A vssd1 vssd1 vccd1 vccd1 _27304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22628_ _22638_/A _22554_/A _22624_/X _22638_/C vssd1 vssd1 vccd1 vccd1 _22631_/A
+ sky130_fd_sc_hd__o31a_1
X_26396_ _27267_/CLK _26396_/D vssd1 vssd1 vccd1 vccd1 _26396_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13361_ _16022_/A vssd1 vssd1 vccd1 vccd1 _15776_/A sky130_fd_sc_hd__buf_2
XFILLER_139_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25347_ _25347_/A vssd1 vssd1 vccd1 vccd1 _27273_/D sky130_fd_sc_hd__clkbuf_1
X_22559_ _22553_/X _22558_/Y _22547_/X vssd1 vssd1 vccd1 vccd1 _26299_/D sky130_fd_sc_hd__a21oi_1
XFILLER_6_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15100_ _14744_/A _25784_/Q _15221_/S _26870_/Q _15120_/S vssd1 vssd1 vccd1 vccd1
+ _15100_/X sky130_fd_sc_hd__o221a_1
X_13292_ _15394_/A _13283_/X _13290_/X _13291_/X vssd1 vssd1 vccd1 vccd1 _13292_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16080_ _16074_/X _16076_/X _16079_/X _15647_/S _12703_/A vssd1 vssd1 vccd1 vccd1
+ _16080_/X sky130_fd_sc_hd__o221a_1
X_25278_ _23725_/X _27243_/Q _25282_/S vssd1 vssd1 vccd1 vccd1 _25279_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27017_ _27049_/CLK _27017_/D vssd1 vssd1 vccd1 vccd1 _27017_/Q sky130_fd_sc_hd__dfxtp_1
X_15031_ _15031_/A vssd1 vssd1 vccd1 vccd1 _16308_/S sky130_fd_sc_hd__clkbuf_4
X_24229_ _26966_/Q _24225_/B _24228_/Y vssd1 vssd1 vccd1 vccd1 _26966_/D sky130_fd_sc_hd__o21a_1
XFILLER_108_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19770_ _19824_/B _19768_/Y _19663_/X _19769_/X vssd1 vssd1 vccd1 vccd1 _19770_/X
+ sky130_fd_sc_hd__o31a_1
X_16982_ _17856_/A _16982_/B _16982_/C vssd1 vssd1 vccd1 vccd1 _16982_/X sky130_fd_sc_hd__and3b_1
XFILLER_123_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18721_ _18721_/A vssd1 vssd1 vccd1 vccd1 _19252_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15933_ _13330_/A _15930_/X _15932_/X _13340_/A vssd1 vssd1 vccd1 vccd1 _15933_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18652_ _17268_/X _18439_/X _18441_/X _25543_/Q vssd1 vssd1 vccd1 vccd1 _18652_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _15860_/X _15863_/X _13530_/X vssd1 vssd1 vccd1 vccd1 _15864_/Y sky130_fd_sc_hd__o21ai_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ _17615_/A _17603_/B vssd1 vssd1 vccd1 vccd1 _25582_/D sky130_fd_sc_hd__nor2_1
XFILLER_224_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14815_ _14755_/X _14813_/X _14814_/X _14794_/X vssd1 vssd1 vccd1 vccd1 _14815_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18583_ _18579_/X _18581_/X _18582_/X _18377_/A _18005_/A vssd1 vssd1 vccd1 vccd1
+ _18583_/X sky130_fd_sc_hd__a221o_1
XFILLER_252_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15795_ _25612_/Q _14595_/A _15794_/X _14616_/A vssd1 vssd1 vccd1 vccd1 _15833_/A
+ sky130_fd_sc_hd__o22a_4
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ _17653_/A vssd1 vssd1 vccd1 vccd1 _17534_/X sky130_fd_sc_hd__buf_2
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14746_ _14746_/A vssd1 vssd1 vccd1 vccd1 _14747_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_251_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17465_ _17465_/A _17708_/B vssd1 vssd1 vccd1 vccd1 _17471_/A sky130_fd_sc_hd__or2_1
X_14677_ _14677_/A vssd1 vssd1 vccd1 vccd1 _14678_/A sky130_fd_sc_hd__clkbuf_4
X_19204_ _26964_/Q _18569_/X _18570_/X _26996_/Q vssd1 vssd1 vccd1 vccd1 _19204_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16416_ _19828_/A _16284_/S _16415_/Y vssd1 vssd1 vccd1 vccd1 _17780_/A sky130_fd_sc_hd__o21ai_2
X_13628_ _12769_/A _26693_/Q _26821_/Q _15961_/B _13049_/A vssd1 vssd1 vccd1 vccd1
+ _13628_/X sky130_fd_sc_hd__a221o_1
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17396_ _17395_/X _17399_/C _17366_/X vssd1 vssd1 vccd1 vccd1 _17396_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19135_ _27058_/Q _19055_/X _19132_/X _19134_/X _19066_/X vssd1 vssd1 vccd1 vccd1
+ _19135_/X sky130_fd_sc_hd__o221a_2
XFILLER_34_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16347_ _25854_/Q _26054_/Q _16347_/S vssd1 vssd1 vccd1 vccd1 _16347_/X sky130_fd_sc_hd__mux2_1
X_13559_ _14025_/B _13559_/B vssd1 vssd1 vccd1 vccd1 _15708_/B sky130_fd_sc_hd__nor2_1
XFILLER_185_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19066_ _19066_/A vssd1 vssd1 vccd1 vccd1 _19066_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16278_ _16276_/X _16277_/X _16278_/S vssd1 vssd1 vccd1 vccd1 _16278_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18017_ _19087_/A vssd1 vssd1 vccd1 vccd1 _18976_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput403 _17011_/X vssd1 vssd1 vccd1 vccd1 din0[5] sky130_fd_sc_hd__buf_2
X_15229_ _15308_/S vssd1 vssd1 vccd1 vccd1 _16360_/S sky130_fd_sc_hd__clkbuf_4
Xoutput414 _25949_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[13] sky130_fd_sc_hd__buf_2
Xoutput425 _25959_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[23] sky130_fd_sc_hd__buf_2
Xoutput436 _25940_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[4] sky130_fd_sc_hd__buf_2
Xoutput447 _26234_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[2] sky130_fd_sc_hd__buf_2
XFILLER_5_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput458 _25741_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[17] sky130_fd_sc_hd__buf_2
Xoutput469 _25751_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[27] sky130_fd_sc_hd__buf_2
XFILLER_259_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19968_ _19968_/A vssd1 vssd1 vccd1 vccd1 _20089_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18919_ _27052_/Q _19055_/A _18916_/X _18918_/X _19066_/A vssd1 vssd1 vccd1 vccd1
+ _18919_/X sky130_fd_sc_hd__o221a_1
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19899_ _19895_/X _19896_/Y _19898_/Y vssd1 vssd1 vccd1 vccd1 _19899_/Y sky130_fd_sc_hd__a21oi_1
X_21930_ _21930_/A vssd1 vssd1 vccd1 vccd1 _26081_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_283_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21861_ _21861_/A vssd1 vssd1 vccd1 vccd1 _26058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_271_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20812_ _25802_/Q vssd1 vssd1 vccd1 vccd1 _20813_/A sky130_fd_sc_hd__clkbuf_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23600_ _23600_/A vssd1 vssd1 vccd1 vccd1 _23600_/X sky130_fd_sc_hd__clkbuf_2
X_24580_ _24619_/A vssd1 vssd1 vccd1 vccd1 _24580_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_21792_ _21792_/A vssd1 vssd1 vccd1 vccd1 _26028_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20743_ _20743_/A vssd1 vssd1 vccd1 vccd1 _25768_/D sky130_fd_sc_hd__clkbuf_1
X_23531_ _26690_/Q _23530_/X _23540_/S vssd1 vssd1 vccd1 vccd1 _23532_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23462_ _23462_/A vssd1 vssd1 vccd1 vccd1 _26662_/D sky130_fd_sc_hd__clkbuf_1
X_26250_ _26250_/CLK _26250_/D vssd1 vssd1 vccd1 vccd1 _26250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20674_ _20674_/A vssd1 vssd1 vccd1 vccd1 _20683_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_51_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22413_ _22361_/A _22379_/X _22405_/B _22412_/Y _22402_/X vssd1 vssd1 vccd1 vccd1
+ _26240_/D sky130_fd_sc_hd__o221a_1
X_25201_ _24693_/B _25198_/X _25196_/X _27211_/Q _25199_/X vssd1 vssd1 vccd1 vccd1
+ _27211_/D sky130_fd_sc_hd__o221a_1
X_26181_ _26319_/CLK _26181_/D vssd1 vssd1 vccd1 vccd1 _26181_/Q sky130_fd_sc_hd__dfxtp_1
X_23393_ _26632_/Q _23076_/X _23397_/S vssd1 vssd1 vccd1 vccd1 _23394_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22344_ _22337_/X _17078_/X _26227_/Q vssd1 vssd1 vccd1 vccd1 _22344_/X sky130_fd_sc_hd__a21o_1
XFILLER_163_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25132_ _27190_/Q _25112_/X _25131_/X vssd1 vssd1 vccd1 vccd1 _27190_/D sky130_fd_sc_hd__o21ba_1
XFILLER_275_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25063_ _24686_/Y _25043_/X _25062_/Y _25055_/X vssd1 vssd1 vccd1 vccd1 _25063_/X
+ sky130_fd_sc_hd__a31o_1
X_22275_ _26203_/Q _22264_/X _22270_/X _26304_/Q _22271_/X vssd1 vssd1 vccd1 vccd1
+ _22275_/X sky130_fd_sc_hd__a221o_1
X_24014_ _24014_/A vssd1 vssd1 vccd1 vccd1 _26879_/D sky130_fd_sc_hd__clkbuf_1
X_21226_ _21603_/A vssd1 vssd1 vccd1 vccd1 _21407_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21157_ _25924_/Q _21148_/X _21149_/X input24/X vssd1 vssd1 vccd1 vccd1 _21158_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_132_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20108_ _27149_/Q _20219_/B vssd1 vssd1 vccd1 vccd1 _20108_/Y sky130_fd_sc_hd__nand2_1
XFILLER_259_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25965_ _26995_/CLK _25965_/D vssd1 vssd1 vccd1 vccd1 _25965_/Q sky130_fd_sc_hd__dfxtp_1
X_21088_ _25905_/Q _21074_/X _21077_/X input35/X vssd1 vssd1 vccd1 vccd1 _21089_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_59_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12930_ _15245_/A _12926_/X _12929_/X vssd1 vssd1 vccd1 vccd1 _12930_/X sky130_fd_sc_hd__a21o_1
X_24916_ _27136_/Q _24913_/X _24915_/Y _24631_/X vssd1 vssd1 vccd1 vccd1 _27136_/D
+ sky130_fd_sc_hd__o211a_1
X_20039_ _20039_/A _20039_/B vssd1 vssd1 vccd1 vccd1 _20039_/X sky130_fd_sc_hd__and2_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25896_ _26900_/CLK _25896_/D vssd1 vssd1 vccd1 vccd1 _25896_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _12835_/Y _15704_/A _12849_/X _12857_/X _12933_/B vssd1 vssd1 vccd1 vccd1
+ _12911_/A sky130_fd_sc_hd__a2111oi_4
X_24847_ _27118_/Q _24856_/B vssd1 vssd1 vccd1 vccd1 _24847_/Y sky130_fd_sc_hd__nand2_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14600_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14601_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _16261_/S _15578_/X _15579_/X _13274_/A vssd1 vssd1 vccd1 vccd1 _15581_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24778_ _24801_/A vssd1 vssd1 vccd1 vccd1 _24779_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _25579_/Q _17218_/A _17978_/A vssd1 vssd1 vccd1 vccd1 _17971_/C sky130_fd_sc_hd__o21bai_2
XFILLER_233_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _13344_/A _14529_/X _14530_/X _13309_/B vssd1 vssd1 vccd1 vccd1 _14535_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_214_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26517_ _27321_/CLK _26517_/D vssd1 vssd1 vccd1 vccd1 _26517_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23729_ _23728_/X _26761_/Q _23732_/S vssd1 vssd1 vccd1 vccd1 _23730_/A sky130_fd_sc_hd__mux2_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _18338_/A vssd1 vssd1 vccd1 vccd1 _20973_/A sky130_fd_sc_hd__clkbuf_8
X_14462_ _13955_/A _14458_/X _14461_/X _13210_/A vssd1 vssd1 vccd1 vccd1 _14462_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26448_ _27287_/CLK _26448_/D vssd1 vssd1 vccd1 vccd1 _26448_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16201_ _16185_/X _16200_/X _14722_/A vssd1 vssd1 vccd1 vccd1 _16201_/Y sky130_fd_sc_hd__a21oi_2
X_13413_ _26918_/Q _15471_/S vssd1 vssd1 vccd1 vccd1 _13413_/X sky130_fd_sc_hd__or2_1
X_17181_ _17181_/A _17195_/B vssd1 vssd1 vccd1 vccd1 _17181_/Y sky130_fd_sc_hd__nand2_1
X_14393_ _14064_/X _14391_/X _14392_/X _14067_/X vssd1 vssd1 vccd1 vccd1 _14393_/X
+ sky130_fd_sc_hd__o211a_1
X_26379_ _26796_/CLK _26379_/D vssd1 vssd1 vccd1 vccd1 _26379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16132_ _25619_/Q _14596_/A _16131_/X _14617_/A vssd1 vssd1 vccd1 vccd1 _23578_/A
+ sky130_fd_sc_hd__o22a_4
X_13344_ _13344_/A vssd1 vssd1 vccd1 vccd1 _13512_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_183_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16063_ _14870_/A _16060_/X _16062_/X _15039_/A vssd1 vssd1 vccd1 vccd1 _16063_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_155_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13275_ _16348_/S _13264_/X _13268_/X _13274_/X vssd1 vssd1 vccd1 vccd1 _13276_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_154_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15014_ _27321_/Q _26578_/Q _15014_/S vssd1 vssd1 vccd1 vccd1 _15014_/X sky130_fd_sc_hd__mux2_1
XFILLER_269_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19822_ _22483_/A _19721_/X _19813_/X _19821_/X _19758_/X vssd1 vssd1 vccd1 vccd1
+ _25666_/D sky130_fd_sc_hd__o221a_1
XFILLER_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16965_ _16980_/A _16965_/B _16965_/C vssd1 vssd1 vccd1 vccd1 _16966_/A sky130_fd_sc_hd__and3_2
X_19753_ _19753_/A _19753_/B vssd1 vssd1 vccd1 vccd1 _19753_/Y sky130_fd_sc_hd__xnor2_1
X_15916_ _15916_/A _15916_/B vssd1 vssd1 vccd1 vccd1 _15916_/X sky130_fd_sc_hd__or2_1
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18704_ _18435_/X _18702_/X _18703_/Y vssd1 vssd1 vccd1 vccd1 _18704_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_237_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19684_ _27136_/Q _27070_/Q vssd1 vssd1 vccd1 vccd1 _19686_/B sky130_fd_sc_hd__xor2_1
XFILLER_237_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16896_ _16896_/A _16932_/B vssd1 vssd1 vccd1 vccd1 _16896_/X sky130_fd_sc_hd__or2_1
XFILLER_253_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18635_ _18635_/A _18635_/B vssd1 vssd1 vccd1 vccd1 _19574_/A sky130_fd_sc_hd__and2_1
X_15847_ _14727_/A _15845_/X _15846_/X _13367_/A vssd1 vssd1 vccd1 vccd1 _15847_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_209_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18566_ _27013_/Q _18514_/X _18564_/X _18565_/X vssd1 vssd1 vccd1 vccd1 _18566_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15778_ _13488_/A _26923_/Q _26407_/Q _15485_/S _16015_/A vssd1 vssd1 vccd1 vccd1
+ _15778_/X sky130_fd_sc_hd__a221o_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17517_ _17597_/A vssd1 vssd1 vccd1 vccd1 _17517_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14729_ _14729_/A vssd1 vssd1 vccd1 vccd1 _15227_/S sky130_fd_sc_hd__clkbuf_4
X_18497_ _18547_/S _18496_/Y _17988_/A vssd1 vssd1 vccd1 vccd1 _18497_/X sky130_fd_sc_hd__a21bo_2
XFILLER_232_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17448_ _26325_/Q vssd1 vssd1 vccd1 vccd1 _22633_/A sky130_fd_sc_hd__clkinv_2
XFILLER_177_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ _25544_/Q _25545_/Q _17379_/C vssd1 vssd1 vccd1 vccd1 _17381_/B sky130_fd_sc_hd__and3_1
XFILLER_118_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27315_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19118_ _19252_/A _19118_/B vssd1 vssd1 vccd1 vccd1 _19118_/X sky130_fd_sc_hd__or2_1
X_20390_ _20370_/A _20367_/Y _20369_/B vssd1 vssd1 vccd1 vccd1 _20391_/B sky130_fd_sc_hd__o21ai_1
XFILLER_174_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19049_ _19049_/A _19579_/B vssd1 vssd1 vccd1 vccd1 _19049_/X sky130_fd_sc_hd__or2_1
XFILLER_134_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22060_ _26139_/Q _20907_/X _22066_/S vssd1 vssd1 vccd1 vccd1 _22061_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21011_ _25876_/Q _20894_/X _21015_/S vssd1 vssd1 vccd1 vccd1 _21012_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput288 _17066_/X vssd1 vssd1 vccd1 vccd1 addr0[3] sky130_fd_sc_hd__buf_2
Xoutput299 _16997_/X vssd1 vssd1 vccd1 vccd1 addr1[5] sky130_fd_sc_hd__buf_2
XFILLER_141_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_6 _22368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25750_ _26292_/CLK _25750_/D vssd1 vssd1 vccd1 vccd1 _25750_/Q sky130_fd_sc_hd__dfxtp_4
X_22962_ _22962_/A _25321_/B vssd1 vssd1 vccd1 vccd1 _23019_/A sky130_fd_sc_hd__nor2_8
XFILLER_256_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24701_ _24701_/A vssd1 vssd1 vccd1 vccd1 _24701_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_283_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21913_ _21959_/S vssd1 vssd1 vccd1 vccd1 _21922_/S sky130_fd_sc_hd__buf_2
XFILLER_243_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25681_ _25690_/CLK _25681_/D vssd1 vssd1 vccd1 vccd1 _25681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22893_ _26424_/Q _22640_/X _22901_/S vssd1 vssd1 vccd1 vccd1 _22894_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24632_ _27068_/Q _24553_/B _24629_/Y _24631_/X vssd1 vssd1 vccd1 vccd1 _27068_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21844_ _21844_/A vssd1 vssd1 vccd1 vccd1 _26050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24563_ _24920_/A _24569_/B vssd1 vssd1 vccd1 vccd1 _24563_/Y sky130_fd_sc_hd__nand2_1
X_21775_ _21775_/A vssd1 vssd1 vccd1 vccd1 _26020_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26302_ _26327_/CLK _26302_/D vssd1 vssd1 vccd1 vccd1 _26302_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_169_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20726_ _20504_/X _25761_/Q _20728_/S vssd1 vssd1 vccd1 vccd1 _20727_/A sky130_fd_sc_hd__mux2_1
X_23514_ _23514_/A vssd1 vssd1 vccd1 vccd1 _23514_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27282_ _27282_/CLK _27282_/D vssd1 vssd1 vccd1 vccd1 _27282_/Q sky130_fd_sc_hd__dfxtp_1
X_24494_ _24494_/A vssd1 vssd1 vccd1 vccd1 _24518_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_211_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26233_ _27297_/CLK _26233_/D vssd1 vssd1 vccd1 vccd1 _26233_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_211_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23445_ _26655_/Q _23047_/X _23447_/S vssd1 vssd1 vccd1 vccd1 _23446_/A sky130_fd_sc_hd__mux2_1
X_20657_ _20657_/A vssd1 vssd1 vccd1 vccd1 _21878_/A sky130_fd_sc_hd__buf_8
XFILLER_139_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26164_ _27264_/CLK _26164_/D vssd1 vssd1 vccd1 vccd1 _26164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23376_ _23376_/A vssd1 vssd1 vccd1 vccd1 _26624_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20588_ _23760_/A vssd1 vssd1 vccd1 vccd1 _20588_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25115_ _22513_/A _25092_/X _25114_/X _19118_/B _25106_/X vssd1 vssd1 vccd1 vccd1
+ _25115_/X sky130_fd_sc_hd__a221o_1
X_22327_ _26221_/Q _22154_/A _22316_/X _26322_/Q _22317_/X vssd1 vssd1 vccd1 vccd1
+ _22327_/X sky130_fd_sc_hd__a221o_1
XFILLER_165_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26095_ _27326_/CLK _26095_/D vssd1 vssd1 vccd1 vccd1 _26095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13060_ _15474_/S vssd1 vssd1 vccd1 vccd1 _15557_/S sky130_fd_sc_hd__buf_2
X_22258_ _22288_/A vssd1 vssd1 vccd1 vccd1 _22258_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_180_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25046_ _24671_/Y _25043_/X _25045_/Y _25027_/X vssd1 vssd1 vccd1 vccd1 _25046_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_140_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21209_ _21214_/A _21209_/B _21212_/B _21218_/D vssd1 vssd1 vccd1 vccd1 _21210_/B
+ sky130_fd_sc_hd__or4b_1
X_22189_ _26180_/Q _22185_/X _22188_/X _22181_/X vssd1 vssd1 vccd1 vccd1 _26180_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_239_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26997_ _27001_/CLK _26997_/D vssd1 vssd1 vccd1 vccd1 _26997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16750_ _25676_/Q vssd1 vssd1 vccd1 vccd1 _22505_/A sky130_fd_sc_hd__buf_2
X_13962_ _25803_/Q _27237_/Q _14310_/S vssd1 vssd1 vccd1 vccd1 _13962_/X sky130_fd_sc_hd__mux2_1
X_25948_ _25985_/CLK _25948_/D vssd1 vssd1 vccd1 vccd1 _25948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15701_ _17837_/A _15701_/B vssd1 vssd1 vccd1 vccd1 _15702_/A sky130_fd_sc_hd__nor2_1
XFILLER_247_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_79_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27298_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12913_ _12913_/A vssd1 vssd1 vccd1 vccd1 _15245_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_219_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16681_ _16660_/A _17020_/A _17060_/A _25980_/Q vssd1 vssd1 vccd1 vccd1 _16681_/Y
+ sky130_fd_sc_hd__a22oi_4
X_25879_ _27277_/CLK _25879_/D vssd1 vssd1 vccd1 vccd1 _25879_/Q sky130_fd_sc_hd__dfxtp_1
X_13893_ _14257_/A vssd1 vssd1 vccd1 vccd1 _15980_/S sky130_fd_sc_hd__buf_6
XFILLER_235_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18420_ _18898_/A _18415_/X _18419_/X vssd1 vssd1 vccd1 vccd1 _18421_/B sky130_fd_sc_hd__o21ai_1
XFILLER_206_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15632_ _26504_/Q _26376_/Q _15643_/S vssd1 vssd1 vccd1 vccd1 _15632_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _25861_/Q _25790_/Q vssd1 vssd1 vccd1 vccd1 _14403_/A sky130_fd_sc_hd__nand2_4
XFILLER_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _18547_/S _18346_/X _18350_/X vssd1 vssd1 vccd1 vccd1 _18352_/B sky130_fd_sc_hd__o21ai_2
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _13086_/X _26893_/Q _26765_/Q _15653_/S vssd1 vssd1 vccd1 vccd1 _15563_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _12775_/A vssd1 vssd1 vccd1 vccd1 _12776_/A sky130_fd_sc_hd__buf_2
XFILLER_202_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17299_/X _17303_/C _25521_/Q vssd1 vssd1 vccd1 vccd1 _17304_/B sky130_fd_sc_hd__a21oi_1
XFILLER_187_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14514_ _26520_/Q _26128_/Q _14514_/S vssd1 vssd1 vccd1 vccd1 _14514_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ _14317_/X _18013_/X _18281_/Y _18022_/X _25601_/Q vssd1 vssd1 vccd1 vccd1
+ _18283_/B sky130_fd_sc_hd__a32o_1
X_15494_ _16183_/S _15489_/X _15493_/X _14228_/X vssd1 vssd1 vccd1 vccd1 _15495_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17233_ _25176_/A vssd1 vssd1 vccd1 vccd1 _24208_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_174_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14445_ _25573_/Q _14443_/A _14193_/B vssd1 vssd1 vccd1 vccd1 _14445_/X sky130_fd_sc_hd__o21a_1
X_17164_ _19455_/B _20689_/A vssd1 vssd1 vccd1 vccd1 _17164_/X sky130_fd_sc_hd__or2_2
X_14376_ _12736_/A _25760_/Q _14539_/S _26846_/Q _14473_/S vssd1 vssd1 vccd1 vccd1
+ _14376_/X sky130_fd_sc_hd__o221a_1
XFILLER_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16115_ _13255_/A _26863_/Q _25777_/Q _16260_/S _13335_/A vssd1 vssd1 vccd1 vccd1
+ _16115_/X sky130_fd_sc_hd__a221o_1
X_13327_ _16342_/S _13325_/X _13326_/X _13274_/X vssd1 vssd1 vccd1 vccd1 _13327_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17095_ _26238_/Q _26237_/Q vssd1 vssd1 vccd1 vccd1 _22387_/B sky130_fd_sc_hd__or2_1
XFILLER_142_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16046_ _25649_/Q _16130_/B vssd1 vssd1 vccd1 vccd1 _16046_/X sky130_fd_sc_hd__and2_1
X_13258_ _14551_/S vssd1 vssd1 vccd1 vccd1 _14308_/S sky130_fd_sc_hd__buf_2
XFILLER_282_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13189_ _14459_/S vssd1 vssd1 vccd1 vccd1 _14452_/S sky130_fd_sc_hd__buf_4
XFILLER_111_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19805_ _19805_/A _19805_/B vssd1 vssd1 vccd1 vccd1 _19805_/X sky130_fd_sc_hd__or2_1
XFILLER_215_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17997_ _17997_/A vssd1 vssd1 vccd1 vccd1 _19393_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_215_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19736_ _19853_/A _19736_/B vssd1 vssd1 vccd1 vccd1 _19777_/B sky130_fd_sc_hd__nor2_1
X_16948_ _16948_/A _16948_/B vssd1 vssd1 vccd1 vccd1 _16949_/B sky130_fd_sc_hd__nor2_4
XFILLER_284_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19667_ _19943_/B _19670_/A vssd1 vssd1 vccd1 vccd1 _19727_/A sky130_fd_sc_hd__nor2_1
X_16879_ _16855_/A _16877_/X _16878_/X _16842_/A vssd1 vssd1 vccd1 vccd1 _16880_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18618_ _27046_/Q _18503_/A _18613_/X _18617_/X _18519_/A vssd1 vssd1 vccd1 vccd1
+ _18618_/X sky130_fd_sc_hd__o221a_1
XFILLER_252_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19598_ _19769_/B vssd1 vssd1 vccd1 vccd1 _20227_/B sky130_fd_sc_hd__buf_2
XFILLER_252_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18549_ _18368_/X _18371_/X _18549_/S vssd1 vssd1 vccd1 vccd1 _18549_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21560_ _21284_/A _19230_/X _21286_/A _25821_/Q _21547_/A vssd1 vssd1 vccd1 vccd1
+ _21560_/X sky130_fd_sc_hd__a221o_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20511_ _23526_/A vssd1 vssd1 vccd1 vccd1 _23702_/A sky130_fd_sc_hd__buf_4
XFILLER_166_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21491_ _21488_/X _21462_/X _21490_/Y _21451_/X vssd1 vssd1 vccd1 vccd1 _21491_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_193_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23230_ _23230_/A vssd1 vssd1 vccd1 vccd1 _26559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20442_ _22533_/A _20467_/C vssd1 vssd1 vccd1 vccd1 _20442_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_118_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23161_ _26529_/Q _23066_/X _23161_/S vssd1 vssd1 vccd1 vccd1 _23162_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20373_ _22526_/A _20003_/X _20365_/X _20372_/X _20346_/X vssd1 vssd1 vccd1 vccd1
+ _25686_/D sky130_fd_sc_hd__o221a_1
XFILLER_256_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22112_ _22170_/A vssd1 vssd1 vccd1 vccd1 _22310_/A sky130_fd_sc_hd__buf_2
XFILLER_161_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23092_ _23565_/A vssd1 vssd1 vccd1 vccd1 _23092_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22043_ _22043_/A vssd1 vssd1 vccd1 vccd1 _26131_/D sky130_fd_sc_hd__clkbuf_1
X_26920_ _26920_/CLK _26920_/D vssd1 vssd1 vccd1 vccd1 _26920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26851_ _26917_/CLK _26851_/D vssd1 vssd1 vccd1 vccd1 _26851_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_87_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25802_ _26520_/CLK _25802_/D vssd1 vssd1 vccd1 vccd1 _25802_/Q sky130_fd_sc_hd__dfxtp_4
X_26782_ _27295_/CLK _26782_/D vssd1 vssd1 vccd1 vccd1 _26782_/Q sky130_fd_sc_hd__dfxtp_1
X_23994_ _26871_/Q _23597_/X _23998_/S vssd1 vssd1 vccd1 vccd1 _23995_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25733_ _26271_/CLK _25733_/D vssd1 vssd1 vccd1 vccd1 _25733_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_228_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22945_ _26448_/Q _22720_/X _22945_/S vssd1 vssd1 vccd1 vccd1 _22946_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25664_ _25670_/CLK _25664_/D vssd1 vssd1 vccd1 vccd1 _25664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22876_ _26417_/Q _22723_/X _22884_/S vssd1 vssd1 vccd1 vccd1 _22877_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24615_ _24615_/A vssd1 vssd1 vccd1 vccd1 _24615_/X sky130_fd_sc_hd__clkbuf_2
X_21827_ _26043_/Q _20916_/X _21827_/S vssd1 vssd1 vccd1 vccd1 _21828_/A sky130_fd_sc_hd__mux2_1
XPHY_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25595_ _25596_/CLK _25595_/D vssd1 vssd1 vccd1 vccd1 _25595_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24546_ _24629_/B vssd1 vssd1 vccd1 vccd1 _24546_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21758_ _21758_/A vssd1 vssd1 vccd1 vccd1 _26012_/D sky130_fd_sc_hd__clkbuf_1
XPHY_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27265_ _27265_/CLK _27265_/D vssd1 vssd1 vccd1 vccd1 _27265_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_197_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26900_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20709_ _25757_/Q _20712_/B vssd1 vssd1 vccd1 vccd1 _20709_/Y sky130_fd_sc_hd__nand2_1
X_24477_ _24725_/B vssd1 vssd1 vccd1 vccd1 _24600_/A sky130_fd_sc_hd__clkinv_2
X_21689_ _21689_/A vssd1 vssd1 vccd1 vccd1 _25983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26216_ _26319_/CLK _26216_/D vssd1 vssd1 vccd1 vccd1 _26216_/Q sky130_fd_sc_hd__dfxtp_1
X_14230_ _13367_/X _14204_/X _14211_/X _13509_/A _14229_/X vssd1 vssd1 vccd1 vccd1
+ _14230_/X sky130_fd_sc_hd__a311o_2
Xclkbuf_leaf_126_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25518_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23428_ _26648_/Q _23127_/X _23430_/S vssd1 vssd1 vccd1 vccd1 _23429_/A sky130_fd_sc_hd__mux2_1
X_27196_ _27196_/CLK _27196_/D vssd1 vssd1 vccd1 vccd1 _27196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14161_ _14159_/X _14160_/X _15903_/S vssd1 vssd1 vccd1 vccd1 _14161_/X sky130_fd_sc_hd__mux2_1
X_26147_ _26673_/CLK _26147_/D vssd1 vssd1 vccd1 vccd1 _26147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23359_ _20617_/X _26618_/Q _23361_/S vssd1 vssd1 vccd1 vccd1 _23360_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13112_ _13112_/A vssd1 vssd1 vccd1 vccd1 _14713_/A sky130_fd_sc_hd__buf_2
XFILLER_152_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26078_ _27277_/CLK _26078_/D vssd1 vssd1 vccd1 vccd1 _26078_/Q sky130_fd_sc_hd__dfxtp_2
X_14092_ _14090_/X _14091_/X _14115_/S vssd1 vssd1 vccd1 vccd1 _14093_/B sky130_fd_sc_hd__mux2_1
XFILLER_113_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13043_ _13043_/A vssd1 vssd1 vccd1 vccd1 _15459_/S sky130_fd_sc_hd__buf_2
X_17920_ _18729_/A vssd1 vssd1 vccd1 vccd1 _17920_/X sky130_fd_sc_hd__clkbuf_2
X_25029_ _27171_/Q _25000_/X _25028_/X vssd1 vssd1 vccd1 vccd1 _27171_/D sky130_fd_sc_hd__o21ba_1
XFILLER_79_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17851_ _17851_/A _17851_/B vssd1 vssd1 vccd1 vccd1 _19389_/C sky130_fd_sc_hd__nand2_1
XFILLER_67_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16802_ _16906_/A vssd1 vssd1 vccd1 vccd1 _16910_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17782_ _17782_/A _17782_/B vssd1 vssd1 vccd1 vccd1 _19276_/A sky130_fd_sc_hd__nand2_1
X_14994_ _20119_/A _14990_/X _14993_/X _14787_/X vssd1 vssd1 vccd1 vccd1 _14994_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19521_ _25643_/Q _19523_/B vssd1 vssd1 vccd1 vccd1 _19521_/X sky130_fd_sc_hd__or2_1
X_16733_ _22489_/A _16726_/X _16727_/X _16732_/X vssd1 vssd1 vccd1 vccd1 _16733_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13945_ _13945_/A vssd1 vssd1 vccd1 vccd1 _13945_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19452_ _19452_/A _19452_/B vssd1 vssd1 vccd1 vccd1 _19582_/B sky130_fd_sc_hd__xnor2_2
XFILLER_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16664_ _16669_/A vssd1 vssd1 vccd1 vccd1 _21562_/B sky130_fd_sc_hd__buf_6
XFILLER_234_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13876_ _14523_/A vssd1 vssd1 vccd1 vccd1 _13876_/X sky130_fd_sc_hd__buf_2
XFILLER_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18403_ _25506_/Q _18559_/A _18400_/X _18402_/X _18574_/A vssd1 vssd1 vccd1 vccd1
+ _18403_/X sky130_fd_sc_hd__o221a_1
X_15615_ _25741_/Q _15614_/Y _15615_/S vssd1 vssd1 vccd1 vccd1 _16620_/B sky130_fd_sc_hd__mux2_1
X_12827_ _25471_/Q _12973_/A _12825_/Y _12826_/X vssd1 vssd1 vccd1 vccd1 _12975_/A
+ sky130_fd_sc_hd__o22a_1
X_19383_ _19087_/X _19378_/X _19382_/X _18891_/X vssd1 vssd1 vccd1 vccd1 _19384_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_234_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16595_ _16962_/A vssd1 vssd1 vccd1 vccd1 _19571_/A sky130_fd_sc_hd__inv_2
XFILLER_250_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18334_ _18968_/A _18334_/B vssd1 vssd1 vccd1 vccd1 _18334_/Y sky130_fd_sc_hd__nand2_1
X_15546_ _15544_/X _15545_/X _15546_/S vssd1 vssd1 vccd1 vccd1 _15546_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12758_ _12758_/A vssd1 vssd1 vccd1 vccd1 _17444_/D sky130_fd_sc_hd__buf_4
XFILLER_277_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18265_ _18057_/X _18069_/X _18265_/S vssd1 vssd1 vccd1 vccd1 _18265_/X sky130_fd_sc_hd__mux2_1
X_15477_ _15547_/A _15474_/X _15476_/X _13159_/A vssd1 vssd1 vccd1 vccd1 _15477_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_202_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12689_ _12808_/A _25570_/Q vssd1 vssd1 vccd1 vccd1 _12799_/A sky130_fd_sc_hd__and2_1
X_17216_ _17222_/A _17216_/B vssd1 vssd1 vccd1 vccd1 _17217_/A sky130_fd_sc_hd__and2_1
X_14428_ _26621_/Q _26717_/Q _26653_/Q _25693_/Q _14520_/S _13121_/B vssd1 vssd1 vccd1
+ vccd1 _14428_/X sky130_fd_sc_hd__mux4_1
X_18196_ _17958_/X _17948_/X _18197_/S vssd1 vssd1 vccd1 vccd1 _18196_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17147_ _23363_/A _17105_/X _17146_/X _25574_/Q vssd1 vssd1 vccd1 vccd1 _17148_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_155_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14359_ _17504_/B _17971_/A _17504_/C _14359_/D vssd1 vssd1 vccd1 vccd1 _21195_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_116_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17078_ _22390_/B vssd1 vssd1 vccd1 vccd1 _17078_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16029_ _13465_/A _16012_/Y _16028_/Y _14826_/A vssd1 vssd1 vccd1 vccd1 _16029_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_257_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19719_ _19683_/X _19690_/X _19717_/X _19718_/X vssd1 vssd1 vccd1 vccd1 _19719_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_284_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20991_ _25249_/C vssd1 vssd1 vccd1 vccd1 _23211_/A sky130_fd_sc_hd__buf_6
XFILLER_225_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22730_ _23773_/A vssd1 vssd1 vccd1 vccd1 _22730_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22661_ _26333_/Q _22659_/X _22673_/S vssd1 vssd1 vccd1 vccd1 _22662_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24400_ _26299_/Q _24393_/X _24394_/X input243/X _24395_/X vssd1 vssd1 vccd1 vccd1
+ _24400_/X sky130_fd_sc_hd__a221o_1
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21612_ _21610_/X _21611_/X _21589_/X vssd1 vssd1 vccd1 vccd1 _21612_/X sky130_fd_sc_hd__a21o_1
XFILLER_80_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25380_ _25380_/A vssd1 vssd1 vccd1 vccd1 _27288_/D sky130_fd_sc_hd__clkbuf_1
X_22592_ _22580_/X _22591_/Y _22587_/X vssd1 vssd1 vccd1 vccd1 _26312_/D sky130_fd_sc_hd__a21oi_1
XFILLER_178_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24331_ _27002_/Q _27001_/Q _24331_/C vssd1 vssd1 vccd1 vccd1 _24334_/B sky130_fd_sc_hd__and3_1
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21543_ _25958_/Q _21506_/X _21542_/Y _21531_/X vssd1 vssd1 vccd1 vccd1 _25958_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_193_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27050_ _27062_/CLK _27050_/D vssd1 vssd1 vccd1 vccd1 _27050_/Q sky130_fd_sc_hd__dfxtp_1
X_24262_ _26977_/Q _24260_/B _24261_/Y vssd1 vssd1 vccd1 vccd1 _26977_/D sky130_fd_sc_hd__o21a_1
XFILLER_193_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21474_ _21414_/X _21472_/X _21473_/X vssd1 vssd1 vccd1 vccd1 _21474_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_154_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26001_ _26592_/CLK _26001_/D vssd1 vssd1 vccd1 vccd1 _26001_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_181_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23213_ _23281_/S vssd1 vssd1 vccd1 vccd1 _23222_/S sky130_fd_sc_hd__clkbuf_8
X_20425_ _20699_/A _20355_/X _20424_/X _20357_/X vssd1 vssd1 vccd1 vccd1 _20426_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_112_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24193_ _26954_/Q _24188_/B _24192_/Y vssd1 vssd1 vccd1 vccd1 _26954_/D sky130_fd_sc_hd__o21a_1
XFILLER_146_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23144_ _26521_/Q _23041_/X _23150_/S vssd1 vssd1 vccd1 vccd1 _23145_/A sky130_fd_sc_hd__mux2_1
X_20356_ _19309_/A _18092_/A _19315_/Y _20328_/X vssd1 vssd1 vccd1 vccd1 _20356_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_150_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23075_ _23075_/A vssd1 vssd1 vccd1 vccd1 _26499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_283_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20287_ _22518_/A _20286_/C _22520_/A vssd1 vssd1 vccd1 vccd1 _20287_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_122_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22026_ _22026_/A vssd1 vssd1 vccd1 vccd1 _26124_/D sky130_fd_sc_hd__clkbuf_1
X_26903_ _26903_/CLK _26903_/D vssd1 vssd1 vccd1 vccd1 _26903_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26834_ _26932_/CLK _26834_/D vssd1 vssd1 vccd1 vccd1 _26834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26765_ _27312_/CLK _26765_/D vssd1 vssd1 vccd1 vccd1 _26765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23977_ _23977_/A vssd1 vssd1 vccd1 vccd1 _26863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13730_ _25805_/Q _27239_/Q _15630_/A vssd1 vssd1 vccd1 vccd1 _13730_/X sky130_fd_sc_hd__mux2_1
X_25716_ _27329_/A _25716_/D vssd1 vssd1 vccd1 vccd1 _25716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22928_ _26440_/Q _22695_/X _22934_/S vssd1 vssd1 vccd1 vccd1 _22929_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26696_ _27310_/CLK _26696_/D vssd1 vssd1 vccd1 vccd1 _26696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25647_ _26297_/CLK _25647_/D vssd1 vssd1 vccd1 vccd1 _25647_/Q sky130_fd_sc_hd__dfxtp_1
X_13661_ _15916_/A _13653_/X _13660_/X _13529_/A vssd1 vssd1 vccd1 vccd1 _13661_/X
+ sky130_fd_sc_hd__o211a_1
X_22859_ _22859_/A vssd1 vssd1 vccd1 vccd1 _26409_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15400_ _26084_/Q _25889_/Q _16433_/S vssd1 vssd1 vccd1 vccd1 _15400_/X sky130_fd_sc_hd__mux2_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16380_ _26935_/Q _16380_/B vssd1 vssd1 vccd1 vccd1 _16380_/X sky130_fd_sc_hd__or2_1
X_13592_ _15808_/B vssd1 vssd1 vccd1 vccd1 _15820_/B sky130_fd_sc_hd__buf_2
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25578_ _26683_/CLK _25578_/D vssd1 vssd1 vccd1 vccd1 _25578_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_197_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15331_ _15331_/A vssd1 vssd1 vccd1 vccd1 _15406_/A sky130_fd_sc_hd__clkbuf_4
X_27317_ _27317_/CLK _27317_/D vssd1 vssd1 vccd1 vccd1 _27317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24529_ _27034_/Q _24506_/X _24528_/Y _24523_/X vssd1 vssd1 vccd1 vccd1 _27034_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18050_ _18048_/X _18049_/X _18050_/S vssd1 vssd1 vccd1 vccd1 _18050_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27248_ _27311_/CLK _27248_/D vssd1 vssd1 vccd1 vccd1 _27248_/Q sky130_fd_sc_hd__dfxtp_1
X_15262_ _26510_/Q _26382_/Q _15276_/S vssd1 vssd1 vccd1 vccd1 _15262_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17001_ _17042_/A vssd1 vssd1 vccd1 vccd1 _17001_/X sky130_fd_sc_hd__clkbuf_2
X_14213_ _14539_/S vssd1 vssd1 vccd1 vccd1 _14289_/S sky130_fd_sc_hd__buf_4
XFILLER_184_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15193_ _16476_/S _14833_/A _14718_/X _15192_/X vssd1 vssd1 vccd1 vccd1 _17782_/A
+ sky130_fd_sc_hd__a22o_2
X_27179_ _27196_/CLK _27179_/D vssd1 vssd1 vccd1 vccd1 _27179_/Q sky130_fd_sc_hd__dfxtp_1
X_14144_ _14602_/A _14144_/B vssd1 vssd1 vccd1 vccd1 _14144_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14075_ _14064_/X _14073_/X _14074_/X _13309_/B vssd1 vssd1 vccd1 vccd1 _14076_/C
+ sky130_fd_sc_hd__o211a_1
X_18952_ _27149_/Q _18952_/B vssd1 vssd1 vccd1 vccd1 _18952_/X sky130_fd_sc_hd__or2_1
XFILLER_140_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_94_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26297_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13026_ _13026_/A vssd1 vssd1 vccd1 vccd1 _13027_/A sky130_fd_sc_hd__clkbuf_2
X_17903_ _16043_/B _16040_/B _17933_/S vssd1 vssd1 vccd1 vccd1 _17903_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18883_ _25738_/Q _18892_/C vssd1 vssd1 vccd1 vccd1 _18883_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_79_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_23_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27259_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17834_ _18593_/B _17817_/X _17827_/Y _17833_/Y vssd1 vssd1 vccd1 vccd1 _18941_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_267_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14977_ _14593_/X _14941_/Y _14976_/Y _15079_/A vssd1 vssd1 vccd1 vccd1 _14977_/X
+ sky130_fd_sc_hd__a211o_4
X_17765_ _18138_/A _18077_/A vssd1 vssd1 vccd1 vccd1 _18303_/S sky130_fd_sc_hd__nor2_2
XFILLER_207_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19504_ _25636_/Q _19510_/B vssd1 vssd1 vccd1 vccd1 _19504_/X sky130_fd_sc_hd__or2_1
X_13928_ _13928_/A _13928_/B vssd1 vssd1 vccd1 vccd1 _13928_/Y sky130_fd_sc_hd__nand2_1
X_16716_ _25665_/Q vssd1 vssd1 vccd1 vccd1 _22480_/A sky130_fd_sc_hd__clkbuf_4
X_17696_ _17762_/B _17736_/A vssd1 vssd1 vccd1 vccd1 _17732_/A sky130_fd_sc_hd__nor2_4
XFILLER_281_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_400 _17036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_411 _17047_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_422 _12781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19435_ _27163_/Q _19465_/B vssd1 vssd1 vccd1 vccd1 _19435_/X sky130_fd_sc_hd__or2_1
X_16647_ _17597_/A _21070_/A vssd1 vssd1 vccd1 vccd1 _16647_/X sky130_fd_sc_hd__or2b_1
X_13859_ _26851_/Q _25765_/Q _14004_/S vssd1 vssd1 vccd1 vccd1 _13859_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_433 _25724_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_444 _25732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_455 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_466 _19283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_477 _14725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16578_ _17776_/A _16578_/B vssd1 vssd1 vccd1 vccd1 _19639_/A sky130_fd_sc_hd__nor2_4
X_19366_ _27129_/Q _18812_/X _19364_/X _19365_/X vssd1 vssd1 vccd1 vccd1 _19366_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_250_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_488 _23587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_499 _16792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18317_ _18315_/X _18729_/B _18317_/S vssd1 vssd1 vccd1 vccd1 _18317_/X sky130_fd_sc_hd__mux2_1
X_15529_ _15529_/A vssd1 vssd1 vccd1 vccd1 _15530_/B sky130_fd_sc_hd__inv_2
X_19297_ _19289_/X _19293_/Y _19296_/X _18738_/A vssd1 vssd1 vccd1 vccd1 _19297_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18248_ _18741_/A _18246_/X _18247_/X vssd1 vssd1 vccd1 vccd1 _18250_/B sky130_fd_sc_hd__a21oi_1
Xclkbuf_opt_12_0_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_57_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_163_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18179_ _18741_/A _18177_/X _18178_/X vssd1 vssd1 vccd1 vccd1 _18181_/B sky130_fd_sc_hd__a21oi_1
X_20210_ _25680_/Q _20233_/C vssd1 vssd1 vccd1 vccd1 _20210_/X sky130_fd_sc_hd__or2_1
XFILLER_116_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21190_ _21190_/A _21709_/B vssd1 vssd1 vccd1 vccd1 _21195_/C sky130_fd_sc_hd__or2_1
XFILLER_143_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20141_ _20141_/A _20141_/B vssd1 vssd1 vccd1 vccd1 _20141_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20072_ _20069_/Y _20070_/X _20046_/X _20049_/Y vssd1 vssd1 vccd1 vccd1 _20072_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_253_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23900_ _23741_/X _26829_/Q _23904_/S vssd1 vssd1 vccd1 vccd1 _23901_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24880_ _24878_/Y _24879_/X _24871_/X vssd1 vssd1 vccd1 vccd1 _27126_/D sky130_fd_sc_hd__a21oi_1
XFILLER_58_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23831_ _23831_/A vssd1 vssd1 vccd1 vccd1 _26798_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26550_ _27259_/CLK _26550_/D vssd1 vssd1 vccd1 vccd1 _26550_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23762_ _23762_/A vssd1 vssd1 vccd1 vccd1 _26771_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20974_ _20974_/A vssd1 vssd1 vccd1 vccd1 _25861_/D sky130_fd_sc_hd__clkinv_2
X_25501_ _25501_/CLK _25501_/D vssd1 vssd1 vccd1 vccd1 _25501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22713_ _22713_/A vssd1 vssd1 vccd1 vccd1 _26349_/D sky130_fd_sc_hd__clkbuf_1
X_26481_ _27288_/CLK _26481_/D vssd1 vssd1 vccd1 vccd1 _26481_/Q sky130_fd_sc_hd__dfxtp_1
X_23693_ _23693_/A vssd1 vssd1 vccd1 vccd1 _23693_/X sky130_fd_sc_hd__buf_2
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25432_ _25432_/A vssd1 vssd1 vccd1 vccd1 _27311_/D sky130_fd_sc_hd__clkbuf_1
X_22644_ _22743_/S vssd1 vssd1 vccd1 vccd1 _22657_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_213_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25363_ _27281_/Q _23744_/A _25365_/S vssd1 vssd1 vccd1 vccd1 _25364_/A sky130_fd_sc_hd__mux2_1
X_22575_ _22567_/X _22573_/Y _22574_/X vssd1 vssd1 vccd1 vccd1 _26305_/D sky130_fd_sc_hd__a21oi_1
XFILLER_178_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27102_ _27173_/CLK _27102_/D vssd1 vssd1 vccd1 vccd1 _27102_/Q sky130_fd_sc_hd__dfxtp_2
X_24314_ _24938_/A vssd1 vssd1 vccd1 vccd1 _24314_/X sky130_fd_sc_hd__buf_4
XFILLER_222_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21526_ _21480_/X _21525_/X _21473_/X vssd1 vssd1 vccd1 vccd1 _21526_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_139_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25294_ _25294_/A vssd1 vssd1 vccd1 vccd1 _27250_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27033_ _27133_/CLK _27033_/D vssd1 vssd1 vccd1 vccd1 _27033_/Q sky130_fd_sc_hd__dfxtp_1
X_24245_ _26971_/Q _24243_/B _24244_/Y vssd1 vssd1 vccd1 vccd1 _26971_/D sky130_fd_sc_hd__o21a_1
X_21457_ _21455_/X _21456_/X _21290_/A vssd1 vssd1 vccd1 vccd1 _21457_/X sky130_fd_sc_hd__a21o_1
XFILLER_182_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20408_ _19796_/X _20407_/Y _20208_/A vssd1 vssd1 vccd1 vccd1 _20408_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24176_ _24188_/A _24176_/B vssd1 vssd1 vccd1 vccd1 _24176_/Y sky130_fd_sc_hd__nor2_1
X_21388_ _21383_/Y _21387_/X _21359_/X vssd1 vssd1 vccd1 vccd1 _21388_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_162_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23127_ _23600_/A vssd1 vssd1 vccd1 vccd1 _23127_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20339_ _20339_/A _20339_/B vssd1 vssd1 vccd1 vccd1 _20343_/A sky130_fd_sc_hd__or2_1
XFILLER_122_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23058_ _26494_/Q _23057_/X _23067_/S vssd1 vssd1 vccd1 vccd1 _23059_/A sky130_fd_sc_hd__mux2_1
XTAP_5311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput100 dout0[61] vssd1 vssd1 vccd1 vccd1 input100/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput111 dout1[13] vssd1 vssd1 vccd1 vccd1 input111/X sky130_fd_sc_hd__clkbuf_1
XTAP_5333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput122 dout1[23] vssd1 vssd1 vccd1 vccd1 input122/X sky130_fd_sc_hd__clkbuf_1
X_14900_ _15003_/S vssd1 vssd1 vccd1 vccd1 _14981_/S sky130_fd_sc_hd__buf_2
XTAP_5344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22009_ _22009_/A vssd1 vssd1 vccd1 vccd1 _26116_/D sky130_fd_sc_hd__clkbuf_1
Xinput133 dout1[33] vssd1 vssd1 vccd1 vccd1 input133/X sky130_fd_sc_hd__clkbuf_2
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _13890_/X _26109_/Q _26010_/Q _13706_/A _13611_/A vssd1 vssd1 vccd1 vccd1
+ _15880_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput144 dout1[43] vssd1 vssd1 vccd1 vccd1 input144/X sky130_fd_sc_hd__clkbuf_2
XTAP_5355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput155 dout1[53] vssd1 vssd1 vccd1 vccd1 input155/X sky130_fd_sc_hd__clkbuf_2
XTAP_5366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput166 dout1[63] vssd1 vssd1 vccd1 vccd1 input166/X sky130_fd_sc_hd__clkbuf_2
XTAP_5377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput177 irq[15] vssd1 vssd1 vccd1 vccd1 input177/X sky130_fd_sc_hd__buf_6
X_14831_ _14831_/A _17779_/A vssd1 vssd1 vccd1 vccd1 _14832_/B sky130_fd_sc_hd__and2_1
XFILLER_248_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26817_ _27303_/CLK _26817_/D vssd1 vssd1 vccd1 vccd1 _26817_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput188 jtag_tdi vssd1 vssd1 vccd1 vccd1 input188/X sky130_fd_sc_hd__buf_12
Xinput199 localMemory_wb_adr_i[18] vssd1 vssd1 vccd1 vccd1 input199/X sky130_fd_sc_hd__clkbuf_1
XFILLER_236_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17550_ _17634_/A vssd1 vssd1 vccd1 vccd1 _17575_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26748_ _26813_/CLK _26748_/D vssd1 vssd1 vccd1 vccd1 _26748_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14762_ _16336_/A vssd1 vssd1 vccd1 vccd1 _14763_/A sky130_fd_sc_hd__buf_2
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16501_ _25900_/Q _16501_/B vssd1 vssd1 vccd1 vccd1 _16501_/X sky130_fd_sc_hd__or2_1
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _26660_/Q _25700_/Q _15548_/S vssd1 vssd1 vccd1 vccd1 _13713_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17481_ _26063_/Q _21209_/B _21212_/B vssd1 vssd1 vccd1 vccd1 _17482_/B sky130_fd_sc_hd__or3b_1
XFILLER_44_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26679_ _26903_/CLK _26679_/D vssd1 vssd1 vccd1 vccd1 _26679_/Q sky130_fd_sc_hd__dfxtp_1
X_14693_ _14691_/X _14692_/X _14693_/S vssd1 vssd1 vccd1 vccd1 _14693_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19220_ _25525_/Q _18439_/A _18441_/A _25557_/Q vssd1 vssd1 vccd1 vccd1 _19220_/X
+ sky130_fd_sc_hd__a22o_1
X_16432_ _14818_/A _16421_/X _16424_/X _16431_/X vssd1 vssd1 vccd1 vccd1 _16432_/X
+ sky130_fd_sc_hd__a31o_1
X_13644_ _13644_/A vssd1 vssd1 vccd1 vccd1 _13644_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_141_wb_clk_i clkbuf_opt_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25599_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_260_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19151_ _12760_/B _18972_/X _18973_/X _19150_/Y vssd1 vssd1 vccd1 vccd1 _19151_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_198_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _15085_/A _16361_/X _16362_/X _15333_/X vssd1 vssd1 vccd1 vccd1 _16363_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_197_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13575_ _12868_/Y _12941_/Y _14325_/S vssd1 vssd1 vccd1 vccd1 _13575_/X sky130_fd_sc_hd__a21o_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18102_ _18102_/A _18119_/A vssd1 vssd1 vccd1 vccd1 _18103_/A sky130_fd_sc_hd__or2_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _25819_/Q _27253_/Q _16433_/S vssd1 vssd1 vccd1 vccd1 _15314_/X sky130_fd_sc_hd__mux2_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19082_ _19146_/C _19082_/B vssd1 vssd1 vccd1 vccd1 _19082_/X sky130_fd_sc_hd__or2_2
XFILLER_8_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16294_ _14601_/A _16292_/Y _16293_/X vssd1 vssd1 vccd1 vccd1 _16294_/X sky130_fd_sc_hd__o21a_1
XFILLER_75_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18033_ _17979_/Y _17971_/X _17978_/A _17219_/A vssd1 vssd1 vccd1 vccd1 _18356_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_185_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15245_ _15245_/A vssd1 vssd1 vccd1 vccd1 _15245_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15176_ _15172_/X _15173_/X _16397_/S vssd1 vssd1 vccd1 vccd1 _15176_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14127_ _17801_/B _14127_/B vssd1 vssd1 vccd1 vccd1 _14128_/B sky130_fd_sc_hd__nor2_1
XFILLER_114_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19984_ _20080_/A _19984_/B vssd1 vssd1 vccd1 vccd1 _20007_/B sky130_fd_sc_hd__nor2_2
XFILLER_140_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14058_ _16006_/A _14053_/X _14057_/X _13210_/A vssd1 vssd1 vccd1 vccd1 _14058_/X
+ sky130_fd_sc_hd__o211a_1
X_18935_ _25613_/Q _18719_/X _18934_/X _18790_/X vssd1 vssd1 vccd1 vccd1 _25613_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13009_ _13009_/A vssd1 vssd1 vccd1 vccd1 _13010_/A sky130_fd_sc_hd__clkbuf_2
X_18866_ _25515_/Q _18807_/X _18808_/X _17384_/X vssd1 vssd1 vccd1 vccd1 _18866_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_255_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17817_ _16735_/A _17816_/X _18593_/A _17817_/D vssd1 vssd1 vccd1 vccd1 _17817_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_282_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18797_ _18799_/A _18211_/X _17988_/A _18681_/A vssd1 vssd1 vccd1 vccd1 _18803_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_54_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17748_ _18102_/A _17749_/B vssd1 vssd1 vccd1 vccd1 _18234_/A sky130_fd_sc_hd__nor2_2
XFILLER_54_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_230 _19971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17679_ _17679_/A _17679_/B _17670_/C vssd1 vssd1 vccd1 vccd1 _18094_/A sky130_fd_sc_hd__or3b_2
XFILLER_23_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_241 _21070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_252 _16822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19418_ _17443_/A _18720_/X _18788_/X _19417_/Y vssd1 vssd1 vccd1 vccd1 _19418_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_250_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_263 _22535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20690_ _20690_/A _20703_/B vssd1 vssd1 vccd1 vccd1 _20690_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_274 _25484_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_285 _25818_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_296 _25827_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19349_ _18929_/X _19345_/X _19348_/X _18782_/X vssd1 vssd1 vccd1 vccd1 _19349_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22360_ _22393_/A _26237_/Q _22360_/C vssd1 vssd1 vccd1 vccd1 _22388_/A sky130_fd_sc_hd__and3_1
XFILLER_248_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21311_ _25473_/Q _21332_/B vssd1 vssd1 vccd1 vccd1 _21311_/X sky130_fd_sc_hd__or2_1
XFILLER_108_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22291_ _26209_/Q _22284_/X _22290_/X _22288_/X vssd1 vssd1 vccd1 vccd1 _26209_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_190_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24030_ _24030_/A vssd1 vssd1 vccd1 vccd1 _26886_/D sky130_fd_sc_hd__clkbuf_1
X_21242_ _24871_/A vssd1 vssd1 vccd1 vccd1 _21242_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_144_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21173_ _21173_/A vssd1 vssd1 vccd1 vccd1 _25928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20124_ _20125_/A _20125_/B _20125_/D _20125_/C vssd1 vssd1 vccd1 vccd1 _20126_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_131_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25981_ _25985_/CLK _25981_/D vssd1 vssd1 vccd1 vccd1 _25981_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24932_ _24932_/A _24951_/B vssd1 vssd1 vccd1 vccd1 _24932_/Y sky130_fd_sc_hd__nand2_1
X_20055_ _20055_/A _20055_/B vssd1 vssd1 vccd1 vccd1 _20055_/X sky130_fd_sc_hd__or2_1
XFILLER_86_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24863_ _27122_/Q _24873_/B vssd1 vssd1 vccd1 vccd1 _24863_/Y sky130_fd_sc_hd__nand2_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26602_ _27305_/CLK _26602_/D vssd1 vssd1 vccd1 vccd1 _26602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23814_ _23814_/A vssd1 vssd1 vccd1 vccd1 _26790_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24794_ _27104_/Q _24798_/B vssd1 vssd1 vccd1 vccd1 _24794_/Y sky130_fd_sc_hd__nand2_1
XFILLER_273_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26533_ _27304_/CLK _26533_/D vssd1 vssd1 vccd1 vccd1 _26533_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23745_ _23744_/X _26766_/Q _23748_/S vssd1 vssd1 vccd1 vccd1 _23746_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20957_ _20957_/A vssd1 vssd1 vccd1 vccd1 _25855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26464_ _27275_/CLK _26464_/D vssd1 vssd1 vccd1 vccd1 _26464_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_242_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23676_ _26744_/Q _23600_/X _23678_/S vssd1 vssd1 vccd1 vccd1 _23677_/A sky130_fd_sc_hd__mux2_1
X_20888_ _20971_/S vssd1 vssd1 vccd1 vccd1 _20901_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25415_ _23715_/X _27304_/Q _25415_/S vssd1 vssd1 vccd1 vccd1 _25416_/A sky130_fd_sc_hd__mux2_1
X_22627_ _17447_/B _22625_/X _22419_/D _22629_/A vssd1 vssd1 vccd1 vccd1 _22638_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_201_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26395_ _27267_/CLK _26395_/D vssd1 vssd1 vccd1 vccd1 _26395_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_139_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25346_ _27273_/Q _23718_/A _25354_/S vssd1 vssd1 vccd1 vccd1 _25347_/A sky130_fd_sc_hd__mux2_1
X_13360_ _14741_/A _26919_/Q _26403_/Q _15299_/S _13359_/X vssd1 vssd1 vccd1 vccd1
+ _13360_/X sky130_fd_sc_hd__a221o_1
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22558_ _26299_/Q _22565_/B vssd1 vssd1 vccd1 vccd1 _22558_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21509_ _21586_/A vssd1 vssd1 vccd1 vccd1 _21509_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25277_ _25277_/A vssd1 vssd1 vccd1 vccd1 _27242_/D sky130_fd_sc_hd__clkbuf_1
X_13291_ _13291_/A vssd1 vssd1 vccd1 vccd1 _13291_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22489_ _22489_/A _22491_/B vssd1 vssd1 vccd1 vccd1 _22490_/A sky130_fd_sc_hd__and2_1
X_27016_ _27049_/CLK _27016_/D vssd1 vssd1 vccd1 vccd1 _27016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15030_ _26514_/Q _26386_/Q _15030_/S vssd1 vssd1 vccd1 vccd1 _15030_/X sky130_fd_sc_hd__mux2_1
X_24228_ _24237_/A _24233_/C vssd1 vssd1 vccd1 vccd1 _24228_/Y sky130_fd_sc_hd__nor2_1
XFILLER_181_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24159_ _24159_/A _24159_/B vssd1 vssd1 vccd1 vccd1 _26943_/D sky130_fd_sc_hd__nor2_1
XFILLER_218_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16981_ _16981_/A vssd1 vssd1 vccd1 vccd1 _16981_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18720_ _19218_/A vssd1 vssd1 vccd1 vccd1 _18720_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15932_ _15932_/A _15932_/B vssd1 vssd1 vccd1 vccd1 _15932_/X sky130_fd_sc_hd__or2_1
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_264_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15863_ _14727_/A _15861_/X _15862_/X _13304_/A vssd1 vssd1 vccd1 vccd1 _15863_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_209_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18651_ _18843_/D _18651_/B vssd1 vssd1 vccd1 vccd1 _18651_/Y sky130_fd_sc_hd__nor2_2
XTAP_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17602_ _20119_/A _17551_/X _17553_/X _17601_/Y vssd1 vssd1 vccd1 vccd1 _17603_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14814_ _14747_/A _26618_/Q _16510_/A _26358_/Q _14733_/A vssd1 vssd1 vccd1 vccd1
+ _14814_/X sky130_fd_sc_hd__o221a_1
XFILLER_280_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15794_ _12951_/X _15792_/X _15793_/X vssd1 vssd1 vccd1 vccd1 _15794_/X sky130_fd_sc_hd__o21a_1
X_18582_ _25732_/Q _18588_/C vssd1 vssd1 vccd1 vccd1 _18582_/X sky130_fd_sc_hd__xor2_2
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_264_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _17533_/A vssd1 vssd1 vccd1 vccd1 _17653_/A sky130_fd_sc_hd__clkbuf_2
X_14745_ _14890_/A vssd1 vssd1 vccd1 vccd1 _14746_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17464_ _26253_/Q _17453_/A _17459_/A _25981_/Q vssd1 vssd1 vccd1 vccd1 _17708_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_189_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14676_ _16479_/A _14673_/X _14675_/X _14662_/X vssd1 vssd1 vccd1 vccd1 _14676_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_32_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19203_ _27060_/Q _19055_/X _19200_/X _19202_/X _19066_/X vssd1 vssd1 vccd1 vccd1
+ _19203_/X sky130_fd_sc_hd__o221a_2
X_16415_ _15290_/A _16414_/Y _14718_/A vssd1 vssd1 vccd1 vccd1 _16415_/Y sky130_fd_sc_hd__o21ai_1
X_13627_ _26629_/Q _26725_/Q _15971_/S vssd1 vssd1 vccd1 vccd1 _13627_/X sky130_fd_sc_hd__mux2_1
X_17395_ _25550_/Q vssd1 vssd1 vccd1 vccd1 _17395_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_201_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19134_ _27026_/Q _19063_/X _19133_/X _18565_/X vssd1 vssd1 vccd1 vccd1 _19134_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16346_ _26805_/Q _26449_/Q _16347_/S vssd1 vssd1 vccd1 vccd1 _16346_/X sky130_fd_sc_hd__mux2_1
X_13558_ _13558_/A vssd1 vssd1 vccd1 vccd1 _16639_/A sky130_fd_sc_hd__buf_4
XFILLER_201_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19065_ _27024_/Q _19063_/X _19064_/X _18565_/X vssd1 vssd1 vccd1 vccd1 _19065_/X
+ sky130_fd_sc_hd__a22o_1
X_16277_ _25852_/Q _26052_/Q _16277_/S vssd1 vssd1 vccd1 vccd1 _16277_/X sky130_fd_sc_hd__mux2_1
X_13489_ _14551_/S vssd1 vssd1 vccd1 vccd1 _14307_/S sky130_fd_sc_hd__buf_2
XFILLER_218_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15228_ _26512_/Q _26384_/Q _15228_/S vssd1 vssd1 vccd1 vccd1 _15228_/X sky130_fd_sc_hd__mux2_1
X_18016_ _18016_/A vssd1 vssd1 vccd1 vccd1 _19087_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_145_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput404 _17012_/X vssd1 vssd1 vccd1 vccd1 din0[6] sky130_fd_sc_hd__buf_2
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput415 _25950_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[14] sky130_fd_sc_hd__buf_2
XFILLER_160_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput426 _25960_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[24] sky130_fd_sc_hd__buf_2
Xoutput437 _25941_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_160_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15159_ _27287_/Q _26480_/Q _16402_/S vssd1 vssd1 vccd1 vccd1 _15159_/X sky130_fd_sc_hd__mux2_1
Xoutput448 _26235_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[3] sky130_fd_sc_hd__buf_2
XFILLER_141_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput459 _25742_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[18] sky130_fd_sc_hd__buf_2
XFILLER_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19967_ _20276_/A vssd1 vssd1 vccd1 vccd1 _19967_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18918_ _27020_/Q _19063_/A _18917_/X _18565_/A vssd1 vssd1 vccd1 vccd1 _18918_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19898_ _19897_/Y _19867_/Y _19865_/Y vssd1 vssd1 vccd1 vccd1 _19898_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_267_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18849_ _16591_/A _18720_/X _18847_/Y _18848_/Y _18788_/X vssd1 vssd1 vccd1 vccd1
+ _18849_/X sky130_fd_sc_hd__a221o_4
XFILLER_83_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21860_ _26058_/Q _20964_/X _21860_/S vssd1 vssd1 vccd1 vccd1 _21861_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20811_ _20811_/A vssd1 vssd1 vccd1 vccd1 _25801_/D sky130_fd_sc_hd__clkbuf_1
X_21791_ _20621_/X _26028_/Q _21791_/S vssd1 vssd1 vccd1 vccd1 _21792_/A sky130_fd_sc_hd__mux2_1
X_23530_ _23530_/A vssd1 vssd1 vccd1 vccd1 _23530_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20742_ _20533_/X _25768_/Q _20750_/S vssd1 vssd1 vccd1 vccd1 _20743_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23461_ _26662_/Q _23069_/X _23469_/S vssd1 vssd1 vccd1 vccd1 _23462_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20673_ _20686_/A vssd1 vssd1 vccd1 vccd1 _20673_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25200_ _24690_/B _25198_/X _25196_/X _27210_/Q _25199_/X vssd1 vssd1 vccd1 vccd1
+ _27210_/D sky130_fd_sc_hd__o221a_1
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22412_ _22394_/A _22381_/X _22411_/X _22337_/X vssd1 vssd1 vccd1 vccd1 _22412_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_148_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26180_ _26319_/CLK _26180_/D vssd1 vssd1 vccd1 vccd1 _26180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23392_ _23392_/A vssd1 vssd1 vccd1 vccd1 _26631_/D sky130_fd_sc_hd__clkbuf_1
X_25131_ _24739_/Y _25124_/X _25130_/Y _25109_/X vssd1 vssd1 vccd1 vccd1 _25131_/X
+ sky130_fd_sc_hd__a31o_1
X_22343_ _17085_/A _26226_/Q _22350_/S vssd1 vssd1 vccd1 vccd1 _22343_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25062_ _20650_/A _25059_/X _25061_/X vssd1 vssd1 vccd1 vccd1 _25062_/Y sky130_fd_sc_hd__o21ai_1
X_22274_ _26203_/Q _22269_/X _22272_/X _22273_/X vssd1 vssd1 vccd1 vccd1 _26203_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24013_ _26879_/Q _23520_/X _24015_/S vssd1 vssd1 vccd1 vccd1 _24014_/A sky130_fd_sc_hd__mux2_1
X_21225_ _21885_/A _21866_/B _21244_/B _21224_/X vssd1 vssd1 vccd1 vccd1 _22536_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_137_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21156_ _21174_/A vssd1 vssd1 vccd1 vccd1 _21172_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_132_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20107_ _20069_/Y _20071_/Y _20131_/A _20105_/Y vssd1 vssd1 vccd1 vccd1 _20131_/B
+ sky130_fd_sc_hd__a211oi_1
X_25964_ _26995_/CLK _25964_/D vssd1 vssd1 vccd1 vccd1 _25964_/Q sky130_fd_sc_hd__dfxtp_1
X_21087_ _21087_/A vssd1 vssd1 vccd1 vccd1 _25904_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24915_ _24915_/A _24923_/B vssd1 vssd1 vccd1 vccd1 _24915_/Y sky130_fd_sc_hd__nand2_1
X_20038_ _20039_/A _20039_/B vssd1 vssd1 vccd1 vccd1 _20038_/X sky130_fd_sc_hd__or2_1
XFILLER_59_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_274_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25895_ _26483_/CLK _25895_/D vssd1 vssd1 vccd1 vccd1 _25895_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12860_ _12878_/B _12860_/B vssd1 vssd1 vccd1 vccd1 _12933_/B sky130_fd_sc_hd__or2_2
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24846_ _24844_/Y _24845_/X _24835_/X vssd1 vssd1 vccd1 vccd1 _27117_/D sky130_fd_sc_hd__a21oi_1
XFILLER_274_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24777_ _24777_/A _24777_/B vssd1 vssd1 vccd1 vccd1 _24801_/A sky130_fd_sc_hd__nor2_4
XFILLER_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _25596_/Q _25594_/Q _12790_/X _12808_/A vssd1 vssd1 vccd1 vccd1 _17978_/A
+ sky130_fd_sc_hd__o31a_4
X_21989_ _21989_/A vssd1 vssd1 vccd1 vccd1 _26107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14453_/X _25829_/Q _26029_/Q _13841_/A _13336_/A vssd1 vssd1 vccd1 vccd1
+ _14530_/X sky130_fd_sc_hd__a221o_1
XFILLER_42_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26516_ _27324_/CLK _26516_/D vssd1 vssd1 vccd1 vccd1 _26516_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23728_ _23728_/A vssd1 vssd1 vccd1 vccd1 _23728_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14043_/X _14459_/X _14460_/X _13773_/A vssd1 vssd1 vccd1 vccd1 _14461_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26447_ _27287_/CLK _26447_/D vssd1 vssd1 vccd1 vccd1 _26447_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23659_ _26736_/Q _23574_/X _23667_/S vssd1 vssd1 vccd1 vccd1 _23660_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16200_ _14807_/A _16188_/X _16192_/X _16199_/X _14786_/A vssd1 vssd1 vccd1 vccd1
+ _16200_/X sky130_fd_sc_hd__a311o_1
X_13412_ _15807_/S vssd1 vssd1 vccd1 vccd1 _15471_/S sky130_fd_sc_hd__clkbuf_4
X_17180_ _25486_/Q _17159_/X _17179_/Y _17175_/X vssd1 vssd1 vccd1 vccd1 _25486_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26378_ _27281_/CLK _26378_/D vssd1 vssd1 vccd1 vccd1 _26378_/Q sky130_fd_sc_hd__dfxtp_1
X_14392_ _12736_/A _26878_/Q _26750_/Q _14536_/S _14384_/X vssd1 vssd1 vccd1 vccd1
+ _14392_/X sky130_fd_sc_hd__a221o_1
XFILLER_183_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16131_ _14600_/A _16129_/Y _16130_/X _15135_/A vssd1 vssd1 vccd1 vccd1 _16131_/X
+ sky130_fd_sc_hd__o22a_1
X_25329_ _25329_/A vssd1 vssd1 vccd1 vccd1 _27265_/D sky130_fd_sc_hd__clkbuf_1
X_13343_ _14473_/S vssd1 vssd1 vccd1 vccd1 _13344_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16062_ _26083_/Q _15623_/B _14713_/B _16061_/X vssd1 vssd1 vccd1 vccd1 _16062_/X
+ sky130_fd_sc_hd__o211a_1
X_13274_ _13274_/A vssd1 vssd1 vccd1 vccd1 _13274_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_182_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15013_ _17851_/A _17850_/A vssd1 vssd1 vccd1 vccd1 _16560_/A sky130_fd_sc_hd__nand2_2
XFILLER_269_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19821_ _19748_/X _19820_/X _19755_/X vssd1 vssd1 vccd1 vccd1 _19821_/X sky130_fd_sc_hd__a21o_1
XFILLER_269_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19752_ _19750_/Y _19752_/B vssd1 vssd1 vccd1 vccd1 _19753_/B sky130_fd_sc_hd__and2b_1
XFILLER_231_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16964_ _16862_/X _16954_/X _16956_/X _16860_/X _16963_/X vssd1 vssd1 vccd1 vccd1
+ _16965_/C sky130_fd_sc_hd__a221o_1
XFILLER_77_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18703_ _19947_/A _19268_/B vssd1 vssd1 vccd1 vccd1 _18703_/Y sky130_fd_sc_hd__nor2_1
X_15915_ _26533_/Q _26141_/Q _15915_/S vssd1 vssd1 vccd1 vccd1 _15916_/B sky130_fd_sc_hd__mux2_1
X_19683_ _24810_/A vssd1 vssd1 vccd1 vccd1 _19683_/X sky130_fd_sc_hd__buf_2
XFILLER_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16895_ _16895_/A vssd1 vssd1 vccd1 vccd1 _16924_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18634_ _18634_/A _18634_/B _16735_/A vssd1 vssd1 vccd1 vccd1 _18635_/B sky130_fd_sc_hd__or3b_1
XFILLER_253_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15846_ _15589_/A _27277_/Q _26470_/Q _15914_/S _15859_/A vssd1 vssd1 vccd1 vccd1
+ _15846_/X sky130_fd_sc_hd__a221o_1
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18565_ _18565_/A vssd1 vssd1 vccd1 vccd1 _18565_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_280_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15777_ _13359_/A _15774_/X _15776_/X _13339_/A vssd1 vssd1 vccd1 vccd1 _15777_/X
+ sky130_fd_sc_hd__o211a_1
X_12989_ _12989_/A vssd1 vssd1 vccd1 vccd1 _13139_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17516_ _19636_/A vssd1 vssd1 vccd1 vccd1 _17516_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14728_ _16195_/S vssd1 vssd1 vccd1 vccd1 _14729_/A sky130_fd_sc_hd__clkbuf_4
X_18496_ _17920_/X _17897_/X _18271_/X vssd1 vssd1 vccd1 vccd1 _18496_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_205_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17447_ _26327_/Q _17447_/B vssd1 vssd1 vccd1 vccd1 _21868_/A sky130_fd_sc_hd__and2_2
XFILLER_232_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14659_ _14659_/A vssd1 vssd1 vccd1 vccd1 _14660_/A sky130_fd_sc_hd__buf_4
XFILLER_165_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17378_ _17375_/X _17379_/C _25545_/Q vssd1 vssd1 vccd1 vccd1 _17380_/B sky130_fd_sc_hd__a21oi_1
XFILLER_193_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19117_ _19317_/A _19117_/B vssd1 vssd1 vccd1 vccd1 _19117_/Y sky130_fd_sc_hd__nand2_1
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16329_ _15285_/A _16324_/X _16328_/Y _14706_/A vssd1 vssd1 vccd1 vccd1 _16329_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19048_ _19048_/A _19048_/B vssd1 vssd1 vccd1 vccd1 _19579_/B sky130_fd_sc_hd__xnor2_2
XFILLER_173_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21010_ _21010_/A vssd1 vssd1 vccd1 vccd1 _25875_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput289 _17067_/X vssd1 vssd1 vccd1 vccd1 addr0[4] sky130_fd_sc_hd__buf_2
XFILLER_275_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_7 _22368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22961_ _22961_/A vssd1 vssd1 vccd1 vccd1 _26455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24700_ _24723_/A vssd1 vssd1 vccd1 vccd1 _24722_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21912_ _21912_/A vssd1 vssd1 vccd1 vccd1 _26073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25680_ _26278_/CLK _25680_/D vssd1 vssd1 vccd1 vccd1 _25680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22892_ _22960_/S vssd1 vssd1 vccd1 vccd1 _22901_/S sky130_fd_sc_hd__buf_2
XFILLER_167_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24631_ _25221_/A vssd1 vssd1 vccd1 vccd1 _24631_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21843_ _26050_/Q _20939_/X _21849_/S vssd1 vssd1 vccd1 vccd1 _21844_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24562_ _24615_/A vssd1 vssd1 vccd1 vccd1 _24562_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_169_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21774_ _20588_/X _26020_/Q _21776_/S vssd1 vssd1 vccd1 vccd1 _21775_/A sky130_fd_sc_hd__mux2_1
X_26301_ _26327_/CLK _26301_/D vssd1 vssd1 vccd1 vccd1 _26301_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_24_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23513_ _23513_/A vssd1 vssd1 vccd1 vccd1 _26684_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20725_ _20725_/A vssd1 vssd1 vccd1 vccd1 _25760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27281_ _27281_/CLK _27281_/D vssd1 vssd1 vccd1 vccd1 _27281_/Q sky130_fd_sc_hd__dfxtp_1
X_24493_ _27027_/Q _24480_/X _24492_/Y _24470_/X vssd1 vssd1 vccd1 vccd1 _27027_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26232_ _27297_/CLK _26232_/D vssd1 vssd1 vccd1 vccd1 _26232_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23444_ _23444_/A vssd1 vssd1 vccd1 vccd1 _26654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20656_ _20656_/A _20656_/B vssd1 vssd1 vccd1 vccd1 _20656_/X sky130_fd_sc_hd__or2_1
XFILLER_149_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26163_ _27264_/CLK _26163_/D vssd1 vssd1 vccd1 vccd1 _26163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23375_ _26624_/Q _23050_/X _23375_/S vssd1 vssd1 vccd1 vccd1 _23376_/A sky130_fd_sc_hd__mux2_1
X_20587_ _23584_/A vssd1 vssd1 vccd1 vccd1 _23760_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25114_ _25114_/A vssd1 vssd1 vccd1 vccd1 _25114_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22326_ _26221_/Q _22315_/X _22325_/X _22319_/X vssd1 vssd1 vccd1 vccd1 _26221_/D
+ sky130_fd_sc_hd__o211a_1
X_26094_ _27293_/CLK _26094_/D vssd1 vssd1 vccd1 vccd1 _26094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25045_ _20641_/A _25031_/X _25044_/X vssd1 vssd1 vccd1 vccd1 _25045_/Y sky130_fd_sc_hd__o21ai_1
X_22257_ _26197_/Q _22249_/X _22255_/X _26298_/Q _22256_/X vssd1 vssd1 vccd1 vccd1
+ _22257_/X sky130_fd_sc_hd__a221o_1
XFILLER_152_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21208_ _21208_/A _21208_/B _21219_/A _21208_/D vssd1 vssd1 vccd1 vccd1 _21218_/D
+ sky130_fd_sc_hd__nor4_1
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22188_ _26179_/Q _22186_/X _22179_/X input278/X _22187_/X vssd1 vssd1 vccd1 vccd1
+ _22188_/X sky130_fd_sc_hd__a221o_1
XFILLER_160_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21139_ _25919_/Q _21130_/X _21131_/X input18/X vssd1 vssd1 vccd1 vccd1 _21140_/B
+ sky130_fd_sc_hd__o22a_1
X_26996_ _26996_/CLK _26996_/D vssd1 vssd1 vccd1 vccd1 _26996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_266_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13961_ _13958_/X _13959_/X _14309_/S vssd1 vssd1 vccd1 vccd1 _13961_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25947_ _25985_/CLK _25947_/D vssd1 vssd1 vccd1 vccd1 _25947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12912_ _12912_/A vssd1 vssd1 vccd1 vccd1 _12913_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15700_ _17837_/A _15701_/B vssd1 vssd1 vccd1 vccd1 _18938_/S sky130_fd_sc_hd__nand2_2
XFILLER_111_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16680_ _16676_/A _16676_/B _20978_/B vssd1 vssd1 vccd1 vccd1 _17060_/A sky130_fd_sc_hd__o21a_1
X_25878_ _27307_/CLK _25878_/D vssd1 vssd1 vccd1 vccd1 _25878_/Q sky130_fd_sc_hd__dfxtp_2
X_13892_ _14433_/S vssd1 vssd1 vccd1 vccd1 _14257_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_219_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12843_ _12891_/A _13389_/A _17623_/C _12899_/A _25925_/Q vssd1 vssd1 vccd1 vccd1
+ _15704_/A sky130_fd_sc_hd__o32a_4
X_15631_ _26344_/Q _26604_/Q _15643_/S vssd1 vssd1 vccd1 vccd1 _15631_/X sky130_fd_sc_hd__mux2_1
X_24829_ _24848_/A vssd1 vssd1 vccd1 vccd1 _24829_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15562_ _25709_/Q _16310_/B _15561_/X _15168_/A vssd1 vssd1 vccd1 vccd1 _15562_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18350_ _18362_/A _18350_/B vssd1 vssd1 vccd1 vccd1 _18350_/X sky130_fd_sc_hd__or2_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12774_/A vssd1 vssd1 vccd1 vccd1 _12775_/A sky130_fd_sc_hd__buf_2
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _26096_/Q _25997_/Q _14513_/S vssd1 vssd1 vccd1 vccd1 _14513_/X sky130_fd_sc_hd__mux2_1
X_17301_ _17299_/X _17303_/C _17300_/Y vssd1 vssd1 vccd1 vccd1 _25520_/D sky130_fd_sc_hd__o21a_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_48_wb_clk_i clkbuf_leaf_48_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _27281_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15493_ _15491_/X _26894_/Q _26766_/Q _15834_/S _15852_/A vssd1 vssd1 vccd1 vccd1
+ _15493_/X sky130_fd_sc_hd__a221o_1
X_18281_ _18968_/A _18281_/B vssd1 vssd1 vccd1 vccd1 _18281_/Y sky130_fd_sc_hd__nand2_1
XFILLER_261_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17232_ _25502_/Q vssd1 vssd1 vccd1 vccd1 _17242_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14444_ _16813_/B _16813_/C _16578_/B vssd1 vssd1 vccd1 vccd1 _14444_/X sky130_fd_sc_hd__a21o_1
XFILLER_230_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17163_ _25480_/Q _17159_/X _17162_/Y _17134_/X vssd1 vssd1 vccd1 vccd1 _25480_/D
+ sky130_fd_sc_hd__o211a_1
X_14375_ _25799_/Q _27233_/Q _14375_/S vssd1 vssd1 vccd1 vccd1 _14375_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16114_ _13255_/A _26927_/Q _26411_/Q _16260_/S _13330_/A vssd1 vssd1 vccd1 vccd1
+ _16114_/X sky130_fd_sc_hd__a221o_1
X_13326_ _15321_/A _26107_/Q _26008_/Q _16267_/S _13321_/A vssd1 vssd1 vccd1 vccd1
+ _13326_/X sky130_fd_sc_hd__a221o_1
X_17094_ _22121_/A _17094_/B _26191_/Q vssd1 vssd1 vccd1 vccd1 _17094_/X sky130_fd_sc_hd__and3b_1
XFILLER_170_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16045_ _15245_/X _12926_/X _14603_/A vssd1 vssd1 vccd1 vccd1 _16045_/Y sky130_fd_sc_hd__a21oi_1
X_13257_ _14054_/A vssd1 vssd1 vccd1 vccd1 _14551_/S sky130_fd_sc_hd__buf_2
XFILLER_97_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13188_ _14060_/A vssd1 vssd1 vccd1 vccd1 _14459_/S sky130_fd_sc_hd__buf_2
XFILLER_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19804_ _19805_/A _19805_/B vssd1 vssd1 vccd1 vccd1 _19804_/X sky130_fd_sc_hd__and2_1
XFILLER_111_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17996_ _18308_/B vssd1 vssd1 vccd1 vccd1 _17997_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19735_ _19853_/A _19736_/B vssd1 vssd1 vccd1 vccd1 _19737_/A sky130_fd_sc_hd__and2_1
XFILLER_284_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16947_ _16957_/A _16896_/X _16938_/X _16847_/A _16946_/Y vssd1 vssd1 vccd1 vccd1
+ _16948_/B sky130_fd_sc_hd__o221a_1
XFILLER_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19666_ _19882_/B _18150_/X _19663_/X _19665_/X vssd1 vssd1 vccd1 vccd1 _19666_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_226_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16878_ _16910_/A _16878_/B vssd1 vssd1 vccd1 vccd1 _16878_/X sky130_fd_sc_hd__or2_1
XFILLER_280_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18617_ _27014_/Q _18514_/A _18616_/X _18455_/A vssd1 vssd1 vccd1 vccd1 _18617_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15829_ _15812_/X _15828_/X _13174_/A vssd1 vssd1 vccd1 vccd1 _15830_/B sky130_fd_sc_hd__a21oi_4
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19597_ _20125_/A vssd1 vssd1 vccd1 vccd1 _19676_/A sky130_fd_sc_hd__buf_2
XFILLER_240_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18548_ _18548_/A vssd1 vssd1 vccd1 vccd1 _18548_/X sky130_fd_sc_hd__buf_4
XFILLER_52_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18479_ _18630_/A _18479_/B vssd1 vssd1 vccd1 vccd1 _18480_/A sky130_fd_sc_hd__and2_1
XFILLER_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20510_ _20510_/A vssd1 vssd1 vccd1 vccd1 _25696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21490_ _21490_/A vssd1 vssd1 vccd1 vccd1 _21490_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20441_ _25690_/Q vssd1 vssd1 vccd1 vccd1 _22533_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23160_ _23160_/A vssd1 vssd1 vccd1 vccd1 _26528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20372_ _20179_/X _20371_/X _20186_/X vssd1 vssd1 vccd1 vccd1 _20372_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22111_ _26230_/Q _22236_/C vssd1 vssd1 vccd1 vccd1 _22170_/A sky130_fd_sc_hd__nand2_2
XFILLER_133_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23091_ _23091_/A vssd1 vssd1 vccd1 vccd1 _26504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22042_ _26131_/Q _20881_/X _22044_/S vssd1 vssd1 vccd1 vccd1 _22043_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26850_ _26917_/CLK _26850_/D vssd1 vssd1 vccd1 vccd1 _26850_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25801_ _26520_/CLK _25801_/D vssd1 vssd1 vccd1 vccd1 _25801_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26781_ _27295_/CLK _26781_/D vssd1 vssd1 vccd1 vccd1 _26781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23993_ _23993_/A vssd1 vssd1 vccd1 vccd1 _26870_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25732_ _26271_/CLK _25732_/D vssd1 vssd1 vccd1 vccd1 _25732_/Q sky130_fd_sc_hd__dfxtp_4
X_22944_ _22944_/A vssd1 vssd1 vccd1 vccd1 _26447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25663_ _26264_/CLK _25663_/D vssd1 vssd1 vccd1 vccd1 _25663_/Q sky130_fd_sc_hd__dfxtp_1
X_22875_ _22875_/A vssd1 vssd1 vccd1 vccd1 _22884_/S sky130_fd_sc_hd__buf_4
XFILLER_245_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24614_ _27061_/Q _24602_/X _24613_/Y _24606_/X vssd1 vssd1 vccd1 vccd1 _27061_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21826_ _21826_/A vssd1 vssd1 vccd1 vccd1 _26042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25594_ _25596_/CLK _25594_/D vssd1 vssd1 vccd1 vccd1 _25594_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24545_ _24561_/A vssd1 vssd1 vccd1 vccd1 _24629_/B sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21757_ _20554_/X _26012_/Q _21765_/S vssd1 vssd1 vccd1 vccd1 _21758_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27264_ _27264_/CLK _27264_/D vssd1 vssd1 vccd1 vccd1 _27264_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20708_ _20712_/B _26261_/D _20707_/X _19991_/X vssd1 vssd1 vccd1 vccd1 _25756_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24476_ _24472_/X _25617_/Q _24475_/X vssd1 vssd1 vccd1 vccd1 _24725_/B sky130_fd_sc_hd__o21a_4
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21688_ _25983_/Q input195/X _21696_/S vssd1 vssd1 vccd1 vccd1 _21689_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26215_ _26319_/CLK _26215_/D vssd1 vssd1 vccd1 vccd1 _26215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23427_ _23427_/A vssd1 vssd1 vccd1 vccd1 _26647_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20639_ _20639_/A _20643_/B vssd1 vssd1 vccd1 vccd1 _20639_/X sky130_fd_sc_hd__or2_1
X_27195_ _27198_/CLK _27195_/D vssd1 vssd1 vccd1 vccd1 _27195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14160_ _25833_/Q _26033_/Q _15902_/S vssd1 vssd1 vccd1 vccd1 _14160_/X sky130_fd_sc_hd__mux2_1
X_26146_ _26531_/CLK _26146_/D vssd1 vssd1 vccd1 vccd1 _26146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23358_ _23358_/A vssd1 vssd1 vccd1 vccd1 _26617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13111_ _14354_/S vssd1 vssd1 vccd1 vccd1 _13112_/A sky130_fd_sc_hd__buf_2
XFILLER_137_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22309_ _26215_/Q _22299_/X _22308_/X _22304_/X vssd1 vssd1 vccd1 vccd1 _26215_/D
+ sky130_fd_sc_hd__o211a_1
X_26077_ _26601_/CLK _26077_/D vssd1 vssd1 vccd1 vccd1 _26077_/Q sky130_fd_sc_hd__dfxtp_1
X_14091_ _25834_/Q _26034_/Q _14114_/S vssd1 vssd1 vccd1 vccd1 _14091_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23289_ _26587_/Q input250/X _23289_/S vssd1 vssd1 vccd1 vccd1 _23290_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_166_wb_clk_i clkbuf_opt_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26286_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13042_ _15888_/S vssd1 vssd1 vccd1 vccd1 _13043_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25028_ _24659_/Y _25014_/X _25026_/Y _25027_/X vssd1 vssd1 vccd1 vccd1 _25028_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17850_ _17850_/A vssd1 vssd1 vccd1 vccd1 _17851_/B sky130_fd_sc_hd__inv_2
XFILLER_266_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16801_ _16801_/A vssd1 vssd1 vccd1 vccd1 _16906_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17781_ _17781_/A vssd1 vssd1 vccd1 vccd1 _17782_/B sky130_fd_sc_hd__inv_2
X_26979_ _26980_/CLK _26979_/D vssd1 vssd1 vccd1 vccd1 _26979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_254_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14993_ _14766_/A _14991_/X _14992_/X _14760_/A vssd1 vssd1 vccd1 vccd1 _14993_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19520_ _19512_/X _18772_/X _19519_/X _19515_/X vssd1 vssd1 vccd1 vccd1 _25642_/D
+ sky130_fd_sc_hd__o211a_1
X_16732_ _18593_/A _16732_/B vssd1 vssd1 vccd1 vccd1 _16732_/X sky130_fd_sc_hd__xor2_4
XFILLER_247_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13944_ _13937_/X _26690_/Q _26818_/Q _15759_/S _13943_/X vssd1 vssd1 vccd1 vccd1
+ _13944_/X sky130_fd_sc_hd__a221o_1
XFILLER_74_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19451_ _25628_/Q _18719_/A _19450_/X _19352_/X vssd1 vssd1 vccd1 vccd1 _25628_/D
+ sky130_fd_sc_hd__o211a_1
X_13875_ _13857_/X _13868_/X _13874_/X _13163_/A vssd1 vssd1 vccd1 vccd1 _13875_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_223_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16663_ _25996_/Q _25995_/Q vssd1 vssd1 vccd1 vccd1 _16669_/A sky130_fd_sc_hd__or2_1
XFILLER_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18402_ _17356_/X _18568_/A _18401_/X _17688_/A _18572_/A vssd1 vssd1 vccd1 vccd1
+ _18402_/X sky130_fd_sc_hd__a221o_1
XFILLER_250_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12826_ _12953_/A _21300_/A _25473_/Q _21320_/A vssd1 vssd1 vccd1 vccd1 _12826_/X
+ sky130_fd_sc_hd__or4bb_1
X_15614_ _20120_/A vssd1 vssd1 vccd1 vccd1 _15614_/Y sky130_fd_sc_hd__inv_2
XFILLER_250_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19382_ _19414_/B _19382_/B vssd1 vssd1 vccd1 vccd1 _19382_/X sky130_fd_sc_hd__or2_2
XFILLER_15_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16594_ _16594_/A _16788_/A vssd1 vssd1 vccd1 vccd1 _16597_/A sky130_fd_sc_hd__nand2_1
XFILLER_222_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18333_ _18027_/X _18288_/Y _18332_/X _19087_/A vssd1 vssd1 vccd1 vccd1 _18334_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15545_ _26505_/Q _26377_/Q _15557_/S vssd1 vssd1 vccd1 vccd1 _15545_/X sky130_fd_sc_hd__mux2_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _12757_/A vssd1 vssd1 vccd1 vccd1 _12758_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15476_ _26082_/Q _15453_/A _13135_/A _15475_/X vssd1 vssd1 vccd1 vccd1 _15476_/X
+ sky130_fd_sc_hd__o211a_1
X_18264_ _18070_/X _18066_/X _18265_/S vssd1 vssd1 vccd1 vccd1 _18264_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12688_ _13641_/A vssd1 vssd1 vccd1 vccd1 _12808_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_187_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14427_ _14254_/S _14425_/X _14426_/X _14100_/A _14440_/S vssd1 vssd1 vccd1 vccd1
+ _14427_/X sky130_fd_sc_hd__o311a_1
X_17215_ _25497_/Q _17529_/A _17146_/A _17443_/A vssd1 vssd1 vccd1 vccd1 _17216_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18195_ _18314_/A vssd1 vssd1 vccd1 vccd1 _18269_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14358_ _25579_/Q _14358_/B _17133_/A vssd1 vssd1 vccd1 vccd1 _14359_/D sky130_fd_sc_hd__or3_1
X_17146_ _17146_/A vssd1 vssd1 vccd1 vccd1 _17146_/X sky130_fd_sc_hd__buf_2
XFILLER_190_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13309_ _13309_/A _13309_/B vssd1 vssd1 vccd1 vccd1 _13310_/A sky130_fd_sc_hd__nor2_1
XFILLER_183_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17077_ _22361_/B _22393_/A _22361_/A vssd1 vssd1 vccd1 vccd1 _22390_/B sky130_fd_sc_hd__and3b_2
X_14289_ _26623_/Q _26719_/Q _14289_/S vssd1 vssd1 vccd1 vccd1 _14289_/X sky130_fd_sc_hd__mux2_1
XFILLER_226_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16028_ _16016_/X _16019_/X _16027_/Y vssd1 vssd1 vccd1 vccd1 _16028_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_226_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17979_ _18001_/B vssd1 vssd1 vccd1 vccd1 _17979_/Y sky130_fd_sc_hd__inv_2
XFILLER_285_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19718_ _20186_/A vssd1 vssd1 vccd1 vccd1 _19718_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_238_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20990_ _21709_/A _20990_/B vssd1 vssd1 vccd1 vccd1 _25868_/D sky130_fd_sc_hd__nor2_1
XFILLER_238_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19649_ _19649_/A _19686_/A vssd1 vssd1 vccd1 vccd1 _19649_/Y sky130_fd_sc_hd__nand2_1
XFILLER_226_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22660_ _22743_/S vssd1 vssd1 vccd1 vccd1 _22673_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_213_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21611_ _21586_/X _19373_/X _21587_/X _25825_/Q _21547_/X vssd1 vssd1 vccd1 vccd1
+ _21611_/X sky130_fd_sc_hd__a221o_1
XFILLER_244_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22591_ _26312_/Q _22591_/B vssd1 vssd1 vccd1 vccd1 _22591_/Y sky130_fd_sc_hd__nand2_1
XFILLER_222_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24330_ _27001_/Q _24331_/C _24329_/Y vssd1 vssd1 vccd1 vccd1 _27001_/D sky130_fd_sc_hd__o21a_1
X_21542_ _21538_/Y _21541_/X _21492_/X vssd1 vssd1 vccd1 vccd1 _21542_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_178_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24261_ _24269_/A _24266_/C vssd1 vssd1 vccd1 vccd1 _24261_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21473_ _21603_/A vssd1 vssd1 vccd1 vccd1 _21473_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26000_ _26592_/CLK _26000_/D vssd1 vssd1 vccd1 vccd1 _26000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23212_ _23268_/A vssd1 vssd1 vccd1 vccd1 _23281_/S sky130_fd_sc_hd__buf_4
X_20424_ _20328_/X _19415_/Y _18019_/X _14931_/Y vssd1 vssd1 vccd1 vccd1 _20424_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_107_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24192_ _24216_/A _24197_/C vssd1 vssd1 vccd1 vccd1 _24192_/Y sky130_fd_sc_hd__nor2_1
XFILLER_162_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23143_ _23143_/A vssd1 vssd1 vccd1 vccd1 _26520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20355_ _20355_/A vssd1 vssd1 vccd1 vccd1 _20355_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23074_ _26499_/Q _23073_/X _23083_/S vssd1 vssd1 vccd1 vccd1 _23075_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20286_ _25683_/Q _25682_/Q _20286_/C vssd1 vssd1 vccd1 vccd1 _20334_/C sky130_fd_sc_hd__and3_1
XFILLER_115_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26902_ _27322_/CLK _26902_/D vssd1 vssd1 vccd1 vccd1 _26902_/Q sky130_fd_sc_hd__dfxtp_1
X_22025_ _26124_/Q _20961_/X _22027_/S vssd1 vssd1 vccd1 vccd1 _22026_/A sky130_fd_sc_hd__mux2_1
XTAP_5504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26833_ _27252_/CLK _26833_/D vssd1 vssd1 vccd1 vccd1 _26833_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26764_ _27314_/CLK _26764_/D vssd1 vssd1 vccd1 vccd1 _26764_/Q sky130_fd_sc_hd__dfxtp_1
X_23976_ _26863_/Q _23571_/X _23976_/S vssd1 vssd1 vccd1 vccd1 _23977_/A sky130_fd_sc_hd__mux2_1
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22927_ _22927_/A vssd1 vssd1 vccd1 vccd1 _26439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25715_ _27329_/A _25715_/D vssd1 vssd1 vccd1 vccd1 _25715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26695_ _26797_/CLK _26695_/D vssd1 vssd1 vccd1 vccd1 _26695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13660_ _13644_/X _13655_/X _13659_/X _13821_/A vssd1 vssd1 vccd1 vccd1 _13660_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25646_ _25661_/CLK _25646_/D vssd1 vssd1 vccd1 vccd1 _25646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22858_ _26409_/Q _22698_/X _22862_/S vssd1 vssd1 vccd1 vccd1 _22859_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21809_ _21809_/A vssd1 vssd1 vccd1 vccd1 _26034_/D sky130_fd_sc_hd__clkbuf_1
X_13591_ _14173_/B vssd1 vssd1 vccd1 vccd1 _15808_/B sky130_fd_sc_hd__clkbuf_4
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25577_ _26683_/CLK _25577_/D vssd1 vssd1 vccd1 vccd1 _25577_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22789_ _26379_/Q _22704_/X _22789_/S vssd1 vssd1 vccd1 vccd1 _22790_/A sky130_fd_sc_hd__mux2_1
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _26510_/Q _26382_/Q _16086_/S vssd1 vssd1 vccd1 vccd1 _15330_/X sky130_fd_sc_hd__mux2_1
XFILLER_197_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24528_ _24538_/A _24625_/A vssd1 vssd1 vccd1 vccd1 _24528_/Y sky130_fd_sc_hd__nand2_1
X_27316_ _27316_/CLK _27316_/D vssd1 vssd1 vccd1 vccd1 _27316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15261_ _26350_/Q _26610_/Q _15276_/S vssd1 vssd1 vccd1 vccd1 _15261_/X sky130_fd_sc_hd__mux2_1
X_24459_ _24454_/X _25614_/Q _24458_/X vssd1 vssd1 vccd1 vccd1 _24948_/A sky130_fd_sc_hd__o21ai_4
XFILLER_157_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27247_ _27311_/CLK _27247_/D vssd1 vssd1 vccd1 vccd1 _27247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14212_ _14474_/S vssd1 vssd1 vccd1 vccd1 _14539_/S sky130_fd_sc_hd__buf_2
XFILLER_177_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17000_ _22491_/A _16996_/X _16990_/A _16735_/X vssd1 vssd1 vccd1 vccd1 _17000_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_177_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15192_ _15290_/A _15192_/B vssd1 vssd1 vccd1 vccd1 _15192_/X sky130_fd_sc_hd__or2_1
X_27178_ _27198_/CLK _27178_/D vssd1 vssd1 vccd1 vccd1 _27178_/Q sky130_fd_sc_hd__dfxtp_1
X_26129_ _26240_/CLK _26129_/D vssd1 vssd1 vccd1 vccd1 _26129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14143_ _13911_/X _14489_/A _14142_/X _12916_/X _25906_/Q vssd1 vssd1 vccd1 vccd1
+ _14144_/B sky130_fd_sc_hd__o32a_1
XFILLER_152_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14074_ _13250_/A _26101_/Q _26002_/Q _13657_/A _12731_/A vssd1 vssd1 vccd1 vccd1
+ _14074_/X sky130_fd_sc_hd__a221o_1
XFILLER_180_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18951_ _27117_/Q _19056_/A _18949_/X _18950_/X vssd1 vssd1 vccd1 vccd1 _18951_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_180_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13025_ _13025_/A vssd1 vssd1 vccd1 vccd1 _13026_/A sky130_fd_sc_hd__buf_2
XFILLER_140_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17902_ _15701_/B _15788_/B _17950_/S vssd1 vssd1 vccd1 vccd1 _17902_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18882_ _18552_/X _18865_/Y _18881_/X _18779_/X vssd1 vssd1 vccd1 vccd1 _18882_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_239_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17833_ _18906_/A _17833_/B vssd1 vssd1 vccd1 vccd1 _17833_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17764_ _18436_/A _17724_/X _17763_/X vssd1 vssd1 vccd1 vccd1 _17764_/X sky130_fd_sc_hd__a21o_4
XFILLER_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14976_ _14958_/X _14975_/X _14593_/X vssd1 vssd1 vccd1 vccd1 _14976_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_270_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19503_ _19499_/X _18404_/X _19501_/X _19502_/X vssd1 vssd1 vccd1 vccd1 _25635_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_63_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27276_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_235_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16715_ _22478_/A _16703_/X _16705_/X _18329_/A vssd1 vssd1 vccd1 vccd1 _16715_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_263_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13927_ _17592_/B _13927_/B vssd1 vssd1 vccd1 vccd1 _13928_/B sky130_fd_sc_hd__nor2_2
X_17695_ _17708_/A _19828_/A _17694_/Y vssd1 vssd1 vccd1 vccd1 _17736_/A sky130_fd_sc_hd__a21o_1
XFILLER_228_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_401 _17038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_412 _17048_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19434_ _27131_/Q _18748_/X _19432_/X _19433_/X vssd1 vssd1 vccd1 vccd1 _19434_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_207_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_423 _12781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16646_ _25796_/Q _17533_/A vssd1 vssd1 vccd1 vccd1 _17597_/A sky130_fd_sc_hd__nand2_2
XFILLER_250_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13858_ _13135_/A _13854_/X _13856_/X _13857_/X vssd1 vssd1 vccd1 vccd1 _13858_/X
+ sky130_fd_sc_hd__a211o_1
XINSDIODE2_434 _25726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_445 _25732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_456 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_467 _20628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12809_ _25569_/Q _17504_/C _17992_/B vssd1 vssd1 vccd1 vccd1 _12810_/D sky130_fd_sc_hd__or3b_1
X_19365_ _27097_/Q _18815_/X _18816_/X _27195_/Q _18817_/X vssd1 vssd1 vccd1 vccd1
+ _19365_/X sky130_fd_sc_hd__a221o_1
XFILLER_188_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_478 _16419_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16577_ _16594_/A vssd1 vssd1 vccd1 vccd1 _16833_/A sky130_fd_sc_hd__buf_2
XINSDIODE2_489 _16028_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13789_ _13472_/X _26884_/Q _26756_/Q _15496_/S _13494_/X vssd1 vssd1 vccd1 vccd1
+ _13789_/X sky130_fd_sc_hd__a221o_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18316_ _17959_/X _17905_/X _18318_/S vssd1 vssd1 vccd1 vccd1 _18729_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15528_ _17840_/A _15528_/B vssd1 vssd1 vccd1 vccd1 _15529_/A sky130_fd_sc_hd__nor2_1
X_19296_ _18936_/A _18352_/B _18365_/Y _18597_/X _19295_/X vssd1 vssd1 vccd1 vccd1
+ _19296_/X sky130_fd_sc_hd__o221a_1
XFILLER_188_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18247_ _19700_/A _15441_/X _18577_/A vssd1 vssd1 vccd1 vccd1 _18247_/X sky130_fd_sc_hd__mux2_1
X_15459_ _26114_/Q _26015_/Q _15459_/S vssd1 vssd1 vccd1 vccd1 _15459_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18178_ _19665_/A _16521_/A _18303_/S vssd1 vssd1 vccd1 vccd1 _18178_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17129_ _17129_/A _17131_/B vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__nand2_2
XFILLER_128_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20140_ _15441_/X _18016_/A _19589_/A _20092_/B _20125_/B vssd1 vssd1 vccd1 vccd1
+ _20144_/A sky130_fd_sc_hd__o221a_1
XFILLER_144_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20071_ _20046_/X _20049_/Y _20069_/Y _20070_/X vssd1 vssd1 vccd1 vccd1 _20071_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_98_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23830_ _23744_/X _26798_/Q _23832_/S vssd1 vssd1 vccd1 vccd1 _23831_/A sky130_fd_sc_hd__mux2_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23761_ _23760_/X _26771_/Q _23764_/S vssd1 vssd1 vccd1 vccd1 _23762_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20973_ _20973_/A _20973_/B vssd1 vssd1 vccd1 vccd1 _20974_/A sky130_fd_sc_hd__nand2_1
XFILLER_199_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25500_ _25598_/CLK _25500_/D vssd1 vssd1 vccd1 vccd1 _25500_/Q sky130_fd_sc_hd__dfxtp_1
X_22712_ _26349_/Q _22711_/X _22721_/S vssd1 vssd1 vccd1 vccd1 _22713_/A sky130_fd_sc_hd__mux2_1
X_26480_ _27287_/CLK _26480_/D vssd1 vssd1 vccd1 vccd1 _26480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23692_ _23692_/A vssd1 vssd1 vccd1 vccd1 _26749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25431_ _23738_/X _27311_/Q _25437_/S vssd1 vssd1 vccd1 vccd1 _25432_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22643_ _22724_/A vssd1 vssd1 vccd1 vccd1 _22743_/S sky130_fd_sc_hd__buf_8
XFILLER_80_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25362_ _25362_/A vssd1 vssd1 vccd1 vccd1 _27280_/D sky130_fd_sc_hd__clkbuf_1
X_22574_ _22600_/A vssd1 vssd1 vccd1 vccd1 _22574_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_278_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24313_ _26995_/Q _24311_/B _24312_/Y vssd1 vssd1 vccd1 vccd1 _26995_/D sky130_fd_sc_hd__o21a_1
X_27101_ _27173_/CLK _27101_/D vssd1 vssd1 vccd1 vccd1 _27101_/Q sky130_fd_sc_hd__dfxtp_1
X_21525_ _20679_/A _21481_/X _21459_/A _21524_/X vssd1 vssd1 vccd1 vccd1 _21525_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_194_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25293_ _23747_/X _27250_/Q _25293_/S vssd1 vssd1 vccd1 vccd1 _25294_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27032_ _27154_/CLK _27032_/D vssd1 vssd1 vccd1 vccd1 _27032_/Q sky130_fd_sc_hd__dfxtp_1
X_24244_ _24269_/A _24250_/C vssd1 vssd1 vccd1 vccd1 _24244_/Y sky130_fd_sc_hd__nor2_1
XFILLER_193_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21456_ _21284_/A _18958_/X _21286_/A _25813_/Q _21346_/X vssd1 vssd1 vccd1 vccd1
+ _21456_/X sky130_fd_sc_hd__a221o_1
XFILLER_108_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20407_ _20443_/B _20443_/C vssd1 vssd1 vccd1 vccd1 _20407_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_107_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24175_ _26949_/Q _26948_/Q _24175_/C vssd1 vssd1 vccd1 vccd1 _24176_/B sky130_fd_sc_hd__and3_1
XFILLER_108_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21387_ _21354_/X _21355_/X _21385_/Y _21386_/X vssd1 vssd1 vccd1 vccd1 _21387_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_162_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23126_ _23126_/A vssd1 vssd1 vccd1 vccd1 _26515_/D sky130_fd_sc_hd__clkbuf_1
X_20338_ _27126_/Q _20248_/X _20276_/X _20337_/Y vssd1 vssd1 vccd1 vccd1 _20338_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23057_ _23530_/A vssd1 vssd1 vccd1 vccd1 _23057_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20269_ _27155_/Q _27089_/Q vssd1 vssd1 vccd1 vccd1 _20269_/Y sky130_fd_sc_hd__nor2_1
XTAP_5312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput101 dout0[62] vssd1 vssd1 vccd1 vccd1 input101/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput112 dout1[14] vssd1 vssd1 vccd1 vccd1 input112/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22008_ _26116_/Q _20935_/X _22016_/S vssd1 vssd1 vccd1 vccd1 _22009_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput123 dout1[24] vssd1 vssd1 vccd1 vccd1 input123/X sky130_fd_sc_hd__clkbuf_1
XTAP_5345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput134 dout1[34] vssd1 vssd1 vccd1 vccd1 input134/X sky130_fd_sc_hd__clkbuf_2
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput145 dout1[44] vssd1 vssd1 vccd1 vccd1 input145/X sky130_fd_sc_hd__clkbuf_2
XTAP_5356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput156 dout1[54] vssd1 vssd1 vccd1 vccd1 input156/X sky130_fd_sc_hd__clkbuf_2
XFILLER_237_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput167 dout1[6] vssd1 vssd1 vccd1 vccd1 input167/X sky130_fd_sc_hd__clkbuf_1
X_26816_ _27299_/CLK _26816_/D vssd1 vssd1 vccd1 vccd1 _26816_/Q sky130_fd_sc_hd__dfxtp_1
X_14830_ _14831_/A _17779_/A vssd1 vssd1 vccd1 vccd1 _19427_/S sky130_fd_sc_hd__nor2_2
XFILLER_263_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput178 irq[1] vssd1 vssd1 vccd1 vccd1 input178/X sky130_fd_sc_hd__buf_6
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 jtag_tms vssd1 vssd1 vccd1 vccd1 _22390_/A sky130_fd_sc_hd__buf_12
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26747_ _26904_/CLK _26747_/D vssd1 vssd1 vccd1 vccd1 _26747_/Q sky130_fd_sc_hd__dfxtp_1
X_14761_ _16524_/A _14740_/X _14756_/X _14760_/X vssd1 vssd1 vccd1 vccd1 _14776_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23959_ _26855_/Q _23546_/X _23965_/S vssd1 vssd1 vccd1 vccd1 _23960_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16500_ _27294_/Q _26487_/Q _16500_/S vssd1 vssd1 vccd1 vccd1 _16500_/X sky130_fd_sc_hd__mux2_1
XFILLER_232_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _16071_/S _13709_/X _13710_/X _13031_/A _15646_/A vssd1 vssd1 vccd1 vccd1
+ _13717_/B sky130_fd_sc_hd__o2111a_1
XFILLER_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17480_ _26257_/Q _17458_/B _17459_/A _25985_/Q vssd1 vssd1 vccd1 vccd1 _21212_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_189_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14692_ _26126_/Q _26027_/Q _14692_/S vssd1 vssd1 vccd1 vccd1 _14692_/X sky130_fd_sc_hd__mux2_1
XFILLER_232_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26678_ _27321_/CLK _26678_/D vssd1 vssd1 vccd1 vccd1 _26678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16431_ _14793_/A _16427_/X _16430_/X _14808_/A vssd1 vssd1 vccd1 vccd1 _16431_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13643_ _25878_/Q _16419_/B vssd1 vssd1 vccd1 vccd1 _13643_/X sky130_fd_sc_hd__or2_1
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25629_ _27327_/CLK _25629_/D vssd1 vssd1 vccd1 vccd1 _25629_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_32_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19150_ _19448_/A _19121_/Y _19149_/X vssd1 vssd1 vccd1 vccd1 _19150_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_158_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13574_ _25911_/Q _12902_/A _15874_/A _13573_/Y vssd1 vssd1 vccd1 vccd1 _13574_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16362_ _15111_/A _26613_/Q _16441_/S _26353_/Q _16278_/S vssd1 vssd1 vccd1 vccd1
+ _16362_/X sky130_fd_sc_hd__o221a_1
XFILLER_9_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18101_ _18443_/A vssd1 vssd1 vccd1 vccd1 _18559_/A sky130_fd_sc_hd__clkbuf_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15313_ _15313_/A vssd1 vssd1 vccd1 vccd1 _15313_/X sky130_fd_sc_hd__clkbuf_2
X_16293_ _25655_/Q _14609_/A _15135_/X vssd1 vssd1 vccd1 vccd1 _16293_/X sky130_fd_sc_hd__a21o_1
X_19081_ _25743_/Q _19081_/B vssd1 vssd1 vccd1 vccd1 _19082_/B sky130_fd_sc_hd__nor2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_181_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26904_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_185_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18032_ _18227_/C _18032_/B vssd1 vssd1 vccd1 vccd1 _18032_/Y sky130_fd_sc_hd__nand2_1
XFILLER_258_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15244_ _15244_/A vssd1 vssd1 vccd1 vccd1 _15244_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_110_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27004_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_166_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15175_ _15384_/S vssd1 vssd1 vccd1 vccd1 _16397_/S sky130_fd_sc_hd__buf_4
XFILLER_153_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14126_ _17801_/B _14127_/B vssd1 vssd1 vccd1 vccd1 _18372_/S sky130_fd_sc_hd__and2_1
XFILLER_181_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_9_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_153_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19983_ _20080_/A _19984_/B vssd1 vssd1 vccd1 vccd1 _19983_/X sky130_fd_sc_hd__and2_1
X_14057_ _14043_/X _14055_/X _14056_/X _13277_/A vssd1 vssd1 vccd1 vccd1 _14057_/X
+ sky130_fd_sc_hd__a211o_1
X_18934_ _13641_/B _18890_/X _18931_/Y _18932_/X _18933_/X vssd1 vssd1 vccd1 vccd1
+ _18934_/X sky130_fd_sc_hd__a221o_4
XFILLER_279_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13008_ _13008_/A vssd1 vssd1 vccd1 vccd1 _13009_/A sky130_fd_sc_hd__buf_2
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18865_ _18852_/Y _18856_/X _18864_/X vssd1 vssd1 vccd1 vccd1 _18865_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_239_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17816_ _18906_/A _17816_/B _17816_/C _18726_/A vssd1 vssd1 vccd1 vccd1 _17816_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_227_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18796_ _18795_/Y _16635_/C _19453_/S vssd1 vssd1 vccd1 vccd1 _18796_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17747_ _17762_/A _17747_/B _17747_/C _17722_/B vssd1 vssd1 vccd1 vccd1 _17749_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_282_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14959_ _27323_/Q _26580_/Q _14963_/S vssd1 vssd1 vccd1 vccd1 _14959_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17678_ _17738_/A vssd1 vssd1 vccd1 vccd1 _21203_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_220 _20055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_231 _20168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19417_ _18144_/A _19388_/A _19416_/X vssd1 vssd1 vccd1 vccd1 _19417_/Y sky130_fd_sc_hd__o21ai_1
XINSDIODE2_242 _21070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16629_ _17816_/B vssd1 vssd1 vccd1 vccd1 _18855_/A sky130_fd_sc_hd__buf_4
XINSDIODE2_253 _16829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_264 _20686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_275 _25487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_286 _25818_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_297 _25801_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19348_ _19381_/B _19348_/B vssd1 vssd1 vccd1 vccd1 _19348_/X sky130_fd_sc_hd__or2_2
XFILLER_176_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19279_ _19274_/X _19275_/X _19278_/X _18792_/X vssd1 vssd1 vccd1 vccd1 _19279_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
X_21310_ _21573_/A vssd1 vssd1 vccd1 vccd1 _21310_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22290_ _26208_/Q _22279_/X _22285_/X _26309_/Q _22286_/X vssd1 vssd1 vccd1 vccd1
+ _22290_/X sky130_fd_sc_hd__a221o_1
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21241_ _25027_/A vssd1 vssd1 vccd1 vccd1 _24871_/A sky130_fd_sc_hd__buf_6
XFILLER_191_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21172_ _21172_/A _21172_/B vssd1 vssd1 vccd1 vccd1 _21173_/A sky130_fd_sc_hd__or2_1
XFILLER_116_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20123_ _20115_/A _20121_/X _19698_/X _20668_/A vssd1 vssd1 vccd1 vccd1 _20125_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_259_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25980_ _27022_/CLK _25980_/D vssd1 vssd1 vccd1 vccd1 _25980_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_86_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24931_ _24954_/A vssd1 vssd1 vccd1 vccd1 _24951_/B sky130_fd_sc_hd__clkbuf_2
X_20054_ _22500_/A _19876_/X _20045_/X _20053_/Y _19874_/X vssd1 vssd1 vccd1 vccd1
+ _25674_/D sky130_fd_sc_hd__o221a_1
XFILLER_98_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24862_ _24860_/Y _24861_/X _24854_/X vssd1 vssd1 vccd1 vccd1 _27121_/D sky130_fd_sc_hd__a21oi_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26601_ _26601_/CLK _26601_/D vssd1 vssd1 vccd1 vccd1 _26601_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23813_ _23718_/X _26790_/Q _23821_/S vssd1 vssd1 vccd1 vccd1 _23814_/A sky130_fd_sc_hd__mux2_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24793_ _24788_/Y _24792_/X _22634_/X vssd1 vssd1 vccd1 vccd1 _27103_/D sky130_fd_sc_hd__a21oi_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26532_ _27276_/CLK _26532_/D vssd1 vssd1 vccd1 vccd1 _26532_/Q sky130_fd_sc_hd__dfxtp_1
X_23744_ _23744_/A vssd1 vssd1 vccd1 vccd1 _23744_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20956_ _25855_/Q _20955_/X _20965_/S vssd1 vssd1 vccd1 vccd1 _20957_/A sky130_fd_sc_hd__mux2_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26463_ _26465_/CLK _26463_/D vssd1 vssd1 vccd1 vccd1 _26463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23675_ _23675_/A vssd1 vssd1 vccd1 vccd1 _26743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20887_ _23702_/A vssd1 vssd1 vccd1 vccd1 _20887_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22626_ _26327_/Q vssd1 vssd1 vccd1 vccd1 _22629_/A sky130_fd_sc_hd__inv_2
X_25414_ _25414_/A vssd1 vssd1 vccd1 vccd1 _27303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26394_ _27264_/CLK _26394_/D vssd1 vssd1 vccd1 vccd1 _26394_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_201_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25345_ _25391_/S vssd1 vssd1 vccd1 vccd1 _25354_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_139_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22557_ _22553_/X _22556_/Y _22547_/X vssd1 vssd1 vccd1 vccd1 _26298_/D sky130_fd_sc_hd__a21oi_1
XFILLER_194_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21508_ _25488_/Q _21574_/B vssd1 vssd1 vccd1 vccd1 _21508_/X sky130_fd_sc_hd__or2_1
X_13290_ _13321_/A _13290_/B vssd1 vssd1 vccd1 vccd1 _13290_/X sky130_fd_sc_hd__or2_1
X_25276_ _23722_/X _27242_/Q _25282_/S vssd1 vssd1 vccd1 vccd1 _25277_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22488_ _22488_/A vssd1 vssd1 vccd1 vccd1 _26269_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24227_ _26966_/Q _26965_/Q _24227_/C vssd1 vssd1 vccd1 vccd1 _24233_/C sky130_fd_sc_hd__and3_1
X_27015_ _27049_/CLK _27015_/D vssd1 vssd1 vccd1 vccd1 _27015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21439_ _21439_/A vssd1 vssd1 vccd1 vccd1 _21439_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24158_ _26943_/Q _24160_/C _17137_/A vssd1 vssd1 vccd1 vccd1 _24159_/B sky130_fd_sc_hd__o21ai_1
XFILLER_135_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23109_ _26510_/Q _23108_/X _23115_/S vssd1 vssd1 vccd1 vccd1 _23110_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24089_ _24146_/S vssd1 vssd1 vccd1 vccd1 _24098_/S sky130_fd_sc_hd__buf_2
X_16980_ _16980_/A _16980_/B _16980_/C vssd1 vssd1 vccd1 vccd1 _16981_/A sky130_fd_sc_hd__and3_2
XFILLER_111_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15931_ _26633_/Q _26729_/Q _15931_/S vssd1 vssd1 vccd1 vccd1 _15932_/B sky130_fd_sc_hd__mux2_1
XFILLER_89_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18650_ _25734_/Q _18650_/B vssd1 vssd1 vccd1 vccd1 _18651_/B sky130_fd_sc_hd__nor2_1
XTAP_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15862_ _15589_/A _26858_/Q _25772_/Q _15582_/A _15859_/A vssd1 vssd1 vccd1 vccd1
+ _15862_/X sky130_fd_sc_hd__a221o_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17601_ _17560_/X _17623_/B _13565_/X _17554_/X _25919_/Q vssd1 vssd1 vccd1 vccd1
+ _17601_/Y sky130_fd_sc_hd__o32ai_1
XFILLER_97_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14813_ _26518_/Q _26390_/Q _14813_/S vssd1 vssd1 vccd1 vccd1 _14813_/X sky130_fd_sc_hd__mux2_1
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ _18382_/X _18580_/Y _18010_/C vssd1 vssd1 vccd1 vccd1 _18581_/X sky130_fd_sc_hd__o21a_1
XFILLER_236_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _25644_/Q _15443_/B _14612_/A vssd1 vssd1 vccd1 vccd1 _15793_/X sky130_fd_sc_hd__a21o_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17532_ _17548_/A _17532_/B vssd1 vssd1 vccd1 vccd1 _25567_/D sky130_fd_sc_hd__nor2_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14744_ _14744_/A vssd1 vssd1 vccd1 vccd1 _14890_/A sky130_fd_sc_hd__buf_2
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_opt_4_0_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25824_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_44_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17463_ _26254_/Q _17454_/A _17460_/A _25982_/Q vssd1 vssd1 vccd1 vccd1 _17465_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_232_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14675_ _26094_/Q _14652_/S _14700_/S _14674_/X vssd1 vssd1 vccd1 vccd1 _14675_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19202_ _27028_/Q _19063_/X _19201_/X _18565_/X vssd1 vssd1 vccd1 vccd1 _19202_/X
+ sky130_fd_sc_hd__a22o_1
X_16414_ _14593_/A _16408_/X _16413_/X vssd1 vssd1 vccd1 vccd1 _16414_/Y sky130_fd_sc_hd__o21ai_4
X_13626_ _13884_/S vssd1 vssd1 vccd1 vccd1 _15818_/S sky130_fd_sc_hd__clkbuf_4
X_17394_ _25549_/Q _17392_/B _17393_/Y vssd1 vssd1 vccd1 vccd1 _25549_/D sky130_fd_sc_hd__o21a_1
XFILLER_220_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19133_ _27154_/Q _19334_/B vssd1 vssd1 vccd1 vccd1 _19133_/X sky130_fd_sc_hd__or2_1
XFILLER_158_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16345_ _16336_/X _16343_/X _16344_/X vssd1 vssd1 vccd1 vccd1 _16345_/X sky130_fd_sc_hd__o21a_1
X_13557_ _13557_/A vssd1 vssd1 vccd1 vccd1 _13558_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19064_ _27152_/Q _19334_/B vssd1 vssd1 vccd1 vccd1 _19064_/X sky130_fd_sc_hd__or2_1
X_13488_ _13488_/A vssd1 vssd1 vccd1 vccd1 _15109_/A sky130_fd_sc_hd__buf_4
X_16276_ _26803_/Q _26447_/Q _16277_/S vssd1 vssd1 vccd1 vccd1 _16276_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18015_ _19914_/A vssd1 vssd1 vccd1 vccd1 _18016_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15227_ _15225_/X _15226_/X _15227_/S vssd1 vssd1 vccd1 vccd1 _15227_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput405 _17014_/X vssd1 vssd1 vccd1 vccd1 din0[7] sky130_fd_sc_hd__buf_2
Xoutput416 _25951_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[15] sky130_fd_sc_hd__buf_2
XFILLER_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput427 _25961_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[25] sky130_fd_sc_hd__buf_2
Xoutput438 _25942_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[6] sky130_fd_sc_hd__buf_2
X_15158_ _15351_/B vssd1 vssd1 vccd1 vccd1 _16402_/S sky130_fd_sc_hd__buf_2
XFILLER_5_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput449 _26236_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[4] sky130_fd_sc_hd__buf_2
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14109_ _26593_/Q _14109_/B vssd1 vssd1 vccd1 vccd1 _14109_/X sky130_fd_sc_hd__or2_1
XFILLER_271_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15089_ _14890_/A _26614_/Q _14891_/A _26354_/Q _15095_/S vssd1 vssd1 vccd1 vccd1
+ _15089_/X sky130_fd_sc_hd__o221a_1
X_19966_ _22494_/A _19638_/X _19964_/X _19965_/X vssd1 vssd1 vccd1 vccd1 _25671_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_234_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18917_ _27148_/Q _18952_/B vssd1 vssd1 vccd1 vccd1 _18917_/X sky130_fd_sc_hd__or2_1
XFILLER_86_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19897_ _27141_/Q _27075_/Q vssd1 vssd1 vccd1 vccd1 _19897_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18848_ _19042_/A _18848_/B vssd1 vssd1 vccd1 vccd1 _18848_/Y sky130_fd_sc_hd__nand2_1
XFILLER_267_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18779_ _18927_/A vssd1 vssd1 vccd1 vccd1 _18779_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_283_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20810_ _25801_/Q vssd1 vssd1 vccd1 vccd1 _20811_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_209_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21790_ _21790_/A vssd1 vssd1 vccd1 vccd1 _26027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20741_ _20787_/S vssd1 vssd1 vccd1 vccd1 _20750_/S sky130_fd_sc_hd__buf_2
XFILLER_51_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23460_ _23506_/S vssd1 vssd1 vccd1 vccd1 _23469_/S sky130_fd_sc_hd__buf_6
XFILLER_23_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20672_ _26279_/Q _20660_/X _20670_/X _20671_/X vssd1 vssd1 vccd1 vccd1 _25742_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22411_ _22405_/A _22395_/Y _22406_/X _22410_/X vssd1 vssd1 vccd1 vccd1 _22411_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_149_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23391_ _26631_/Q _23073_/X _23397_/S vssd1 vssd1 vccd1 vccd1 _23392_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25130_ _20683_/A _25113_/X _25129_/X vssd1 vssd1 vccd1 vccd1 _25130_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_109_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22342_ _22335_/Y _22340_/X _22341_/X _22330_/X vssd1 vssd1 vccd1 vccd1 _26226_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25061_ _22491_/A _25038_/X _25060_/X _16735_/X _25052_/X vssd1 vssd1 vccd1 vccd1
+ _25061_/X sky130_fd_sc_hd__a221o_1
X_22273_ _22288_/A vssd1 vssd1 vccd1 vccd1 _22273_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24012_ _24012_/A vssd1 vssd1 vccd1 vccd1 _26878_/D sky130_fd_sc_hd__clkbuf_1
X_21224_ _20624_/A _21277_/A _21222_/X _21279_/A vssd1 vssd1 vccd1 vccd1 _21224_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21155_ _21155_/A vssd1 vssd1 vccd1 vccd1 _25923_/D sky130_fd_sc_hd__clkbuf_1
X_20106_ _20131_/A _20105_/Y _20069_/Y _20071_/Y vssd1 vssd1 vccd1 vccd1 _20106_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_259_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25963_ _26995_/CLK _25963_/D vssd1 vssd1 vccd1 vccd1 _25963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21086_ _21100_/A _21086_/B vssd1 vssd1 vccd1 vccd1 _21087_/A sky130_fd_sc_hd__or2_1
XFILLER_101_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24914_ _24954_/A vssd1 vssd1 vccd1 vccd1 _24923_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_19_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20037_ _20061_/A _20061_/B vssd1 vssd1 vccd1 vccd1 _20082_/A sky130_fd_sc_hd__xnor2_2
XFILLER_246_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25894_ _26677_/CLK _25894_/D vssd1 vssd1 vccd1 vccd1 _25894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24845_ _20666_/A _24829_/X _24711_/Y _24830_/X vssd1 vssd1 vccd1 vccd1 _24845_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_262_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _25591_/Q _25590_/Q _12790_/C vssd1 vssd1 vccd1 vccd1 _12790_/X sky130_fd_sc_hd__or3_1
X_21988_ _26107_/Q _20907_/X _21994_/S vssd1 vssd1 vccd1 vccd1 _21989_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24776_ _24341_/A _24900_/C _24776_/C vssd1 vssd1 vccd1 vccd1 _24777_/B sky130_fd_sc_hd__and3b_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26515_ _27322_/CLK _26515_/D vssd1 vssd1 vccd1 vccd1 _26515_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23727_ _23727_/A vssd1 vssd1 vccd1 vccd1 _26760_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939_ _23754_/A vssd1 vssd1 vccd1 vccd1 _20939_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14460_ _13250_/A _25759_/Q _14551_/S _26845_/Q _14047_/A vssd1 vssd1 vccd1 vccd1
+ _14460_/X sky130_fd_sc_hd__o221a_1
XFILLER_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26446_ _26611_/CLK _26446_/D vssd1 vssd1 vccd1 vccd1 _26446_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23658_ _23669_/A vssd1 vssd1 vccd1 vccd1 _23667_/S sky130_fd_sc_hd__buf_6
XFILLER_224_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13411_ _14252_/S vssd1 vssd1 vccd1 vccd1 _15807_/S sky130_fd_sc_hd__clkbuf_4
X_22609_ _22606_/X _22608_/Y _22600_/X vssd1 vssd1 vccd1 vccd1 _26318_/D sky130_fd_sc_hd__a21oi_1
X_14391_ _26654_/Q _25694_/Q _14391_/S vssd1 vssd1 vccd1 vccd1 _14391_/X sky130_fd_sc_hd__mux2_1
X_26377_ _27280_/CLK _26377_/D vssd1 vssd1 vccd1 vccd1 _26377_/Q sky130_fd_sc_hd__dfxtp_1
X_23589_ _23589_/A vssd1 vssd1 vccd1 vccd1 _26708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13342_ _14047_/A vssd1 vssd1 vccd1 vccd1 _14473_/S sky130_fd_sc_hd__clkbuf_4
X_16130_ _25651_/Q _16130_/B vssd1 vssd1 vccd1 vccd1 _16130_/X sky130_fd_sc_hd__and2_1
X_25328_ _27265_/Q _23693_/A _25332_/S vssd1 vssd1 vccd1 vccd1 _25329_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13273_ _13545_/A vssd1 vssd1 vccd1 vccd1 _13274_/A sky130_fd_sc_hd__buf_4
XFILLER_183_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16061_ _25888_/Q _16061_/B vssd1 vssd1 vccd1 vccd1 _16061_/X sky130_fd_sc_hd__or2_1
X_25259_ _25259_/A vssd1 vssd1 vccd1 vccd1 _27234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15012_ _20696_/A _19374_/A _15012_/S vssd1 vssd1 vccd1 vccd1 _17850_/A sky130_fd_sc_hd__mux2_2
XFILLER_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19820_ _19819_/Y _27139_/Q _19820_/S vssd1 vssd1 vccd1 vccd1 _19820_/X sky130_fd_sc_hd__mux2_4
XFILLER_69_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19751_ _27137_/Q _27071_/Q vssd1 vssd1 vccd1 vccd1 _19752_/B sky130_fd_sc_hd__nand2_1
XFILLER_78_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16963_ _16983_/A _16973_/B _16963_/C vssd1 vssd1 vccd1 vccd1 _16963_/X sky130_fd_sc_hd__and3_1
XFILLER_96_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18702_ _18437_/X _18691_/X _18701_/X vssd1 vssd1 vccd1 vccd1 _18702_/X sky130_fd_sc_hd__a21o_4
XFILLER_209_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15914_ _26793_/Q _26437_/Q _15914_/S vssd1 vssd1 vccd1 vccd1 _15914_/X sky130_fd_sc_hd__mux2_1
XFILLER_231_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19682_ _24777_/A vssd1 vssd1 vccd1 vccd1 _24810_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_249_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16894_ _16894_/A vssd1 vssd1 vccd1 vccd1 _16894_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_265_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18633_ _18634_/A _18634_/B _16735_/A vssd1 vssd1 vccd1 vccd1 _18635_/A sky130_fd_sc_hd__o21bai_1
XFILLER_280_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15845_ _15589_/A _26342_/Q _26602_/Q _15408_/A _15843_/A vssd1 vssd1 vccd1 vccd1
+ _15845_/X sky130_fd_sc_hd__a221o_1
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18564_ _19870_/A _19261_/B vssd1 vssd1 vccd1 vccd1 _18564_/X sky130_fd_sc_hd__or2_1
XFILLER_80_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15776_ _15776_/A _15776_/B vssd1 vssd1 vccd1 vccd1 _15776_/X sky130_fd_sc_hd__or2_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12988_ _12992_/A _13029_/A vssd1 vssd1 vccd1 vccd1 _12989_/A sky130_fd_sc_hd__nor2_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17515_ _19650_/A vssd1 vssd1 vccd1 vccd1 _19636_/A sky130_fd_sc_hd__buf_4
XFILLER_233_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14727_ _14727_/A vssd1 vssd1 vccd1 vccd1 _16195_/S sky130_fd_sc_hd__buf_6
X_18495_ _18495_/A _18495_/B vssd1 vssd1 vccd1 vccd1 _18495_/Y sky130_fd_sc_hd__nor2_1
XFILLER_220_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17446_ _26326_/Q _26325_/Q vssd1 vssd1 vccd1 vccd1 _17447_/B sky130_fd_sc_hd__nor2_1
XFILLER_221_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14658_ _25827_/Q _14652_/S _14700_/S _14657_/X vssd1 vssd1 vccd1 vccd1 _14658_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13609_ _26661_/Q _25701_/Q _15964_/S vssd1 vssd1 vccd1 vccd1 _13609_/X sky130_fd_sc_hd__mux2_1
X_17377_ _17375_/X _17379_/C _17376_/Y vssd1 vssd1 vccd1 vccd1 _25544_/D sky130_fd_sc_hd__o21a_1
X_14589_ _15290_/A vssd1 vssd1 vccd1 vccd1 _16250_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19116_ _19087_/X _19114_/X _19115_/Y _18884_/X vssd1 vssd1 vccd1 vccd1 _19117_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16328_ _16328_/A _16328_/B vssd1 vssd1 vccd1 vccd1 _16328_/Y sky130_fd_sc_hd__nand2_1
XFILLER_229_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19047_ _19034_/A _19011_/B _17840_/X vssd1 vssd1 vccd1 vccd1 _19048_/B sky130_fd_sc_hd__a21bo_1
X_16259_ _26087_/Q _25892_/Q _16259_/S vssd1 vssd1 vccd1 vccd1 _16259_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_8 _22368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19949_ _20652_/A _19771_/X _19948_/X _19604_/X vssd1 vssd1 vccd1 vccd1 _19977_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22960_ _26455_/Q _22742_/X _22960_/S vssd1 vssd1 vccd1 vccd1 _22961_/A sky130_fd_sc_hd__mux2_1
XFILLER_261_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_261_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21911_ _20529_/X _26073_/Q _21911_/S vssd1 vssd1 vccd1 vccd1 _21912_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22891_ _22947_/A vssd1 vssd1 vccd1 vccd1 _22960_/S sky130_fd_sc_hd__buf_8
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24630_ _24630_/A vssd1 vssd1 vccd1 vccd1 _25221_/A sky130_fd_sc_hd__clkbuf_2
X_21842_ _21842_/A vssd1 vssd1 vccd1 vccd1 _26049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24561_ _24561_/A vssd1 vssd1 vccd1 vccd1 _24615_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_252_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21773_ _21773_/A vssd1 vssd1 vccd1 vccd1 _26019_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_270_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26300_ _26327_/CLK _26300_/D vssd1 vssd1 vccd1 vccd1 _26300_/Q sky130_fd_sc_hd__dfxtp_1
X_20724_ _20500_/X _25760_/Q _20728_/S vssd1 vssd1 vccd1 vccd1 _20725_/A sky130_fd_sc_hd__mux2_1
X_23512_ _26684_/Q _23508_/X _23524_/S vssd1 vssd1 vccd1 vccd1 _23513_/A sky130_fd_sc_hd__mux2_1
X_24492_ _24492_/A hold1/A vssd1 vssd1 vccd1 vccd1 _24492_/Y sky130_fd_sc_hd__nand2_1
X_27280_ _27280_/CLK _27280_/D vssd1 vssd1 vccd1 vccd1 _27280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26231_ _26297_/CLK _26231_/D vssd1 vssd1 vccd1 vccd1 _26231_/Q sky130_fd_sc_hd__dfxtp_1
X_23443_ _26654_/Q _23044_/X _23447_/S vssd1 vssd1 vccd1 vccd1 _23444_/A sky130_fd_sc_hd__mux2_1
X_20655_ _26273_/Q _20646_/X _20654_/X _20644_/X vssd1 vssd1 vccd1 vccd1 _25736_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26162_ _27264_/CLK _26162_/D vssd1 vssd1 vccd1 vccd1 _26162_/Q sky130_fd_sc_hd__dfxtp_1
X_23374_ _23374_/A vssd1 vssd1 vccd1 vccd1 _26623_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20586_ _20586_/A vssd1 vssd1 vccd1 vccd1 _25714_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22325_ _26220_/Q _22154_/A _22316_/X _26321_/Q _22317_/X vssd1 vssd1 vccd1 vccd1
+ _22325_/X sky130_fd_sc_hd__a221o_1
XFILLER_192_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25113_ _25113_/A vssd1 vssd1 vccd1 vccd1 _25113_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26093_ _26905_/CLK _26093_/D vssd1 vssd1 vccd1 vccd1 _26093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25044_ _22485_/A _25038_/X _25033_/X _18483_/A _25024_/X vssd1 vssd1 vccd1 vccd1
+ _25044_/X sky130_fd_sc_hd__a221o_1
XFILLER_279_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22256_ _22271_/A vssd1 vssd1 vccd1 vccd1 _22256_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_180_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21207_ _26584_/Q _21562_/C vssd1 vssd1 vccd1 vccd1 _21866_/B sky130_fd_sc_hd__and2_1
XFILLER_132_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22187_ _22203_/A vssd1 vssd1 vccd1 vccd1 _22187_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_254_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21138_ _21138_/A vssd1 vssd1 vccd1 vccd1 _21154_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_278_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26995_ _26995_/CLK _26995_/D vssd1 vssd1 vccd1 vccd1 _26995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13960_ _14552_/S vssd1 vssd1 vccd1 vccd1 _14309_/S sky130_fd_sc_hd__clkbuf_4
X_25946_ _27022_/CLK _25946_/D vssd1 vssd1 vccd1 vccd1 _25946_/Q sky130_fd_sc_hd__dfxtp_1
X_21069_ _21138_/A vssd1 vssd1 vccd1 vccd1 _21197_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12911_ _12911_/A _12911_/B _15871_/A vssd1 vssd1 vccd1 vccd1 _12912_/A sky130_fd_sc_hd__or3_2
XFILLER_74_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25877_ _26601_/CLK _25877_/D vssd1 vssd1 vccd1 vccd1 _25877_/Q sky130_fd_sc_hd__dfxtp_4
X_13891_ _14344_/S vssd1 vssd1 vccd1 vccd1 _14433_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_19_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15630_ _15630_/A vssd1 vssd1 vccd1 vccd1 _15643_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _25795_/Q _25993_/Q vssd1 vssd1 vccd1 vccd1 _12899_/A sky130_fd_sc_hd__or2b_2
X_24828_ _27113_/Q _24837_/B vssd1 vssd1 vccd1 vccd1 _24828_/Y sky130_fd_sc_hd__nand2_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15561_ _26669_/Q _15561_/B vssd1 vssd1 vccd1 vccd1 _15561_/X sky130_fd_sc_hd__or2_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12773_/A vssd1 vssd1 vccd1 vccd1 _12774_/A sky130_fd_sc_hd__buf_2
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24759_ _20434_/B _24744_/X _25151_/A _24740_/X vssd1 vssd1 vccd1 vccd1 _24760_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_261_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17300_ _17299_/X _17303_/C _17269_/X vssd1 vssd1 vccd1 vccd1 _17300_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14264_/S _14510_/X _14511_/X vssd1 vssd1 vccd1 vccd1 _14512_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _19003_/A _18229_/X _18279_/X _18976_/A vssd1 vssd1 vccd1 vccd1 _18281_/B
+ sky130_fd_sc_hd__a22o_1
X_15492_ _15760_/A vssd1 vssd1 vccd1 vccd1 _15852_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_187_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17231_ _17242_/A _22535_/B vssd1 vssd1 vccd1 vccd1 _25501_/D sky130_fd_sc_hd__nor2_1
XFILLER_203_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26429_ _27267_/CLK _26429_/D vssd1 vssd1 vccd1 vccd1 _26429_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14443_ _14443_/A vssd1 vssd1 vccd1 vccd1 _16578_/B sky130_fd_sc_hd__inv_2
XFILLER_202_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_88_wb_clk_i _25501_/CLK vssd1 vssd1 vccd1 vccd1 _26878_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17162_ _17162_/A _17195_/B vssd1 vssd1 vccd1 vccd1 _17162_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14374_ _14372_/X _14373_/X _14390_/S vssd1 vssd1 vccd1 vccd1 _14374_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16113_ _16113_/A vssd1 vssd1 vccd1 vccd1 _16260_/S sky130_fd_sc_hd__buf_6
XFILLER_128_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13325_ _15321_/A _25840_/Q _26040_/Q _16189_/S _16088_/A vssd1 vssd1 vccd1 vccd1
+ _13325_/X sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26799_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17093_ _22230_/B vssd1 vssd1 vccd1 vccd1 _17094_/B sky130_fd_sc_hd__inv_2
XFILLER_171_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16044_ _16625_/A _16626_/B _16043_/Y _18938_/S vssd1 vssd1 vccd1 vccd1 _16614_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13256_ _13256_/A vssd1 vssd1 vccd1 vccd1 _14054_/A sky130_fd_sc_hd__buf_2
XFILLER_182_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13187_ _13256_/A vssd1 vssd1 vccd1 vccd1 _14060_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19803_ _19823_/A _19803_/B vssd1 vssd1 vccd1 vccd1 _19808_/A sky130_fd_sc_hd__xnor2_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17995_ _17995_/A _17995_/B _19455_/B vssd1 vssd1 vccd1 vccd1 _18308_/B sky130_fd_sc_hd__and3_1
XFILLER_85_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19734_ _19675_/A _19675_/B _19703_/X _19705_/B _19733_/X vssd1 vssd1 vccd1 vccd1
+ _19736_/B sky130_fd_sc_hd__o311a_1
XFILLER_78_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16946_ _16946_/A _16954_/A vssd1 vssd1 vccd1 vccd1 _16946_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19665_ _19665_/A _20055_/B vssd1 vssd1 vccd1 vccd1 _19665_/X sky130_fd_sc_hd__or2_1
XFILLER_64_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16877_ _16463_/X _23555_/A _15830_/Y _16860_/B vssd1 vssd1 vccd1 vccd1 _16877_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_65_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18616_ _19896_/A _19367_/B vssd1 vssd1 vccd1 vccd1 _18616_/X sky130_fd_sc_hd__or2_1
XFILLER_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15828_ _13031_/A _15819_/X _15827_/X _14713_/C vssd1 vssd1 vccd1 vccd1 _15828_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19596_ _19774_/B vssd1 vssd1 vccd1 vccd1 _20125_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18547_ _18496_/Y _18546_/Y _18547_/S vssd1 vssd1 vccd1 vccd1 _18547_/X sky130_fd_sc_hd__mux2_1
X_15759_ _26503_/Q _26375_/Q _15759_/S vssd1 vssd1 vccd1 vccd1 _15760_/B sky130_fd_sc_hd__mux2_1
XFILLER_52_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18478_ _13980_/X _18285_/X _18477_/X _18409_/X _25604_/Q vssd1 vssd1 vccd1 vccd1
+ _18479_/B sky130_fd_sc_hd__a32o_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17429_ _25561_/Q _17434_/C vssd1 vssd1 vccd1 vccd1 _17430_/B sky130_fd_sc_hd__and2_1
XFILLER_166_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20440_ _22531_/A _19638_/X _20439_/X _19965_/X vssd1 vssd1 vccd1 vccd1 _25689_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_277_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20371_ _27159_/Q _20370_/Y _20371_/S vssd1 vssd1 vccd1 vccd1 _20371_/X sky130_fd_sc_hd__mux2_2
XFILLER_277_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22110_ _22152_/A vssd1 vssd1 vccd1 vccd1 _22110_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23090_ _26504_/Q _23089_/X _23099_/S vssd1 vssd1 vccd1 vccd1 _23091_/A sky130_fd_sc_hd__mux2_1
XFILLER_279_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22041_ _22041_/A vssd1 vssd1 vccd1 vccd1 _26130_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25800_ _26520_/CLK _25800_/D vssd1 vssd1 vccd1 vccd1 _25800_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26780_ _27295_/CLK _26780_/D vssd1 vssd1 vccd1 vccd1 _26780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23992_ _26870_/Q _23594_/X _23998_/S vssd1 vssd1 vccd1 vccd1 _23993_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25731_ _26271_/CLK _25731_/D vssd1 vssd1 vccd1 vccd1 _25731_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22943_ _26447_/Q _22717_/X _22945_/S vssd1 vssd1 vccd1 vccd1 _22944_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25662_ _26264_/CLK _25662_/D vssd1 vssd1 vccd1 vccd1 _25662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22874_ _22874_/A vssd1 vssd1 vccd1 vccd1 _26416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24613_ _24969_/A _24621_/B vssd1 vssd1 vccd1 vccd1 _24613_/Y sky130_fd_sc_hd__nand2_1
X_21825_ _26042_/Q _20913_/X _21827_/S vssd1 vssd1 vccd1 vccd1 _21826_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25593_ _27327_/CLK _25593_/D vssd1 vssd1 vccd1 vccd1 _25593_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24544_ _25206_/D _24544_/B vssd1 vssd1 vccd1 vccd1 _24561_/A sky130_fd_sc_hd__nor2_4
XFILLER_70_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21756_ _21778_/A vssd1 vssd1 vccd1 vccd1 _21765_/S sky130_fd_sc_hd__buf_4
XPHY_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20707_ _27101_/Q _22638_/B _20707_/C _20707_/D vssd1 vssd1 vccd1 vccd1 _20707_/X
+ sky130_fd_sc_hd__and4_1
X_27263_ _27265_/CLK _27263_/D vssd1 vssd1 vccd1 vccd1 _27263_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_4_11_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_11_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
X_21687_ _21698_/A vssd1 vssd1 vccd1 vccd1 _21696_/S sky130_fd_sc_hd__clkbuf_2
X_24475_ _26312_/Q _24473_/X _24474_/X input225/X _21885_/A vssd1 vssd1 vccd1 vccd1
+ _24475_/X sky130_fd_sc_hd__a221o_2
XFILLER_11_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26214_ _26980_/CLK _26214_/D vssd1 vssd1 vccd1 vccd1 _26214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23426_ _26647_/Q _23124_/X _23430_/S vssd1 vssd1 vccd1 vccd1 _23427_/A sky130_fd_sc_hd__mux2_1
X_20638_ _26266_/Q _20633_/X _20637_/X _20631_/X vssd1 vssd1 vccd1 vccd1 _25729_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27194_ _27196_/CLK _27194_/D vssd1 vssd1 vccd1 vccd1 _27194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26145_ _27280_/CLK _26145_/D vssd1 vssd1 vccd1 vccd1 _26145_/Q sky130_fd_sc_hd__dfxtp_1
X_23357_ _20613_/X _26617_/Q _23357_/S vssd1 vssd1 vccd1 vccd1 _23358_/A sky130_fd_sc_hd__mux2_1
X_20569_ _20569_/A vssd1 vssd1 vccd1 vccd1 _25710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22308_ _26214_/Q _22294_/X _22300_/X _26315_/Q _22301_/X vssd1 vssd1 vccd1 vccd1
+ _22308_/X sky130_fd_sc_hd__a221o_1
X_13110_ _15187_/A _13072_/X _13104_/X _14708_/A vssd1 vssd1 vccd1 vccd1 _13110_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_124_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14090_ _26785_/Q _26429_/Q _14114_/S vssd1 vssd1 vccd1 vccd1 _14090_/X sky130_fd_sc_hd__mux2_1
X_26076_ _27307_/CLK _26076_/D vssd1 vssd1 vccd1 vccd1 _26076_/Q sky130_fd_sc_hd__dfxtp_1
X_23288_ _23288_/A vssd1 vssd1 vccd1 vccd1 _26586_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13041_ _14269_/S vssd1 vssd1 vccd1 vccd1 _15888_/S sky130_fd_sc_hd__buf_4
XFILLER_4_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22239_ _22239_/A _22239_/B vssd1 vssd1 vccd1 vccd1 _22317_/A sky130_fd_sc_hd__or2_2
X_25027_ _25027_/A vssd1 vssd1 vccd1 vccd1 _25027_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_180_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16800_ _17998_/A _16800_/B vssd1 vssd1 vccd1 vccd1 _16801_/A sky130_fd_sc_hd__or2_2
X_17780_ _17780_/A _17780_/B vssd1 vssd1 vccd1 vccd1 _19355_/A sky130_fd_sc_hd__nand2_1
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26978_ _26980_/CLK _26978_/D vssd1 vssd1 vccd1 vccd1 _26978_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_135_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27137_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14992_ _14890_/X _26124_/Q _26025_/Q _14984_/S _14772_/A vssd1 vssd1 vccd1 vccd1
+ _14992_/X sky130_fd_sc_hd__a221o_1
XFILLER_282_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16731_ _25669_/Q vssd1 vssd1 vccd1 vccd1 _22489_/A sky130_fd_sc_hd__buf_4
X_13943_ _13943_/A vssd1 vssd1 vccd1 vccd1 _13943_/X sky130_fd_sc_hd__buf_2
X_25929_ _27221_/CLK _25929_/D vssd1 vssd1 vccd1 vccd1 _25929_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_47_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19450_ _19916_/A _19218_/X _19448_/Y _19449_/Y _19253_/X vssd1 vssd1 vccd1 vccd1
+ _19450_/X sky130_fd_sc_hd__a221o_2
X_16662_ _25985_/Q _25983_/Q _25984_/Q _25982_/Q vssd1 vssd1 vccd1 vccd1 _16662_/X
+ sky130_fd_sc_hd__or4_1
X_13874_ _13431_/A _13870_/X _13873_/X _13863_/A vssd1 vssd1 vccd1 vccd1 _13874_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_35_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18401_ _26946_/Q _18569_/A _18570_/A _26978_/Q vssd1 vssd1 vccd1 vccd1 _18401_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_223_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15613_ _13466_/X _23565_/A _15612_/Y _13214_/A vssd1 vssd1 vccd1 vccd1 _20120_/A
+ sky130_fd_sc_hd__o211ai_4
X_12825_ _12866_/A _12866_/B _25471_/Q vssd1 vssd1 vccd1 vccd1 _12825_/Y sky130_fd_sc_hd__a21oi_1
X_19381_ _19381_/A _19381_/B vssd1 vssd1 vccd1 vccd1 _19382_/B sky130_fd_sc_hd__nor2_1
XFILLER_201_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16593_ _18077_/B vssd1 vssd1 vccd1 vccd1 _16788_/A sky130_fd_sc_hd__buf_4
XFILLER_234_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18332_ _19078_/A _18289_/Y _18306_/X _18331_/X _18895_/A vssd1 vssd1 vccd1 vccd1
+ _18332_/X sky130_fd_sc_hd__a32o_1
X_15544_ _26345_/Q _26605_/Q _15557_/S vssd1 vssd1 vccd1 vccd1 _15544_/X sky130_fd_sc_hd__mux2_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12756_/A vssd1 vssd1 vccd1 vccd1 _12757_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18263_ _18261_/X _18490_/B _18348_/S vssd1 vssd1 vccd1 vccd1 _18263_/X sky130_fd_sc_hd__mux2_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15475_ _25887_/Q _15820_/B vssd1 vssd1 vccd1 vccd1 _15475_/X sky130_fd_sc_hd__or2_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12687_ _25569_/Q vssd1 vssd1 vccd1 vccd1 _17504_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_230_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17214_ _17214_/A vssd1 vssd1 vccd1 vccd1 _25496_/D sky130_fd_sc_hd__clkbuf_1
X_14426_ _12768_/A _25759_/Q _15890_/S _26845_/Q _14331_/X vssd1 vssd1 vccd1 vccd1
+ _14426_/X sky130_fd_sc_hd__o221a_1
XFILLER_147_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18194_ _19455_/C _18194_/B vssd1 vssd1 vccd1 vccd1 _18314_/A sky130_fd_sc_hd__and2_2
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17145_ _17145_/A vssd1 vssd1 vccd1 vccd1 _17146_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14357_ _13007_/A _23517_/A _14356_/X _13025_/A vssd1 vssd1 vccd1 vccd1 _16816_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_7_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13308_ _13477_/A vssd1 vssd1 vccd1 vccd1 _13309_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_116_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17076_ _26240_/Q vssd1 vssd1 vccd1 vccd1 _22361_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_143_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14288_ _14223_/S _14286_/X _14287_/X _13939_/X vssd1 vssd1 vccd1 vccd1 _14292_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16027_ _16023_/X _16026_/X _14806_/A vssd1 vssd1 vccd1 vccd1 _16027_/Y sky130_fd_sc_hd__o21ai_1
X_13239_ _13239_/A vssd1 vssd1 vccd1 vccd1 _13832_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_143_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17978_ _17978_/A _17978_/B _17978_/C vssd1 vssd1 vccd1 vccd1 _18001_/B sky130_fd_sc_hd__nor3_1
XFILLER_226_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19717_ _27104_/Q _19691_/X _19905_/A _19716_/X vssd1 vssd1 vccd1 vccd1 _19717_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16929_ _16907_/X _16978_/C _16928_/X vssd1 vssd1 vccd1 vccd1 _16930_/B sky130_fd_sc_hd__o21a_2
XFILLER_284_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19648_ _27135_/Q _27069_/Q vssd1 vssd1 vccd1 vccd1 _19686_/A sky130_fd_sc_hd__and2_1
XFILLER_225_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19579_ _19579_/A _19579_/B _19579_/C _19579_/D vssd1 vssd1 vccd1 vccd1 _19579_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21610_ _25496_/Q _21620_/B vssd1 vssd1 vccd1 vccd1 _21610_/X sky130_fd_sc_hd__or2_1
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22590_ _22580_/X _22589_/Y _22587_/X vssd1 vssd1 vccd1 vccd1 _26311_/D sky130_fd_sc_hd__a21oi_1
XFILLER_178_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21541_ _21488_/X _25864_/Q _21540_/Y _21518_/X vssd1 vssd1 vccd1 vccd1 _21541_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_178_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24260_ _26977_/Q _24260_/B vssd1 vssd1 vccd1 vccd1 _24266_/C sky130_fd_sc_hd__and2_1
X_21472_ _20668_/A _21415_/X _21459_/X _21471_/X vssd1 vssd1 vccd1 vccd1 _21472_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_194_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23211_ _23211_/A _25393_/B vssd1 vssd1 vccd1 vccd1 _23268_/A sky130_fd_sc_hd__nor2_4
XFILLER_181_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20423_ _25753_/Q vssd1 vssd1 vccd1 vccd1 _20699_/A sky130_fd_sc_hd__buf_6
X_24191_ _26954_/Q _26953_/Q _24191_/C vssd1 vssd1 vccd1 vccd1 _24197_/C sky130_fd_sc_hd__and3_1
XFILLER_147_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23142_ _26520_/Q _23034_/X _23150_/S vssd1 vssd1 vccd1 vccd1 _23143_/A sky130_fd_sc_hd__mux2_1
X_20354_ _20448_/A _20399_/B vssd1 vssd1 vccd1 vccd1 _20354_/X sky130_fd_sc_hd__and2_1
XFILLER_106_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23073_ _23546_/A vssd1 vssd1 vccd1 vccd1 _23073_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20285_ _19725_/X _20284_/Y _20015_/X vssd1 vssd1 vccd1 vccd1 _20289_/A sky130_fd_sc_hd__a21o_1
XFILLER_150_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22024_ _22024_/A vssd1 vssd1 vccd1 vccd1 _26123_/D sky130_fd_sc_hd__clkbuf_1
X_26901_ _26929_/CLK _26901_/D vssd1 vssd1 vccd1 vccd1 _26901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26832_ _27253_/CLK _26832_/D vssd1 vssd1 vccd1 vccd1 _26832_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26763_ _26827_/CLK _26763_/D vssd1 vssd1 vccd1 vccd1 _26763_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23975_ _23975_/A vssd1 vssd1 vccd1 vccd1 _26862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25714_ _26611_/CLK _25714_/D vssd1 vssd1 vccd1 vccd1 _25714_/Q sky130_fd_sc_hd__dfxtp_1
X_22926_ _26439_/Q _22691_/X _22934_/S vssd1 vssd1 vccd1 vccd1 _22927_/A sky130_fd_sc_hd__mux2_1
X_26694_ _27278_/CLK _26694_/D vssd1 vssd1 vccd1 vccd1 _26694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25645_ _27295_/CLK _25645_/D vssd1 vssd1 vccd1 vccd1 _25645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22857_ _22857_/A vssd1 vssd1 vccd1 vccd1 _26408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_271_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21808_ _26034_/Q _20887_/X _21816_/S vssd1 vssd1 vccd1 vccd1 _21809_/A sky130_fd_sc_hd__mux2_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13590_ _13590_/A vssd1 vssd1 vccd1 vccd1 _14173_/B sky130_fd_sc_hd__clkbuf_4
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25576_ _26683_/CLK _25576_/D vssd1 vssd1 vccd1 vccd1 _25576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22788_ _22788_/A vssd1 vssd1 vccd1 vccd1 _26378_/D sky130_fd_sc_hd__clkbuf_1
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27315_ _27315_/CLK _27315_/D vssd1 vssd1 vccd1 vccd1 _27315_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24527_ _24765_/B vssd1 vssd1 vccd1 vccd1 _24625_/A sky130_fd_sc_hd__inv_2
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21739_ _20521_/X _26004_/Q _21743_/S vssd1 vssd1 vccd1 vccd1 _21740_/A sky130_fd_sc_hd__mux2_1
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27246_ _27310_/CLK _27246_/D vssd1 vssd1 vccd1 vccd1 _27246_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ _16378_/S _15257_/X _15259_/X _15040_/X vssd1 vssd1 vccd1 vccd1 _15260_/X
+ sky130_fd_sc_hd__a211o_1
X_24458_ _26309_/Q _24455_/X _24456_/X input222/X _24457_/X vssd1 vssd1 vccd1 vccd1
+ _24458_/X sky130_fd_sc_hd__a221o_1
XFILLER_138_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14211_ _14777_/A _14211_/B _14211_/C vssd1 vssd1 vccd1 vccd1 _14211_/X sky130_fd_sc_hd__or3_1
XFILLER_137_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23409_ _23409_/A vssd1 vssd1 vccd1 vccd1 _26639_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15191_ _14593_/A _15139_/Y _15190_/Y _15079_/A vssd1 vssd1 vccd1 vccd1 _15192_/B
+ sky130_fd_sc_hd__a211o_2
X_27177_ _27198_/CLK _27177_/D vssd1 vssd1 vccd1 vccd1 _27177_/Q sky130_fd_sc_hd__dfxtp_1
X_24389_ _27009_/Q _24357_/X _24388_/Y _24379_/X vssd1 vssd1 vccd1 vccd1 _27009_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26128_ _26240_/CLK _26128_/D vssd1 vssd1 vccd1 vccd1 _26128_/Q sky130_fd_sc_hd__dfxtp_1
X_14142_ input151/X input136/X _14240_/S vssd1 vssd1 vccd1 vccd1 _14142_/X sky130_fd_sc_hd__mux2_8
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14073_ _26525_/Q _26133_/Q _14459_/S vssd1 vssd1 vccd1 vccd1 _14073_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26059_ _26938_/CLK _26059_/D vssd1 vssd1 vccd1 vccd1 _26059_/Q sky130_fd_sc_hd__dfxtp_1
X_18950_ _27085_/Q _19058_/A _19059_/A _27183_/Q _19060_/A vssd1 vssd1 vccd1 vccd1
+ _18950_/X sky130_fd_sc_hd__a221o_1
XFILLER_140_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13024_ _14522_/S _13431_/A _14355_/A _14713_/D vssd1 vssd1 vccd1 vccd1 _13025_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_152_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17901_ _17947_/S vssd1 vssd1 vccd1 vccd1 _17950_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_112_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18881_ _18740_/X _18879_/Y _18880_/X _18887_/B _18777_/X vssd1 vssd1 vccd1 vccd1
+ _18881_/X sky130_fd_sc_hd__o32a_2
XFILLER_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17832_ _18855_/A _17830_/X _18905_/A vssd1 vssd1 vccd1 vccd1 _17833_/B sky130_fd_sc_hd__o21a_1
XFILLER_86_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17763_ _25501_/Q _18443_/A _17733_/X _17761_/X _18468_/A vssd1 vssd1 vccd1 vccd1
+ _17763_/X sky130_fd_sc_hd__o221a_1
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14975_ _17197_/A _14962_/X _14966_/X _14974_/X _14683_/X vssd1 vssd1 vccd1 vccd1
+ _14975_/X sky130_fd_sc_hd__a311o_1
XFILLER_48_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19502_ _19541_/A vssd1 vssd1 vccd1 vccd1 _19502_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16714_ _16714_/A _16714_/B vssd1 vssd1 vccd1 vccd1 _18329_/A sky130_fd_sc_hd__xnor2_4
X_13926_ input112/X input147/X _14488_/S vssd1 vssd1 vccd1 vccd1 _13927_/B sky130_fd_sc_hd__mux2_8
XFILLER_47_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17694_ _17708_/A _17694_/B vssd1 vssd1 vccd1 vccd1 _17694_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_402 _17041_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19433_ _27099_/Q _18751_/X _18752_/X _27197_/Q _18753_/X vssd1 vssd1 vccd1 vccd1
+ _19433_/X sky130_fd_sc_hd__a221o_1
XINSDIODE2_413 _17009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16645_ _12916_/X _16642_/Y _16644_/X vssd1 vssd1 vccd1 vccd1 _16645_/X sky130_fd_sc_hd__o21a_1
X_13857_ _13857_/A vssd1 vssd1 vccd1 vccd1 _13857_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_223_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_424 _12781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_435 _25754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_446 _25733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_457 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19364_ _27227_/Q _19364_/B vssd1 vssd1 vccd1 vccd1 _19364_/X sky130_fd_sc_hd__and2_1
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12808_ _12808_/A _25579_/Q vssd1 vssd1 vccd1 vccd1 _17992_/B sky130_fd_sc_hd__nand2_2
X_16576_ _17055_/A _17055_/B _17055_/C vssd1 vssd1 vccd1 vccd1 _16604_/A sky130_fd_sc_hd__nor3_4
XFILLER_250_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13788_ _26660_/Q _25700_/Q _15408_/A vssd1 vssd1 vccd1 vccd1 _13788_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_468 _20635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_479 _19882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18315_ _17940_/X _17952_/X _18347_/S vssd1 vssd1 vccd1 vccd1 _18315_/X sky130_fd_sc_hd__mux2_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15527_ _17840_/A _15528_/B vssd1 vssd1 vccd1 vccd1 _19016_/S sky130_fd_sc_hd__nand2_2
XFILLER_37_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26917_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19295_ _17787_/A _17786_/A _18733_/X _19294_/X vssd1 vssd1 vccd1 vccd1 _19295_/X
+ sky130_fd_sc_hd__a22o_1
X_12739_ _16591_/A _17995_/B _17669_/B _12738_/X vssd1 vssd1 vccd1 vccd1 _12740_/C
+ sky130_fd_sc_hd__or4b_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18246_ _18806_/A _18231_/X _18245_/X vssd1 vssd1 vccd1 vccd1 _18246_/X sky130_fd_sc_hd__a21o_4
XFILLER_176_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15458_ _26538_/Q _26146_/Q _15459_/S vssd1 vssd1 vccd1 vccd1 _15458_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14409_ _25631_/Q _13933_/A _14401_/B _13557_/A vssd1 vssd1 vccd1 vccd1 _14409_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_237_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18177_ _18806_/A _18157_/X _18176_/X vssd1 vssd1 vccd1 vccd1 _18177_/X sky130_fd_sc_hd__a21o_4
XFILLER_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15389_ _16463_/A _23574_/A _15387_/X _15388_/X vssd1 vssd1 vccd1 vccd1 _16916_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_117_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17128_ _17612_/A vssd1 vssd1 vccd1 vccd1 _17131_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_237_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17059_ _26587_/Q _17003_/X _20796_/C _17051_/X vssd1 vssd1 vccd1 vccd1 _17059_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_143_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20070_ _27148_/Q _27082_/Q vssd1 vssd1 vccd1 vccd1 _20070_/X sky130_fd_sc_hd__or2_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23760_ _23760_/A vssd1 vssd1 vccd1 vccd1 _23760_/X sky130_fd_sc_hd__buf_2
XFILLER_39_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20972_ _20972_/A vssd1 vssd1 vccd1 vccd1 _25860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_272_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22711_ _23754_/A vssd1 vssd1 vccd1 vccd1 _22711_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_281_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23691_ _23690_/X _26749_/Q _23700_/S vssd1 vssd1 vccd1 vccd1 _23692_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25430_ _25430_/A vssd1 vssd1 vccd1 vccd1 _27310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22642_ _24004_/B _23291_/B vssd1 vssd1 vccd1 vccd1 _22724_/A sky130_fd_sc_hd__nor2_8
XFILLER_90_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22573_ _26305_/Q _22578_/B vssd1 vssd1 vccd1 vccd1 _22573_/Y sky130_fd_sc_hd__nand2_1
X_25361_ _27280_/Q _23741_/A _25365_/S vssd1 vssd1 vccd1 vccd1 _25362_/A sky130_fd_sc_hd__mux2_1
XFILLER_278_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27100_ _27176_/CLK _27100_/D vssd1 vssd1 vccd1 vccd1 _27100_/Q sky130_fd_sc_hd__dfxtp_1
X_24312_ _24312_/A _24318_/C vssd1 vssd1 vccd1 vccd1 _24312_/Y sky130_fd_sc_hd__nor2_1
XFILLER_221_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21524_ _21522_/X _21523_/X _21512_/X vssd1 vssd1 vccd1 vccd1 _21524_/X sky130_fd_sc_hd__a21o_1
XFILLER_210_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25292_ _25292_/A vssd1 vssd1 vccd1 vccd1 _27249_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27031_ _27154_/CLK _27031_/D vssd1 vssd1 vccd1 vccd1 _27031_/Q sky130_fd_sc_hd__dfxtp_1
X_24243_ _26971_/Q _24243_/B vssd1 vssd1 vccd1 vccd1 _24250_/C sky130_fd_sc_hd__and2_1
XFILLER_154_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21455_ _25484_/Q _21559_/B vssd1 vssd1 vccd1 vccd1 _21455_/X sky130_fd_sc_hd__or2_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20406_ _20406_/A _20406_/B vssd1 vssd1 vccd1 vccd1 _20443_/C sky130_fd_sc_hd__and2_1
X_24174_ _26948_/Q _24175_/C _24173_/Y vssd1 vssd1 vccd1 vccd1 _26948_/D sky130_fd_sc_hd__o21a_1
XFILLER_108_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21386_ _21581_/A vssd1 vssd1 vccd1 vccd1 _21386_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23125_ _26515_/Q _23124_/X _23131_/S vssd1 vssd1 vccd1 vccd1 _23126_/A sky130_fd_sc_hd__mux2_1
X_20337_ _20337_/A _20337_/B vssd1 vssd1 vccd1 vccd1 _20337_/Y sky130_fd_sc_hd__nand2_1
XFILLER_150_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23056_ _23056_/A vssd1 vssd1 vccd1 vccd1 _26493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_277_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20268_ _27155_/Q _27089_/Q vssd1 vssd1 vccd1 vccd1 _20268_/X sky130_fd_sc_hd__and2_1
XTAP_5302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput102 dout0[63] vssd1 vssd1 vccd1 vccd1 input102/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22007_ _22018_/A vssd1 vssd1 vccd1 vccd1 _22016_/S sky130_fd_sc_hd__buf_4
XTAP_5324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput113 dout1[15] vssd1 vssd1 vccd1 vccd1 input113/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput124 dout1[25] vssd1 vssd1 vccd1 vccd1 input124/X sky130_fd_sc_hd__clkbuf_1
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20199_ _20199_/A _20305_/A vssd1 vssd1 vccd1 vccd1 _20206_/A sky130_fd_sc_hd__nor2_1
XFILLER_49_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput135 dout1[35] vssd1 vssd1 vccd1 vccd1 input135/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput146 dout1[45] vssd1 vssd1 vccd1 vccd1 input146/X sky130_fd_sc_hd__clkbuf_2
XTAP_5357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput157 dout1[55] vssd1 vssd1 vccd1 vccd1 input157/X sky130_fd_sc_hd__clkbuf_2
XFILLER_276_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26815_ _27299_/CLK _26815_/D vssd1 vssd1 vccd1 vccd1 _26815_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput168 dout1[7] vssd1 vssd1 vccd1 vccd1 input168/X sky130_fd_sc_hd__clkbuf_1
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput179 irq[2] vssd1 vssd1 vccd1 vccd1 input179/X sky130_fd_sc_hd__buf_6
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _14760_/A vssd1 vssd1 vccd1 vccd1 _14760_/X sky130_fd_sc_hd__clkbuf_4
X_26746_ _27259_/CLK _26746_/D vssd1 vssd1 vccd1 vccd1 _26746_/Q sky130_fd_sc_hd__dfxtp_1
X_23958_ _23958_/A vssd1 vssd1 vccd1 vccd1 _26854_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13711_ _13711_/A vssd1 vssd1 vccd1 vccd1 _15646_/A sky130_fd_sc_hd__clkbuf_2
X_22909_ _22909_/A vssd1 vssd1 vccd1 vccd1 _26431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26677_ _26677_/CLK _26677_/D vssd1 vssd1 vccd1 vccd1 _26677_/Q sky130_fd_sc_hd__dfxtp_1
X_14691_ _26550_/Q _26158_/Q _14692_/S vssd1 vssd1 vccd1 vccd1 _14691_/X sky130_fd_sc_hd__mux2_1
X_23889_ _23725_/X _26824_/Q _23893_/S vssd1 vssd1 vccd1 vccd1 _23890_/A sky130_fd_sc_hd__mux2_1
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16430_ _14753_/A _16428_/X _16429_/X _14802_/A vssd1 vssd1 vccd1 vccd1 _16430_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_72_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13642_ _14449_/B vssd1 vssd1 vccd1 vccd1 _16419_/B sky130_fd_sc_hd__buf_12
X_25628_ _26940_/CLK _25628_/D vssd1 vssd1 vccd1 vccd1 _25628_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _26513_/Q _26385_/Q _16361_/S vssd1 vssd1 vccd1 vccd1 _16361_/X sky130_fd_sc_hd__mux2_1
X_25559_ _27000_/CLK _25559_/D vssd1 vssd1 vccd1 vccd1 _25559_/Q sky130_fd_sc_hd__dfxtp_1
X_13573_ _14404_/A _13573_/B vssd1 vssd1 vccd1 vccd1 _13573_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18100_ _17242_/B _18556_/A _18557_/A _25534_/Q vssd1 vssd1 vccd1 vccd1 _18100_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _15312_/A vssd1 vssd1 vccd1 vccd1 _15313_/A sky130_fd_sc_hd__buf_4
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19080_ _25743_/Q _19081_/B vssd1 vssd1 vccd1 vccd1 _19146_/C sky130_fd_sc_hd__and2_2
XFILLER_8_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _16292_/A _16292_/B vssd1 vssd1 vccd1 vccd1 _16292_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18031_ _20626_/A _19879_/A vssd1 vssd1 vccd1 vccd1 _18032_/B sky130_fd_sc_hd__nand2_1
XFILLER_258_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15243_ _15243_/A vssd1 vssd1 vccd1 vccd1 _15244_/A sky130_fd_sc_hd__buf_2
X_27229_ _27230_/CLK _27229_/D vssd1 vssd1 vccd1 vccd1 _27229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15174_ _15174_/A vssd1 vssd1 vccd1 vccd1 _15384_/S sky130_fd_sc_hd__buf_4
XFILLER_181_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14125_ _12813_/A _16827_/B _14124_/X _14560_/S vssd1 vssd1 vccd1 vccd1 _14127_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19982_ _19982_/A _19982_/B _19982_/C vssd1 vssd1 vccd1 vccd1 _19984_/B sky130_fd_sc_hd__and3_1
XFILLER_126_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_150_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27228_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_207_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14056_ _13520_/A _25763_/Q _14391_/S _26849_/Q _14458_/S vssd1 vssd1 vccd1 vccd1
+ _14056_/X sky130_fd_sc_hd__o221a_1
X_18933_ _18973_/A vssd1 vssd1 vccd1 vccd1 _18933_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ _13007_/A vssd1 vssd1 vccd1 vccd1 _13008_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_122_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18864_ _19018_/A _18864_/B _18864_/C _18864_/D vssd1 vssd1 vccd1 vccd1 _18864_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_67_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17815_ _18539_/B _18539_/C _18539_/D _18539_/A vssd1 vssd1 vccd1 vccd1 _18593_/B
+ sky130_fd_sc_hd__o31a_4
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18795_ _18838_/A _18795_/B vssd1 vssd1 vccd1 vccd1 _18795_/Y sky130_fd_sc_hd__xnor2_1
XTAP_5880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17746_ _18116_/B _17740_/C vssd1 vssd1 vccd1 vccd1 _18102_/A sky130_fd_sc_hd__or2b_1
X_14958_ _12706_/A _14949_/X _14957_/X _17195_/A vssd1 vssd1 vccd1 vccd1 _14958_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_82_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13909_ _18498_/S _13909_/B vssd1 vssd1 vccd1 vccd1 _17813_/A sky130_fd_sc_hd__or2_2
X_17677_ _17697_/A vssd1 vssd1 vccd1 vccd1 _17738_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14889_ _26809_/Q _26453_/Q _14991_/S vssd1 vssd1 vccd1 vccd1 _14889_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_210 _15190_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_221 _20055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_232 _19268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16628_ _18862_/S _16628_/B vssd1 vssd1 vccd1 vccd1 _17816_/B sky130_fd_sc_hd__nor2_1
X_19416_ _18929_/X _19412_/X _19415_/Y _18782_/X vssd1 vssd1 vccd1 vccd1 _19416_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_243 _16691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_254 _16893_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_265 _20686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_276 _27126_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19347_ _19315_/A _19346_/C _25751_/Q vssd1 vssd1 vccd1 vccd1 _19348_/B sky130_fd_sc_hd__a21oi_1
XINSDIODE2_287 _25819_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16559_ _19388_/A vssd1 vssd1 vccd1 vccd1 _17055_/B sky130_fd_sc_hd__clkinv_2
XINSDIODE2_298 _26143_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19278_ _19577_/A _19256_/B _19328_/S vssd1 vssd1 vccd1 vccd1 _19278_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18229_ _18287_/B _18229_/B vssd1 vssd1 vccd1 vccd1 _18229_/X sky130_fd_sc_hd__or2_1
XFILLER_164_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21240_ _21228_/Y _21238_/Y _21273_/A vssd1 vssd1 vccd1 vccd1 _21240_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_191_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21171_ _25928_/Q _21166_/X _21167_/X input28/X vssd1 vssd1 vccd1 vccd1 _21172_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20122_ _25741_/Q vssd1 vssd1 vccd1 vccd1 _20668_/A sky130_fd_sc_hd__buf_8
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24930_ _24957_/A vssd1 vssd1 vccd1 vccd1 _24930_/X sky130_fd_sc_hd__clkbuf_2
X_20053_ _19991_/X _20051_/X _20052_/X vssd1 vssd1 vccd1 vccd1 _20053_/Y sky130_fd_sc_hd__o21ai_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24861_ _20677_/A _24848_/X _24729_/Y _24849_/X vssd1 vssd1 vccd1 vccd1 _24861_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_85_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26600_ _27307_/CLK _26600_/D vssd1 vssd1 vccd1 vccd1 _26600_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23812_ _23858_/S vssd1 vssd1 vccd1 vccd1 _23821_/S sky130_fd_sc_hd__buf_6
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24792_ _20628_/A _24789_/X _24649_/Y _24791_/X vssd1 vssd1 vccd1 vccd1 _24792_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26531_ _26531_/CLK _26531_/D vssd1 vssd1 vccd1 vccd1 _26531_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23743_ _23743_/A vssd1 vssd1 vccd1 vccd1 _26765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20955_ _23770_/A vssd1 vssd1 vccd1 vccd1 _20955_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26462_ _26462_/CLK _26462_/D vssd1 vssd1 vccd1 vccd1 _26462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23674_ _26743_/Q _23597_/X _23678_/S vssd1 vssd1 vccd1 vccd1 _23675_/A sky130_fd_sc_hd__mux2_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ _20886_/A vssd1 vssd1 vccd1 vccd1 _25833_/D sky130_fd_sc_hd__clkbuf_1
X_25413_ _23712_/X _27303_/Q _25415_/S vssd1 vssd1 vccd1 vccd1 _25414_/A sky130_fd_sc_hd__mux2_1
X_22625_ _26326_/Q _26325_/Q vssd1 vssd1 vccd1 vccd1 _22625_/X sky130_fd_sc_hd__and2_1
X_26393_ _27265_/CLK _26393_/D vssd1 vssd1 vccd1 vccd1 _26393_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25344_ _25344_/A vssd1 vssd1 vccd1 vccd1 _27272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22556_ _26298_/Q _22565_/B vssd1 vssd1 vccd1 vccd1 _22556_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21507_ _21507_/A vssd1 vssd1 vccd1 vccd1 _21574_/B sky130_fd_sc_hd__clkbuf_1
X_25275_ _25275_/A vssd1 vssd1 vccd1 vccd1 _27241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22487_ _22487_/A _22491_/B vssd1 vssd1 vccd1 vccd1 _22488_/A sky130_fd_sc_hd__and2_1
X_27014_ _27014_/CLK _27014_/D vssd1 vssd1 vccd1 vccd1 _27014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24226_ _26965_/Q _24227_/C _24225_/Y vssd1 vssd1 vccd1 vccd1 _26965_/D sky130_fd_sc_hd__o21a_1
X_21438_ input48/X input83/X _21489_/S vssd1 vssd1 vccd1 vccd1 _21439_/A sky130_fd_sc_hd__mux2_8
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24157_ _26943_/Q _26942_/Q _24157_/C vssd1 vssd1 vccd1 vccd1 _24159_/A sky130_fd_sc_hd__and3_1
XFILLER_181_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21369_ _20648_/A _21343_/X _21350_/X _21368_/X vssd1 vssd1 vccd1 vccd1 _21369_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_218_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23108_ _23581_/A vssd1 vssd1 vccd1 vccd1 _23108_/X sky130_fd_sc_hd__clkbuf_2
X_24088_ _24088_/A vssd1 vssd1 vccd1 vccd1 _26912_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15930_ _26665_/Q _25705_/Q _15930_/S vssd1 vssd1 vccd1 vccd1 _15930_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23039_ _26488_/Q _23034_/X _23051_/S vssd1 vssd1 vccd1 vccd1 _23040_/A sky130_fd_sc_hd__mux2_1
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15861_ _15589_/A _26922_/Q _26406_/Q _15582_/A _15843_/A vssd1 vssd1 vccd1 vccd1
+ _15861_/X sky130_fd_sc_hd__a221o_1
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _17615_/A _17600_/B vssd1 vssd1 vccd1 vccd1 _25581_/D sky130_fd_sc_hd__nor2_1
XTAP_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14812_ _14810_/X _14811_/X _16524_/A vssd1 vssd1 vccd1 vccd1 _14812_/X sky130_fd_sc_hd__mux2_1
XFILLER_264_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18580_ _18666_/A _18580_/B vssd1 vssd1 vccd1 vccd1 _18580_/Y sky130_fd_sc_hd__nor2_1
X_15792_ _12871_/A _15790_/Y _15791_/Y _13575_/X _13929_/X vssd1 vssd1 vccd1 vccd1
+ _15792_/X sky130_fd_sc_hd__o32a_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _25567_/Q _17529_/X _17516_/X _17530_/X vssd1 vssd1 vccd1 vccd1 _17532_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_26729_ _26889_/CLK _26729_/D vssd1 vssd1 vccd1 vccd1 _26729_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14743_ _14743_/A vssd1 vssd1 vccd1 vccd1 _14744_/A sky130_fd_sc_hd__buf_2
XFILLER_18_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17462_ _26243_/Q _17455_/X _21206_/A _25971_/Q vssd1 vssd1 vccd1 vccd1 _21208_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14674_ _25899_/Q _16501_/B vssd1 vssd1 vccd1 vccd1 _14674_/X sky130_fd_sc_hd__or2_1
XFILLER_33_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19201_ _27156_/Q _19334_/B vssd1 vssd1 vccd1 vccd1 _19201_/X sky130_fd_sc_hd__or2_1
X_16413_ _16463_/A _23597_/A _15388_/X vssd1 vssd1 vccd1 vccd1 _16413_/X sky130_fd_sc_hd__o21a_1
XFILLER_232_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13625_ _15970_/S _13625_/B vssd1 vssd1 vccd1 vccd1 _13625_/X sky130_fd_sc_hd__or2_1
X_17393_ _17430_/A _17399_/C vssd1 vssd1 vccd1 vccd1 _17393_/Y sky130_fd_sc_hd__nor2_1
XFILLER_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19132_ _27122_/Q _19056_/X _19130_/X _19131_/X vssd1 vssd1 vccd1 vccd1 _19132_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_158_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16344_ _15111_/A _26709_/Q _26837_/Q _16361_/S _14770_/A vssd1 vssd1 vccd1 vccd1
+ _16344_/X sky130_fd_sc_hd__a221o_1
X_13556_ _13556_/A vssd1 vssd1 vccd1 vccd1 _13557_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19063_ _19063_/A vssd1 vssd1 vccd1 vccd1 _19063_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16275_ _14763_/A _16273_/X _16274_/X vssd1 vssd1 vccd1 vccd1 _16275_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13487_ _26630_/Q _26726_/Q _13792_/S vssd1 vssd1 vccd1 vccd1 _13487_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18014_ _18059_/A vssd1 vssd1 vccd1 vccd1 _18721_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15226_ _27287_/Q _26480_/Q _16428_/S vssd1 vssd1 vccd1 vccd1 _15226_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput406 _17018_/X vssd1 vssd1 vccd1 vccd1 din0[8] sky130_fd_sc_hd__buf_2
XFILLER_126_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput417 _25952_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[16] sky130_fd_sc_hd__buf_2
XFILLER_5_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput428 _25962_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[26] sky130_fd_sc_hd__buf_2
XFILLER_172_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15157_ _15155_/X _15156_/X _15263_/S vssd1 vssd1 vccd1 vccd1 _15157_/X sky130_fd_sc_hd__mux2_1
Xoutput439 _25943_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[7] sky130_fd_sc_hd__buf_2
XFILLER_153_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14108_ _26493_/Q _26365_/Q _14257_/A vssd1 vssd1 vccd1 vccd1 _14108_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15088_ _26514_/Q _26386_/Q _15088_/S vssd1 vssd1 vccd1 vccd1 _15088_/X sky130_fd_sc_hd__mux2_1
X_19965_ _20644_/A vssd1 vssd1 vccd1 vccd1 _19965_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14039_ _14028_/X _14036_/X _14038_/X _14325_/S _13557_/A vssd1 vssd1 vccd1 vccd1
+ _14039_/X sky130_fd_sc_hd__o221a_1
XFILLER_141_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18916_ _27116_/Q _19056_/A _18914_/X _18915_/X vssd1 vssd1 vccd1 vccd1 _18916_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_256_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19896_ _19896_/A _19896_/B vssd1 vssd1 vccd1 vccd1 _19896_/Y sky130_fd_sc_hd__nand2_1
XFILLER_267_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18847_ _18967_/A _18847_/B vssd1 vssd1 vccd1 vccd1 _18847_/Y sky130_fd_sc_hd__nand2_2
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18778_ _18740_/X _18774_/Y _18776_/X _18787_/B _18777_/X vssd1 vssd1 vccd1 vccd1
+ _18778_/X sky130_fd_sc_hd__o32a_2
XFILLER_227_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17729_ _17732_/A _17730_/B vssd1 vssd1 vccd1 vccd1 _18460_/A sky130_fd_sc_hd__and2_2
XFILLER_242_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20740_ _20740_/A vssd1 vssd1 vccd1 vccd1 _25767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20671_ _21878_/A vssd1 vssd1 vccd1 vccd1 _20671_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22410_ _22387_/A _22385_/X _22390_/A vssd1 vssd1 vccd1 vccd1 _22410_/X sky130_fd_sc_hd__o21ba_1
X_23390_ _23390_/A vssd1 vssd1 vccd1 vccd1 _26630_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22341_ _22337_/X _17078_/X _26226_/Q vssd1 vssd1 vccd1 vccd1 _22341_/X sky130_fd_sc_hd__a21o_1
XFILLER_176_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22272_ _26202_/Q _22264_/X _22270_/X _26303_/Q _22271_/X vssd1 vssd1 vccd1 vccd1
+ _22272_/X sky130_fd_sc_hd__a221o_1
X_25060_ _25139_/A vssd1 vssd1 vccd1 vccd1 _25060_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24011_ _26878_/Q _23517_/X _24015_/S vssd1 vssd1 vccd1 vccd1 _24012_/A sky130_fd_sc_hd__mux2_1
X_21223_ _21562_/D _21866_/B vssd1 vssd1 vccd1 vccd1 _21279_/A sky130_fd_sc_hd__and2_1
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21154_ _21154_/A _21154_/B vssd1 vssd1 vccd1 vccd1 _21155_/A sky130_fd_sc_hd__or2_1
XFILLER_137_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20105_ _27149_/Q _27083_/Q vssd1 vssd1 vccd1 vccd1 _20105_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25962_ _26995_/CLK _25962_/D vssd1 vssd1 vccd1 vccd1 _25962_/Q sky130_fd_sc_hd__dfxtp_1
X_21085_ _25904_/Q _21074_/X _21077_/X input32/X vssd1 vssd1 vccd1 vccd1 _21086_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_120_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24913_ _24957_/A vssd1 vssd1 vccd1 vccd1 _24913_/X sky130_fd_sc_hd__clkbuf_2
X_20036_ _20662_/A _19708_/A _20035_/Y _19661_/X vssd1 vssd1 vccd1 vccd1 _20061_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25893_ _27287_/CLK _25893_/D vssd1 vssd1 vccd1 vccd1 _25893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_273_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24844_ _27117_/Q _24856_/B vssd1 vssd1 vccd1 vccd1 _24844_/Y sky130_fd_sc_hd__nand2_1
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24775_ _27100_/Q _24636_/X _24774_/X vssd1 vssd1 vccd1 vccd1 _27100_/D sky130_fd_sc_hd__o21ba_1
X_21987_ _21987_/A vssd1 vssd1 vccd1 vccd1 _26106_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26514_ _27321_/CLK _26514_/D vssd1 vssd1 vccd1 vccd1 _26514_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23726_ _23725_/X _26760_/Q _23732_/S vssd1 vssd1 vccd1 vccd1 _23727_/A sky130_fd_sc_hd__mux2_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ _20938_/A vssd1 vssd1 vccd1 vccd1 _25849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26445_ _27284_/CLK _26445_/D vssd1 vssd1 vccd1 vccd1 _26445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23657_ _23657_/A vssd1 vssd1 vccd1 vccd1 _26735_/D sky130_fd_sc_hd__clkbuf_1
X_20869_ _25321_/A vssd1 vssd1 vccd1 vccd1 _24004_/B sky130_fd_sc_hd__buf_4
X_13410_ _15826_/S vssd1 vssd1 vccd1 vccd1 _13410_/X sky130_fd_sc_hd__clkbuf_4
X_22608_ _26318_/Q _22618_/B vssd1 vssd1 vccd1 vccd1 _22608_/Y sky130_fd_sc_hd__nand2_1
X_14390_ _14388_/X _14389_/X _14390_/S vssd1 vssd1 vccd1 vccd1 _14390_/X sky130_fd_sc_hd__mux2_2
X_26376_ _26604_/CLK _26376_/D vssd1 vssd1 vccd1 vccd1 _26376_/Q sky130_fd_sc_hd__dfxtp_1
X_23588_ _26708_/Q _23587_/X _23588_/S vssd1 vssd1 vccd1 vccd1 _23589_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25327_ _25327_/A vssd1 vssd1 vccd1 vccd1 _27264_/D sky130_fd_sc_hd__clkbuf_1
X_13341_ _15333_/A _13331_/X _13335_/X _14751_/A vssd1 vssd1 vccd1 vccd1 _13369_/A
+ sky130_fd_sc_hd__o211a_1
X_22539_ _22554_/A vssd1 vssd1 vccd1 vccd1 _22632_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_194_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16060_ _27282_/Q _26475_/Q _16060_/S vssd1 vssd1 vccd1 vccd1 _16060_/X sky130_fd_sc_hd__mux2_1
X_25258_ _23696_/X _27234_/Q _25260_/S vssd1 vssd1 vccd1 vccd1 _25259_/A sky130_fd_sc_hd__mux2_1
X_13272_ _14228_/A vssd1 vssd1 vccd1 vccd1 _13545_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_185_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15011_ _14724_/X _14941_/Y _15010_/X _14827_/X vssd1 vssd1 vccd1 vccd1 _19374_/A
+ sky130_fd_sc_hd__a211o_4
X_24209_ _24938_/A vssd1 vssd1 vccd1 vccd1 _24209_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_185_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25189_ _25198_/A vssd1 vssd1 vccd1 vccd1 _25189_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19750_ _27137_/Q _27071_/Q vssd1 vssd1 vccd1 vccd1 _19750_/Y sky130_fd_sc_hd__nor2_1
XFILLER_231_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16962_ _16962_/A vssd1 vssd1 vccd1 vccd1 _16983_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_89_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18701_ _25512_/Q _18444_/X _18698_/X _18700_/X _18469_/X vssd1 vssd1 vccd1 vccd1
+ _18701_/X sky130_fd_sc_hd__o221a_1
XFILLER_238_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15913_ _15913_/A vssd1 vssd1 vccd1 vccd1 _23552_/A sky130_fd_sc_hd__clkbuf_4
X_19681_ _22474_/A _19638_/X _19680_/X _19566_/X vssd1 vssd1 vccd1 vccd1 _25662_/D
+ sky130_fd_sc_hd__o211a_1
X_16893_ _16893_/A _16893_/B vssd1 vssd1 vccd1 vccd1 _16894_/A sky130_fd_sc_hd__and2_1
XFILLER_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15844_ _15576_/A _15841_/X _15843_/X _13762_/X vssd1 vssd1 vccd1 vccd1 _15844_/X
+ sky130_fd_sc_hd__o211a_1
X_18632_ _20657_/A vssd1 vssd1 vccd1 vccd1 _22368_/A sky130_fd_sc_hd__buf_6
XFILLER_265_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15775_ _25812_/Q _27246_/Q _15775_/S vssd1 vssd1 vccd1 vccd1 _15776_/B sky130_fd_sc_hd__mux2_1
X_18563_ _27141_/Q vssd1 vssd1 vccd1 vccd1 _19870_/A sky130_fd_sc_hd__clkbuf_4
X_12987_ _25587_/Q vssd1 vssd1 vccd1 vccd1 _13029_/A sky130_fd_sc_hd__inv_2
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _16439_/A vssd1 vssd1 vccd1 vccd1 _16521_/A sky130_fd_sc_hd__clkbuf_4
X_17514_ _17514_/A _20236_/A _17514_/C _17513_/X vssd1 vssd1 vccd1 vccd1 _19650_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_32_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18494_ _18898_/A _18488_/Y _18493_/X vssd1 vssd1 vccd1 vccd1 _18495_/B sky130_fd_sc_hd__o21ai_2
XFILLER_33_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17445_ _19570_/A _19570_/B _19570_/C _19570_/D vssd1 vssd1 vccd1 vccd1 _20236_/A
+ sky130_fd_sc_hd__nor4_4
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14657_ _27261_/Q _16501_/B vssd1 vssd1 vccd1 vccd1 _14657_/X sky130_fd_sc_hd__or2_1
XFILLER_220_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13608_ _15885_/A vssd1 vssd1 vccd1 vccd1 _13608_/X sky130_fd_sc_hd__buf_2
XFILLER_177_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17376_ _17375_/X _17379_/C _17366_/X vssd1 vssd1 vccd1 vccd1 _17376_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14588_ _16170_/A vssd1 vssd1 vccd1 vccd1 _15290_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19115_ _25744_/Q _19146_/C vssd1 vssd1 vccd1 vccd1 _19115_/Y sky130_fd_sc_hd__xnor2_4
X_16327_ _15165_/X _16325_/X _16326_/X vssd1 vssd1 vccd1 vccd1 _16328_/B sky130_fd_sc_hd__o21ai_1
X_13539_ _13955_/A vssd1 vssd1 vccd1 vccd1 _13540_/A sky130_fd_sc_hd__buf_4
XFILLER_174_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19046_ _19046_/A _19046_/B vssd1 vssd1 vccd1 vccd1 _19046_/Y sky130_fd_sc_hd__nand2_1
X_16258_ _15085_/A _16255_/X _16257_/X _15333_/X vssd1 vssd1 vccd1 vccd1 _16258_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15209_ _26644_/Q _26740_/Q _15209_/S vssd1 vssd1 vccd1 vccd1 _15209_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16189_ _27316_/Q _26573_/Q _16189_/S vssd1 vssd1 vccd1 vccd1 _16189_/X sky130_fd_sc_hd__mux2_1
XFILLER_245_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19948_ _19882_/B _18710_/Y _19671_/A _19947_/X vssd1 vssd1 vccd1 vccd1 _19948_/X
+ sky130_fd_sc_hd__o31a_1
XINSDIODE2_9 _18655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19879_ _19879_/A vssd1 vssd1 vccd1 vccd1 _19879_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_255_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21910_ _21910_/A vssd1 vssd1 vccd1 vccd1 _26072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22890_ _23211_/A _23788_/A vssd1 vssd1 vccd1 vccd1 _22947_/A sky130_fd_sc_hd__nor2_8
XFILLER_255_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21841_ _26049_/Q _20935_/X _21849_/S vssd1 vssd1 vccd1 vccd1 _21842_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24560_ _27041_/Q _24546_/X _24559_/Y _24551_/X vssd1 vssd1 vccd1 vccd1 _27041_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_70_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21772_ _20584_/X _26019_/Q _21776_/S vssd1 vssd1 vccd1 vccd1 _21773_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23511_ _23610_/S vssd1 vssd1 vccd1 vccd1 _23524_/S sky130_fd_sc_hd__clkbuf_4
X_20723_ _20723_/A vssd1 vssd1 vccd1 vccd1 _25759_/D sky130_fd_sc_hd__clkbuf_1
X_24491_ _24392_/X _25620_/Q _24490_/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__o21ai_4
XFILLER_168_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26230_ _26297_/CLK _26230_/D vssd1 vssd1 vccd1 vccd1 _26230_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_211_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23442_ _23442_/A vssd1 vssd1 vccd1 vccd1 _26653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20654_ _20654_/A _20656_/B vssd1 vssd1 vccd1 vccd1 _20654_/X sky130_fd_sc_hd__or2_1
XFILLER_165_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26161_ _27264_/CLK _26161_/D vssd1 vssd1 vccd1 vccd1 _26161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23373_ _26623_/Q _23047_/X _23375_/S vssd1 vssd1 vccd1 vccd1 _23374_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20585_ _20584_/X _25714_/Q _20593_/S vssd1 vssd1 vccd1 vccd1 _20586_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25112_ _25137_/A vssd1 vssd1 vccd1 vccd1 _25112_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22324_ _26220_/Q _22315_/X _22323_/X _22319_/X vssd1 vssd1 vccd1 vccd1 _26220_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26092_ _27324_/CLK _26092_/D vssd1 vssd1 vccd1 vccd1 _26092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25043_ _25142_/A vssd1 vssd1 vccd1 vccd1 _25043_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22255_ _22270_/A vssd1 vssd1 vccd1 vccd1 _22255_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21206_ _21206_/A vssd1 vssd1 vccd1 vccd1 _21562_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22186_ _22249_/A vssd1 vssd1 vccd1 vccd1 _22186_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_279_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21137_ _21137_/A vssd1 vssd1 vccd1 vccd1 _25918_/D sky130_fd_sc_hd__clkbuf_1
X_26994_ _26996_/CLK _26994_/D vssd1 vssd1 vccd1 vccd1 _26994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25945_ _27022_/CLK _25945_/D vssd1 vssd1 vccd1 vccd1 _25945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21068_ _21174_/A vssd1 vssd1 vccd1 vccd1 _21138_/A sky130_fd_sc_hd__buf_2
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12910_ _14025_/A _13923_/B _13397_/B vssd1 vssd1 vccd1 vccd1 _15871_/A sky130_fd_sc_hd__nor3_2
XFILLER_150_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20019_ _19833_/X _20030_/B _20018_/Y _20248_/A vssd1 vssd1 vccd1 vccd1 _20020_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25876_ _26595_/CLK _25876_/D vssd1 vssd1 vccd1 vccd1 _25876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13890_ _13890_/A vssd1 vssd1 vccd1 vccd1 _13890_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_273_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12841_ input122/X input157/X _13741_/S vssd1 vssd1 vccd1 vccd1 _17623_/C sky130_fd_sc_hd__mux2_8
X_24827_ _24825_/Y _24826_/X _24816_/X vssd1 vssd1 vccd1 vccd1 _27112_/D sky130_fd_sc_hd__a21oi_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15560_ _15556_/X _15559_/X _16072_/S vssd1 vssd1 vccd1 vccd1 _15560_/X sky130_fd_sc_hd__mux2_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24758_ _24765_/A _24758_/B vssd1 vssd1 vccd1 vccd1 _25151_/A sky130_fd_sc_hd__nand2_4
XFILLER_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _12772_/A vssd1 vssd1 vccd1 vccd1 _12773_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_243_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _12767_/A _25829_/Q _26029_/Q _14169_/B _14515_/S vssd1 vssd1 vccd1 vccd1
+ _14511_/X sky130_fd_sc_hd__a221o_1
XFILLER_187_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23709_ _23709_/A vssd1 vssd1 vccd1 vccd1 _23709_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15491_ _15491_/A vssd1 vssd1 vccd1 vccd1 _15491_/X sky130_fd_sc_hd__buf_2
XFILLER_14_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24689_ _24936_/A vssd1 vssd1 vccd1 vccd1 _24690_/B sky130_fd_sc_hd__clkinv_2
XFILLER_70_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _25466_/A vssd1 vssd1 vccd1 vccd1 _22535_/B sky130_fd_sc_hd__buf_12
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26428_ _27267_/CLK _26428_/D vssd1 vssd1 vccd1 vccd1 _26428_/Q sky130_fd_sc_hd__dfxtp_2
X_14442_ _13172_/A _14421_/X _14441_/X _13025_/A vssd1 vssd1 vccd1 vccd1 _16813_/C
+ sky130_fd_sc_hd__o31a_4
XFILLER_202_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17161_ _20707_/C vssd1 vssd1 vccd1 vccd1 _17195_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14373_ _26910_/Q _26394_/Q _14389_/S vssd1 vssd1 vccd1 vccd1 _14373_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26359_ _26917_/CLK _26359_/D vssd1 vssd1 vccd1 vccd1 _26359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16112_ _13221_/A _16109_/X _16111_/X _14751_/A vssd1 vssd1 vccd1 vccd1 _16117_/A
+ sky130_fd_sc_hd__o211a_1
X_13324_ _16111_/A vssd1 vssd1 vccd1 vccd1 _16088_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17092_ _26235_/Q _17089_/X _22210_/A vssd1 vssd1 vccd1 vccd1 _22121_/A sky130_fd_sc_hd__o21a_1
XFILLER_196_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16043_ _17838_/A _16043_/B vssd1 vssd1 vccd1 vccd1 _16043_/Y sky130_fd_sc_hd__nand2_1
X_13255_ _13255_/A vssd1 vssd1 vccd1 vccd1 _13255_/X sky130_fd_sc_hd__buf_4
XFILLER_170_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_57_wb_clk_i clkbuf_leaf_57_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _26467_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13186_ _25597_/Q _13249_/A vssd1 vssd1 vccd1 vccd1 _13256_/A sky130_fd_sc_hd__nor2_1
XFILLER_43_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19802_ _20639_/A _19708_/A _19801_/X _19661_/X vssd1 vssd1 vccd1 vccd1 _19803_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17994_ _18861_/A vssd1 vssd1 vccd1 vccd1 _18366_/A sky130_fd_sc_hd__buf_4
XFILLER_96_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19733_ _19704_/A _19704_/B _19710_/Y vssd1 vssd1 vccd1 vccd1 _19733_/X sky130_fd_sc_hd__a21o_1
X_16945_ _16332_/X _16952_/A _16887_/A vssd1 vssd1 vccd1 vccd1 _16948_/A sky130_fd_sc_hd__o21a_1
XFILLER_237_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19664_ _19769_/B vssd1 vssd1 vccd1 vccd1 _20055_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16876_ _16876_/A vssd1 vssd1 vccd1 vccd1 _16876_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18615_ _18615_/A vssd1 vssd1 vccd1 vccd1 _19367_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_237_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15827_ _15821_/X _15823_/X _15826_/X _15819_/S _14362_/A vssd1 vssd1 vccd1 vccd1
+ _15827_/X sky130_fd_sc_hd__o221a_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19595_ _20189_/B vssd1 vssd1 vccd1 vccd1 _19774_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_252_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15758_ _26079_/Q _25884_/Q _15758_/S vssd1 vssd1 vccd1 vccd1 _15758_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18546_ _18546_/A vssd1 vssd1 vccd1 vccd1 _18546_/Y sky130_fd_sc_hd__inv_2
XFILLER_252_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14709_ _14709_/A vssd1 vssd1 vccd1 vccd1 _14710_/A sky130_fd_sc_hd__clkbuf_4
X_15689_ _16111_/A _15689_/B vssd1 vssd1 vccd1 vccd1 _15689_/X sky130_fd_sc_hd__or2_1
X_18477_ _19256_/A _18424_/A _18431_/X _18476_/X vssd1 vssd1 vccd1 vccd1 _18477_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_100_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17428_ _17428_/A _17428_/B _17434_/C vssd1 vssd1 vccd1 vccd1 _25560_/D sky130_fd_sc_hd__nor3_1
XFILLER_178_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17359_ _17356_/X _17360_/C _25539_/Q vssd1 vssd1 vccd1 vccd1 _17361_/B sky130_fd_sc_hd__a21oi_1
XFILLER_220_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20370_ _20370_/A _20370_/B vssd1 vssd1 vccd1 vccd1 _20370_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_277_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19029_ _25519_/Q _18810_/X _19026_/X _19028_/X _18832_/X vssd1 vssd1 vccd1 vccd1
+ _19029_/X sky130_fd_sc_hd__o221a_1
XFILLER_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22040_ _26130_/Q _20878_/X _22044_/S vssd1 vssd1 vccd1 vccd1 _22041_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23991_ _23991_/A vssd1 vssd1 vccd1 vccd1 _26869_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25730_ _26271_/CLK _25730_/D vssd1 vssd1 vccd1 vccd1 _25730_/Q sky130_fd_sc_hd__dfxtp_4
X_22942_ _22942_/A vssd1 vssd1 vccd1 vccd1 _26446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25661_ _25661_/CLK _25661_/D vssd1 vssd1 vccd1 vccd1 _25661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22873_ _26416_/Q _22720_/X _22873_/S vssd1 vssd1 vccd1 vccd1 _22874_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24612_ _27060_/Q _24602_/X _24611_/Y _24606_/X vssd1 vssd1 vccd1 vccd1 _27060_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21824_ _21824_/A vssd1 vssd1 vccd1 vccd1 _26041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_271_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25592_ _25596_/CLK _25592_/D vssd1 vssd1 vccd1 vccd1 _25592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24543_ _25206_/B _24543_/B vssd1 vssd1 vccd1 vccd1 _24544_/B sky130_fd_sc_hd__or2_2
XFILLER_93_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21755_ _21755_/A vssd1 vssd1 vccd1 vccd1 _26011_/D sky130_fd_sc_hd__clkbuf_1
XPHY_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27262_ _27326_/CLK _27262_/D vssd1 vssd1 vccd1 vccd1 _27262_/Q sky130_fd_sc_hd__dfxtp_1
X_20706_ _20706_/A vssd1 vssd1 vccd1 vccd1 _26261_/D sky130_fd_sc_hd__clkbuf_1
X_24474_ _24474_/A vssd1 vssd1 vccd1 vccd1 _24474_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_197_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21686_ _21686_/A vssd1 vssd1 vccd1 vccd1 _25982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26213_ _26980_/CLK _26213_/D vssd1 vssd1 vccd1 vccd1 _26213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23425_ _23425_/A vssd1 vssd1 vccd1 vccd1 _26646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20637_ _20637_/A _20643_/B vssd1 vssd1 vccd1 vccd1 _20637_/X sky130_fd_sc_hd__or2_1
X_27193_ _27196_/CLK _27193_/D vssd1 vssd1 vccd1 vccd1 _27193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26144_ _26673_/CLK _26144_/D vssd1 vssd1 vccd1 vccd1 _26144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23356_ _23356_/A vssd1 vssd1 vccd1 vccd1 _26616_/D sky130_fd_sc_hd__clkbuf_1
X_20568_ _20567_/X _25710_/Q _20572_/S vssd1 vssd1 vccd1 vccd1 _20569_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22307_ _26214_/Q _22299_/X _22306_/X _22304_/X vssd1 vssd1 vccd1 vccd1 _26214_/D
+ sky130_fd_sc_hd__o211a_1
X_26075_ _27305_/CLK _26075_/D vssd1 vssd1 vccd1 vccd1 _26075_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_166_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23287_ _26586_/Q input249/X _23289_/S vssd1 vssd1 vccd1 vccd1 _23288_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20499_ _23517_/A vssd1 vssd1 vccd1 vccd1 _23693_/A sky130_fd_sc_hd__buf_2
XFILLER_166_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13040_ _14513_/S vssd1 vssd1 vccd1 vccd1 _14269_/S sky130_fd_sc_hd__clkbuf_2
X_25026_ _20635_/A _25003_/X _25025_/X vssd1 vssd1 vccd1 vccd1 _25026_/Y sky130_fd_sc_hd__o21ai_1
X_22238_ _22270_/A vssd1 vssd1 vccd1 vccd1 _22238_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22169_ _22200_/A vssd1 vssd1 vccd1 vccd1 _22169_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_278_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14991_ _26548_/Q _26156_/Q _14991_/S vssd1 vssd1 vccd1 vccd1 _14991_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26977_ _26980_/CLK _26977_/D vssd1 vssd1 vccd1 vccd1 _26977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13942_ _26626_/Q _26722_/Q _13951_/S vssd1 vssd1 vccd1 vccd1 _13942_/X sky130_fd_sc_hd__mux2_1
X_16730_ _22487_/A _16726_/X _16727_/X _18541_/A vssd1 vssd1 vccd1 vccd1 _16730_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_281_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25928_ _27221_/CLK _25928_/D vssd1 vssd1 vccd1 vccd1 _25928_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_75_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16661_ _16661_/A vssd1 vssd1 vccd1 vccd1 _16661_/X sky130_fd_sc_hd__buf_4
XFILLER_274_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13873_ _26071_/Q _13706_/A _14495_/A _13872_/X vssd1 vssd1 vccd1 vccd1 _13873_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25859_ _26938_/CLK _25859_/D vssd1 vssd1 vccd1 vccd1 _25859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_175_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25607_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18400_ _27042_/Q _18503_/A _18395_/X _18398_/X _18519_/A vssd1 vssd1 vccd1 vccd1
+ _18400_/X sky130_fd_sc_hd__o221a_1
X_15612_ _15581_/Y _15594_/Y _15611_/Y _14817_/A _13207_/A vssd1 vssd1 vccd1 vccd1
+ _15612_/Y sky130_fd_sc_hd__o221ai_4
X_12824_ _25482_/Q _25481_/Q _12953_/A vssd1 vssd1 vccd1 vccd1 _12866_/B sky130_fd_sc_hd__o21bai_2
XFILLER_262_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19380_ _19381_/A _19381_/B vssd1 vssd1 vccd1 vccd1 _19414_/B sky130_fd_sc_hd__and2_1
X_16592_ _17669_/A _17992_/A _17658_/A vssd1 vssd1 vccd1 vccd1 _18077_/B sky130_fd_sc_hd__o21a_1
XFILLER_262_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_104_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26322_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_216_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15543_ _15384_/S _15540_/X _15542_/X _14659_/A vssd1 vssd1 vccd1 vccd1 _15543_/X
+ sky130_fd_sc_hd__a211o_1
X_18331_ _18738_/A _18322_/X _18330_/X vssd1 vssd1 vccd1 vccd1 _18331_/X sky130_fd_sc_hd__a21o_1
XFILLER_203_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12755_ _12755_/A vssd1 vssd1 vccd1 vccd1 _12756_/A sky130_fd_sc_hd__buf_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ _18049_/X _18062_/X _18262_/S vssd1 vssd1 vccd1 vccd1 _18490_/B sky130_fd_sc_hd__mux2_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _27281_/Q _26474_/Q _15474_/S vssd1 vssd1 vccd1 vccd1 _15474_/X sky130_fd_sc_hd__mux2_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12810_/A vssd1 vssd1 vccd1 vccd1 _17971_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14425_ _12768_/A _26393_/Q _15888_/S _26909_/Q _13140_/A vssd1 vssd1 vccd1 vccd1
+ _14425_/X sky130_fd_sc_hd__o221a_1
X_17213_ _17222_/A _17213_/B vssd1 vssd1 vccd1 vccd1 _17214_/A sky130_fd_sc_hd__and2_1
XFILLER_175_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18193_ _19454_/A _18193_/B vssd1 vssd1 vccd1 vccd1 _18193_/Y sky130_fd_sc_hd__nor2_1
X_17144_ _25477_/Q vssd1 vssd1 vccd1 vccd1 _23363_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_190_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14356_ _14421_/A _14341_/X _14355_/X _13171_/A vssd1 vssd1 vccd1 vccd1 _14356_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13307_ _25584_/Q vssd1 vssd1 vccd1 vccd1 _13477_/A sky130_fd_sc_hd__inv_2
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17075_ _26238_/Q vssd1 vssd1 vccd1 vccd1 _22393_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_171_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14287_ _13664_/A _25832_/Q _26032_/Q _15775_/S _13337_/A vssd1 vssd1 vccd1 vccd1
+ _14287_/X sky130_fd_sc_hd__a221o_1
XFILLER_155_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16026_ _13512_/A _16024_/X _16025_/X _14077_/A vssd1 vssd1 vccd1 vccd1 _16026_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13238_ _13644_/A vssd1 vssd1 vccd1 vccd1 _13239_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_170_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13169_ _14621_/A _13128_/X _13145_/X _13165_/X _14681_/A vssd1 vssd1 vccd1 vccd1
+ _13169_/X sky130_fd_sc_hd__a311o_1
XFILLER_124_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17977_ _18271_/B _17974_/Y _18209_/S vssd1 vssd1 vccd1 vccd1 _17977_/X sky130_fd_sc_hd__mux2_1
XFILLER_266_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19716_ _20452_/A _19693_/X _19714_/Y _24986_/B vssd1 vssd1 vccd1 vccd1 _19716_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16928_ _16909_/X _16878_/B _16877_/X _16910_/X _16911_/X vssd1 vssd1 vccd1 vccd1
+ _16928_/X sky130_fd_sc_hd__o221a_1
XFILLER_111_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19647_ _20461_/S vssd1 vssd1 vccd1 vccd1 _19649_/A sky130_fd_sc_hd__buf_2
XFILLER_253_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16859_ _16859_/A vssd1 vssd1 vccd1 vccd1 _16860_/B sky130_fd_sc_hd__buf_4
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19578_ _19389_/X _19390_/Y _19425_/Y _17853_/X vssd1 vssd1 vccd1 vccd1 _19581_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18529_ _25731_/Q _18530_/B vssd1 vssd1 vccd1 vccd1 _18588_/C sky130_fd_sc_hd__and2_2
XFILLER_244_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21540_ _21540_/A vssd1 vssd1 vccd1 vccd1 _21540_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21471_ _21469_/X _21470_/X _21433_/X vssd1 vssd1 vccd1 vccd1 _21471_/X sky130_fd_sc_hd__a21o_1
XFILLER_140_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23210_ _23210_/A vssd1 vssd1 vccd1 vccd1 _26551_/D sky130_fd_sc_hd__clkbuf_1
X_20422_ _20443_/B _20443_/C _20406_/B vssd1 vssd1 vccd1 vccd1 _20427_/A sky130_fd_sc_hd__a21bo_1
X_24190_ _24239_/A vssd1 vssd1 vccd1 vccd1 _24216_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23141_ _23209_/S vssd1 vssd1 vccd1 vccd1 _23150_/S sky130_fd_sc_hd__buf_4
XFILLER_174_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20353_ _20353_/A _20353_/B vssd1 vssd1 vccd1 vccd1 _20399_/B sky130_fd_sc_hd__or2_1
XFILLER_106_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23072_ _23072_/A vssd1 vssd1 vccd1 vccd1 _26498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20284_ _20284_/A _20300_/D vssd1 vssd1 vccd1 vccd1 _20284_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_150_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22023_ _26123_/Q _20958_/X _22027_/S vssd1 vssd1 vccd1 vccd1 _22024_/A sky130_fd_sc_hd__mux2_1
X_26900_ _26900_/CLK _26900_/D vssd1 vssd1 vccd1 vccd1 _26900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26831_ _27314_/CLK _26831_/D vssd1 vssd1 vccd1 vccd1 _26831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_276_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26611_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_69_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26762_ _27309_/CLK _26762_/D vssd1 vssd1 vccd1 vccd1 _26762_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23974_ _26862_/Q _23568_/X _23976_/S vssd1 vssd1 vccd1 vccd1 _23975_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25713_ _26673_/CLK _25713_/D vssd1 vssd1 vccd1 vccd1 _25713_/Q sky130_fd_sc_hd__dfxtp_1
X_22925_ _22947_/A vssd1 vssd1 vccd1 vccd1 _22934_/S sky130_fd_sc_hd__buf_4
X_26693_ _26917_/CLK _26693_/D vssd1 vssd1 vccd1 vccd1 _26693_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25644_ _25661_/CLK _25644_/D vssd1 vssd1 vccd1 vccd1 _25644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22856_ _26408_/Q _22695_/X _22862_/S vssd1 vssd1 vccd1 vccd1 _22857_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21807_ _21864_/S vssd1 vssd1 vccd1 vccd1 _21816_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_231_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25575_ _25590_/CLK _25575_/D vssd1 vssd1 vccd1 vccd1 _25575_/Q sky130_fd_sc_hd__dfxtp_4
X_22787_ _26378_/Q _22701_/X _22789_/S vssd1 vssd1 vccd1 vccd1 _22788_/A sky130_fd_sc_hd__mux2_1
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27314_ _27314_/CLK _27314_/D vssd1 vssd1 vccd1 vccd1 _27314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24526_ _24361_/S _25627_/Q _24525_/X vssd1 vssd1 vccd1 vccd1 _24765_/B sky130_fd_sc_hd__o21a_4
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21738_ _21738_/A vssd1 vssd1 vccd1 vccd1 _26003_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27245_ _27309_/CLK _27245_/D vssd1 vssd1 vccd1 vccd1 _27245_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24457_ _24457_/A vssd1 vssd1 vccd1 vccd1 _24457_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_185_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21669_ _21669_/A vssd1 vssd1 vccd1 vccd1 _25974_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14210_ _13941_/X _14208_/X _14209_/X _13479_/A vssd1 vssd1 vccd1 vccd1 _14211_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23408_ _26639_/Q _23098_/X _23408_/S vssd1 vssd1 vccd1 vccd1 _23409_/A sky130_fd_sc_hd__mux2_1
X_15190_ _15164_/X _15189_/X _15071_/X vssd1 vssd1 vccd1 vccd1 _15190_/Y sky130_fd_sc_hd__a21oi_4
X_27176_ _27176_/CLK _27176_/D vssd1 vssd1 vccd1 vccd1 _27176_/Q sky130_fd_sc_hd__dfxtp_1
X_24388_ _24408_/A _24559_/A vssd1 vssd1 vccd1 vccd1 _24388_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14141_ _14485_/B _14936_/C _12869_/X vssd1 vssd1 vccd1 vccd1 _14141_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_138_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26127_ _26843_/CLK _26127_/D vssd1 vssd1 vccd1 vccd1 _26127_/Q sky130_fd_sc_hd__dfxtp_1
X_23339_ _23339_/A vssd1 vssd1 vccd1 vccd1 _26608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14072_ _14468_/A _14070_/X _14071_/X _14067_/X vssd1 vssd1 vccd1 vccd1 _14076_/B
+ sky130_fd_sc_hd__o211a_1
X_26058_ _26453_/CLK _26058_/D vssd1 vssd1 vccd1 vccd1 _26058_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13023_ _15825_/S _13862_/A vssd1 vssd1 vccd1 vccd1 _14713_/D sky130_fd_sc_hd__nor2_4
X_17900_ _17898_/X _17899_/X _17958_/S vssd1 vssd1 vccd1 vccd1 _17900_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25009_ _27167_/Q _25000_/X _25008_/X vssd1 vssd1 vccd1 vccd1 _27167_/D sky130_fd_sc_hd__o21ba_1
X_18880_ _18775_/X _18878_/Y _18382_/A vssd1 vssd1 vccd1 vccd1 _18880_/X sky130_fd_sc_hd__o21ba_1
XFILLER_266_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17831_ _17831_/A _16040_/B vssd1 vssd1 vccd1 vccd1 _18905_/A sky130_fd_sc_hd__or2b_1
XFILLER_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17762_ _17762_/A _17762_/B _17762_/C vssd1 vssd1 vccd1 vccd1 _18468_/A sky130_fd_sc_hd__or3_4
XFILLER_208_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14974_ _14650_/A _14969_/X _14973_/X _14679_/X vssd1 vssd1 vccd1 vccd1 _14974_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_208_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19501_ _25635_/Q _19510_/B vssd1 vssd1 vccd1 vccd1 _19501_/X sky130_fd_sc_hd__or2_1
XFILLER_47_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16713_ _16713_/A _16713_/B vssd1 vssd1 vccd1 vccd1 _16714_/B sky130_fd_sc_hd__nor2_2
X_13925_ _15954_/A _13925_/B vssd1 vssd1 vccd1 vccd1 _13925_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17693_ _17747_/B _17722_/B vssd1 vssd1 vccd1 vccd1 _17762_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19432_ _27229_/Q _19462_/B vssd1 vssd1 vccd1 vccd1 _19432_/X sky130_fd_sc_hd__and2_1
XFILLER_262_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13856_ _13085_/A _26399_/Q _13431_/A _13855_/X vssd1 vssd1 vccd1 vccd1 _13856_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_403 _17043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16644_ _16657_/A _17533_/A _13911_/X vssd1 vssd1 vccd1 vccd1 _16644_/X sky130_fd_sc_hd__a21o_1
XFILLER_228_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_414 _17009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_425 _12781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_436 _25728_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12807_ _13215_/A _25570_/Q vssd1 vssd1 vccd1 vccd1 _17504_/C sky130_fd_sc_hd__nand2_1
X_19363_ _17327_/X _18439_/A _18441_/A _25561_/Q vssd1 vssd1 vccd1 vccd1 _19363_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_447 _26940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_458 _25983_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13787_ _14725_/A _13787_/B _13787_/C vssd1 vssd1 vccd1 vccd1 _13787_/X sky130_fd_sc_hd__or3_1
X_16575_ _16575_/A _16575_/B _16575_/C _16575_/D vssd1 vssd1 vccd1 vccd1 _17055_/C
+ sky130_fd_sc_hd__or4_2
XINSDIODE2_469 _23699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18314_ _18314_/A vssd1 vssd1 vccd1 vccd1 _18321_/A sky130_fd_sc_hd__clkbuf_2
X_12738_ _25583_/Q _14076_/A _12738_/C _12738_/D vssd1 vssd1 vccd1 vccd1 _12738_/X
+ sky130_fd_sc_hd__and4b_4
X_15526_ _25742_/Q _20141_/A _15526_/S vssd1 vssd1 vccd1 vccd1 _15528_/B sky130_fd_sc_hd__mux2_2
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ _18643_/A _18734_/X _19294_/S vssd1 vssd1 vccd1 vccd1 _19294_/X sky130_fd_sc_hd__mux2_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18245_ _25504_/Q _18810_/A _18242_/X _18244_/X _18832_/A vssd1 vssd1 vccd1 vccd1
+ _18245_/X sky130_fd_sc_hd__o221a_1
X_15457_ _15559_/S _15456_/X _13071_/A vssd1 vssd1 vccd1 vccd1 _15457_/X sky130_fd_sc_hd__a21o_1
XFILLER_230_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14408_ _14594_/A _14406_/X _14407_/X vssd1 vssd1 vccd1 vccd1 _14447_/A sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_72_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26592_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18176_ _25503_/Q _18810_/A _18167_/X _18174_/X _18832_/A vssd1 vssd1 vccd1 vccd1
+ _18176_/X sky130_fd_sc_hd__o221a_1
X_15388_ _15388_/A vssd1 vssd1 vccd1 vccd1 _15388_/X sky130_fd_sc_hd__buf_4
XFILLER_237_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14339_ _14111_/A _14337_/X _14338_/X _14115_/S vssd1 vssd1 vccd1 vccd1 _14339_/X
+ sky130_fd_sc_hd__a211o_1
X_17127_ _17127_/A vssd1 vssd1 vccd1 vccd1 _25471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_274_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17058_ _16604_/A _16804_/Y _16996_/A vssd1 vssd1 vccd1 vccd1 _20796_/C sky130_fd_sc_hd__a21o_2
XFILLER_143_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16009_ _15490_/A _27275_/Q _26468_/Q _15858_/S _13966_/A vssd1 vssd1 vccd1 vccd1
+ _16009_/X sky130_fd_sc_hd__a221o_1
XFILLER_83_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20971_ _25860_/Q _20970_/X _20971_/S vssd1 vssd1 vccd1 vccd1 _20972_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22710_ _22710_/A vssd1 vssd1 vccd1 vccd1 _26348_/D sky130_fd_sc_hd__clkbuf_1
X_23690_ _23690_/A vssd1 vssd1 vccd1 vccd1 _23690_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_214_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22641_ _22817_/B _22641_/B _22817_/C vssd1 vssd1 vccd1 vccd1 _23291_/B sky130_fd_sc_hd__or3_4
XFILLER_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25360_ _25360_/A vssd1 vssd1 vccd1 vccd1 _27279_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22572_ _22567_/X _22571_/Y _22561_/X vssd1 vssd1 vccd1 vccd1 _26304_/D sky130_fd_sc_hd__a21oi_1
XFILLER_210_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24311_ _26995_/Q _24311_/B vssd1 vssd1 vccd1 vccd1 _24318_/C sky130_fd_sc_hd__and2_1
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21523_ _21509_/X _19139_/X _21510_/X _25818_/Q _21483_/X vssd1 vssd1 vccd1 vccd1
+ _21523_/X sky130_fd_sc_hd__a221o_1
XFILLER_22_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25291_ _23744_/X _27249_/Q _25293_/S vssd1 vssd1 vccd1 vccd1 _25292_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27030_ _27062_/CLK _27030_/D vssd1 vssd1 vccd1 vccd1 _27030_/Q sky130_fd_sc_hd__dfxtp_1
X_24242_ _26970_/Q _24237_/B _24241_/Y vssd1 vssd1 vccd1 vccd1 _26970_/D sky130_fd_sc_hd__o21a_1
XFILLER_119_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21454_ _25951_/Q _21443_/X _21453_/Y _21400_/X vssd1 vssd1 vccd1 vccd1 _25951_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_147_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20405_ _20426_/A _20405_/B vssd1 vssd1 vccd1 vccd1 _20406_/B sky130_fd_sc_hd__nand2_1
X_24173_ _24188_/A _24178_/C vssd1 vssd1 vccd1 vccd1 _24173_/Y sky130_fd_sc_hd__nor2_1
X_21385_ _21385_/A vssd1 vssd1 vccd1 vccd1 _21385_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23124_ _23597_/A vssd1 vssd1 vccd1 vccd1 _23124_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20336_ _19657_/X _20382_/C _20335_/Y _20100_/X vssd1 vssd1 vccd1 vccd1 _20337_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_190_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23055_ _26493_/Q _23053_/X _23067_/S vssd1 vssd1 vccd1 vccd1 _23056_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20267_ _27123_/Q _20248_/X _20112_/X _20266_/X vssd1 vssd1 vccd1 vccd1 _20267_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22006_ _22006_/A vssd1 vssd1 vccd1 vccd1 _26115_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_276_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput103 dout0[6] vssd1 vssd1 vccd1 vccd1 input103/X sky130_fd_sc_hd__clkbuf_2
XTAP_5325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput114 dout1[16] vssd1 vssd1 vccd1 vccd1 input114/X sky130_fd_sc_hd__clkbuf_1
X_20198_ _20379_/A _20299_/B vssd1 vssd1 vccd1 vccd1 _20305_/A sky130_fd_sc_hd__and2_1
XFILLER_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput125 dout1[26] vssd1 vssd1 vccd1 vccd1 input125/X sky130_fd_sc_hd__clkbuf_1
XTAP_5347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput136 dout1[36] vssd1 vssd1 vccd1 vccd1 input136/X sky130_fd_sc_hd__clkbuf_2
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput147 dout1[46] vssd1 vssd1 vccd1 vccd1 input147/X sky130_fd_sc_hd__clkbuf_2
X_26814_ _26878_/CLK _26814_/D vssd1 vssd1 vccd1 vccd1 _26814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput158 dout1[56] vssd1 vssd1 vccd1 vccd1 input158/X sky130_fd_sc_hd__clkbuf_2
XTAP_5369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput169 dout1[8] vssd1 vssd1 vccd1 vccd1 input169/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23957_ _26854_/Q _23542_/X _23965_/S vssd1 vssd1 vccd1 vccd1 _23958_/A sky130_fd_sc_hd__mux2_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26745_ _26905_/CLK _26745_/D vssd1 vssd1 vccd1 vccd1 _26745_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13710_ _13086_/X _26692_/Q _26820_/Q _16067_/S _13051_/A vssd1 vssd1 vccd1 vccd1
+ _13710_/X sky130_fd_sc_hd__a221o_1
XFILLER_16_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22908_ _26431_/Q _22666_/X _22912_/S vssd1 vssd1 vccd1 vccd1 _22909_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26676_ _26739_/CLK _26676_/D vssd1 vssd1 vccd1 vccd1 _26676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14690_ _12751_/A _14685_/X _14689_/X vssd1 vssd1 vccd1 vccd1 _14690_/X sky130_fd_sc_hd__o21a_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23888_ _23888_/A vssd1 vssd1 vccd1 vccd1 _26823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13641_ _13641_/A _13641_/B vssd1 vssd1 vccd1 vccd1 _14449_/B sky130_fd_sc_hd__nand2_4
X_22839_ _22839_/A vssd1 vssd1 vccd1 vccd1 _26400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25627_ _27327_/CLK _25627_/D vssd1 vssd1 vccd1 vccd1 _25627_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _16358_/X _16359_/X _16360_/S vssd1 vssd1 vccd1 vccd1 _16360_/X sky130_fd_sc_hd__mux2_1
X_25558_ _25992_/CLK _25558_/D vssd1 vssd1 vccd1 vccd1 _25558_/Q sky130_fd_sc_hd__dfxtp_2
X_13572_ _14031_/A _13572_/B vssd1 vssd1 vccd1 vccd1 _13573_/B sky130_fd_sc_hd__nor2_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _15311_/A vssd1 vssd1 vccd1 vccd1 _15312_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_185_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24509_ _24518_/A _24972_/A vssd1 vssd1 vccd1 vccd1 _24509_/Y sky130_fd_sc_hd__nand2_1
XFILLER_184_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _19156_/A _19156_/B _19191_/B _16290_/X vssd1 vssd1 vccd1 vccd1 _16572_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_9_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25489_ _26683_/CLK _25489_/D vssd1 vssd1 vccd1 vccd1 _25489_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_200_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18030_ _25725_/Q vssd1 vssd1 vccd1 vccd1 _20626_/A sky130_fd_sc_hd__buf_4
X_15242_ _25596_/Q _13636_/B _13179_/A vssd1 vssd1 vccd1 vccd1 _15243_/A sky130_fd_sc_hd__a21o_1
X_27228_ _27228_/CLK _27228_/D vssd1 vssd1 vccd1 vccd1 _27228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27159_ _27160_/CLK _27159_/D vssd1 vssd1 vccd1 vccd1 _27159_/Q sky130_fd_sc_hd__dfxtp_2
X_15173_ _26120_/Q _26021_/Q _16396_/S vssd1 vssd1 vccd1 vccd1 _15173_/X sky130_fd_sc_hd__mux2_1
X_14124_ _25590_/Q _14124_/B vssd1 vssd1 vccd1 vccd1 _14124_/X sky130_fd_sc_hd__or2_1
XFILLER_207_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19981_ _19981_/A _20081_/A vssd1 vssd1 vccd1 vccd1 _19982_/C sky130_fd_sc_hd__or2_1
XFILLER_67_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14055_ _25802_/Q _27236_/Q _14553_/S vssd1 vssd1 vccd1 vccd1 _14055_/X sky130_fd_sc_hd__mux2_1
X_18932_ _18968_/A _18932_/B vssd1 vssd1 vccd1 vccd1 _18932_/X sky130_fd_sc_hd__or2_1
XFILLER_97_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13006_ _20487_/C _13006_/B vssd1 vssd1 vccd1 vccd1 _13007_/A sky130_fd_sc_hd__or2_1
XFILLER_95_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18863_ _18861_/X _18862_/X _16628_/B vssd1 vssd1 vccd1 vccd1 _18864_/D sky130_fd_sc_hd__a21oi_1
XFILLER_239_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_190_wb_clk_i _26681_/CLK vssd1 vssd1 vccd1 vccd1 _27322_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17814_ _18325_/A _18325_/B _17800_/A _16714_/A _17813_/X vssd1 vssd1 vccd1 vccd1
+ _18539_/D sky130_fd_sc_hd__o2111a_1
X_18794_ _18794_/A _18794_/B vssd1 vssd1 vccd1 vccd1 _18795_/B sky130_fd_sc_hd__nand2_1
XTAP_5870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17745_ _17745_/A _17753_/A vssd1 vssd1 vccd1 vccd1 _18116_/B sky130_fd_sc_hd__nand2_2
XFILLER_130_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14957_ _14956_/A _14952_/X _14956_/Y _14706_/X vssd1 vssd1 vccd1 vccd1 _14957_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13908_ _17797_/B _13908_/B vssd1 vssd1 vccd1 vccd1 _13909_/B sky130_fd_sc_hd__nor2_1
XINSDIODE2_200 _14403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17676_ _17691_/A vssd1 vssd1 vccd1 vccd1 _17697_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14888_ _17852_/A vssd1 vssd1 vccd1 vccd1 _16458_/A sky130_fd_sc_hd__inv_2
XFILLER_63_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_211 _15192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19415_ _19421_/B _19415_/B vssd1 vssd1 vccd1 vccd1 _19415_/Y sky130_fd_sc_hd__nand2_2
XINSDIODE2_222 _20034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16627_ _18906_/A _16627_/B vssd1 vssd1 vccd1 vccd1 _16748_/A sky130_fd_sc_hd__xor2_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_233 _16407_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13839_ _13839_/A _13839_/B vssd1 vssd1 vccd1 vccd1 _13839_/Y sky130_fd_sc_hd__nor2_2
XINSDIODE2_244 _18483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_255 _16904_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_266 _20686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19346_ _25751_/Q _25750_/Q _19346_/C vssd1 vssd1 vccd1 vccd1 _19381_/B sky130_fd_sc_hd__and3_1
XINSDIODE2_277 _27107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_288 _25819_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16558_ _16558_/A _19392_/B vssd1 vssd1 vccd1 vccd1 _19388_/A sky130_fd_sc_hd__xnor2_4
XFILLER_188_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_299 _27271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15509_ _15509_/A _15509_/B vssd1 vssd1 vccd1 vccd1 _15509_/X sky130_fd_sc_hd__or2_1
XFILLER_188_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19277_ _19277_/A _19277_/B vssd1 vssd1 vccd1 vccd1 _19577_/A sky130_fd_sc_hd__xnor2_1
XFILLER_241_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16489_ _27326_/Q _26583_/Q _16493_/S vssd1 vssd1 vccd1 vccd1 _16489_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18228_ _19709_/A _18227_/C _25727_/Q vssd1 vssd1 vccd1 vccd1 _18229_/B sky130_fd_sc_hd__a21oi_1
XFILLER_191_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18159_ _27071_/Q _18391_/A _18292_/A _27169_/Q _18293_/A vssd1 vssd1 vccd1 vccd1
+ _18159_/X sky130_fd_sc_hd__a221o_1
XFILLER_117_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21170_ _21170_/A vssd1 vssd1 vccd1 vccd1 _25927_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20121_ _20280_/B _19002_/Y _19589_/B _20120_/X vssd1 vssd1 vccd1 vccd1 _20121_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20052_ _20052_/A vssd1 vssd1 vccd1 vccd1 _20052_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24860_ _27121_/Q _24873_/B vssd1 vssd1 vccd1 vccd1 _24860_/Y sky130_fd_sc_hd__nand2_1
XFILLER_274_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23811_ _23811_/A vssd1 vssd1 vccd1 vccd1 _26789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24791_ _24874_/A vssd1 vssd1 vccd1 vccd1 _24791_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26530_ _27309_/CLK _26530_/D vssd1 vssd1 vccd1 vccd1 _26530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23742_ _23741_/X _26765_/Q _23748_/S vssd1 vssd1 vccd1 vccd1 _23743_/A sky130_fd_sc_hd__mux2_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20954_ _20954_/A vssd1 vssd1 vccd1 vccd1 _25854_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26461_ _26462_/CLK _26461_/D vssd1 vssd1 vccd1 vccd1 _26461_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23673_ _23673_/A vssd1 vssd1 vccd1 vccd1 _26742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20885_ _25833_/Q _20884_/X _20885_/S vssd1 vssd1 vccd1 vccd1 _20886_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25412_ _25412_/A vssd1 vssd1 vccd1 vccd1 _27302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22624_ _26224_/Q _26223_/Q _26219_/Q vssd1 vssd1 vccd1 vccd1 _22624_/X sky130_fd_sc_hd__o21ba_1
X_26392_ _27266_/CLK _26392_/D vssd1 vssd1 vccd1 vccd1 _26392_/Q sky130_fd_sc_hd__dfxtp_2
X_25343_ _27272_/Q _23715_/A _25343_/S vssd1 vssd1 vccd1 vccd1 _25344_/A sky130_fd_sc_hd__mux2_1
X_22555_ _22607_/A vssd1 vssd1 vccd1 vccd1 _22565_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21506_ _21573_/A vssd1 vssd1 vccd1 vccd1 _21506_/X sky130_fd_sc_hd__clkbuf_2
X_25274_ _23718_/X _27241_/Q _25282_/S vssd1 vssd1 vccd1 vccd1 _25275_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22486_ _22486_/A vssd1 vssd1 vccd1 vccd1 _26268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27013_ _27049_/CLK _27013_/D vssd1 vssd1 vccd1 vccd1 _27013_/Q sky130_fd_sc_hd__dfxtp_1
X_24225_ _24237_/A _24225_/B vssd1 vssd1 vccd1 vccd1 _24225_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21437_ _21646_/S vssd1 vssd1 vccd1 vccd1 _21489_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_182_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24156_ _26942_/Q _24157_/C _24155_/Y vssd1 vssd1 vccd1 vccd1 _26942_/D sky130_fd_sc_hd__o21a_1
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21368_ _21363_/X _21366_/X _21367_/X vssd1 vssd1 vccd1 vccd1 _21368_/X sky130_fd_sc_hd__a21o_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23107_ _23107_/A vssd1 vssd1 vccd1 vccd1 _26509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20319_ _27157_/Q _27091_/Q vssd1 vssd1 vccd1 vccd1 _20339_/A sky130_fd_sc_hd__and2_1
XFILLER_123_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24087_ _26912_/Q _23523_/X _24087_/S vssd1 vssd1 vccd1 vccd1 _24088_/A sky130_fd_sc_hd__mux2_1
X_21299_ _25939_/Q _21202_/X _21298_/Y _21262_/X vssd1 vssd1 vccd1 vccd1 _25939_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_150_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23038_ _23137_/S vssd1 vssd1 vccd1 vccd1 _23051_/S sky130_fd_sc_hd__buf_6
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15860_ _15401_/A _15857_/X _15859_/X _13241_/A vssd1 vssd1 vccd1 vccd1 _15860_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_209_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_opt_11_0_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_53_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14811_ _27293_/Q _26486_/Q _14811_/S vssd1 vssd1 vccd1 vccd1 _14811_/X sky130_fd_sc_hd__mux2_1
XTAP_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _15791_/A _15954_/B _15791_/C vssd1 vssd1 vccd1 vccd1 _15791_/Y sky130_fd_sc_hd__nor3_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24989_ _24989_/A _24541_/B vssd1 vssd1 vccd1 vccd1 _24989_/X sky130_fd_sc_hd__or2b_1
XFILLER_18_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17530_ _25904_/Q _17517_/X _14321_/Y _17525_/X vssd1 vssd1 vccd1 vccd1 _17530_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_26728_ _26856_/CLK _26728_/D vssd1 vssd1 vccd1 vccd1 _26728_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14742_ _14742_/A vssd1 vssd1 vccd1 vccd1 _14743_/A sky130_fd_sc_hd__buf_2
XFILLER_83_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17461_ _17461_/A vssd1 vssd1 vccd1 vccd1 _21206_/A sky130_fd_sc_hd__buf_2
X_14673_ _27293_/Q _26486_/Q _16467_/A vssd1 vssd1 vccd1 vccd1 _14673_/X sky130_fd_sc_hd__mux2_1
X_26659_ _27303_/CLK _26659_/D vssd1 vssd1 vccd1 vccd1 _26659_/Q sky130_fd_sc_hd__dfxtp_1
X_19200_ _27124_/Q _19056_/X _19198_/X _19199_/X vssd1 vssd1 vccd1 vccd1 _19200_/X
+ sky130_fd_sc_hd__o22a_2
X_13624_ _25838_/Q _26038_/Q _15725_/S vssd1 vssd1 vccd1 vccd1 _13625_/B sky130_fd_sc_hd__mux2_1
X_16412_ _25625_/Q _14597_/X _16411_/X _14618_/X vssd1 vssd1 vccd1 vccd1 _23597_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17392_ _25549_/Q _17392_/B vssd1 vssd1 vccd1 vccd1 _17399_/C sky130_fd_sc_hd__and2_1
XFILLER_60_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19131_ _27090_/Q _19058_/X _19059_/X _27188_/Q _19060_/X vssd1 vssd1 vccd1 vccd1
+ _19131_/X sky130_fd_sc_hd__a221o_1
X_13555_ _12944_/X _12945_/X _12948_/Y vssd1 vssd1 vccd1 vccd1 _13556_/A sky130_fd_sc_hd__a21oi_1
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16343_ _26645_/Q _26741_/Q _16359_/S vssd1 vssd1 vccd1 vccd1 _16343_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16274_ _13255_/X _26707_/Q _26835_/Q _16347_/S _14770_/A vssd1 vssd1 vccd1 vccd1
+ _16274_/X sky130_fd_sc_hd__a221o_1
X_19062_ _27120_/Q _19056_/X _19057_/X _19061_/X vssd1 vssd1 vccd1 vccd1 _19062_/X
+ sky130_fd_sc_hd__o22a_2
X_13486_ _13829_/S vssd1 vssd1 vccd1 vccd1 _13792_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15225_ _26088_/Q _25893_/Q _16428_/S vssd1 vssd1 vccd1 vccd1 _15225_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18013_ _18285_/A vssd1 vssd1 vccd1 vccd1 _18013_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput407 _17019_/X vssd1 vssd1 vccd1 vccd1 din0[9] sky130_fd_sc_hd__buf_2
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15156_ _26512_/Q _26384_/Q _16395_/S vssd1 vssd1 vccd1 vccd1 _15156_/X sky130_fd_sc_hd__mux2_1
Xoutput418 _25953_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[17] sky130_fd_sc_hd__buf_2
Xoutput429 _25963_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[27] sky130_fd_sc_hd__buf_2
XFILLER_271_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14107_ _14107_/A vssd1 vssd1 vccd1 vccd1 _14107_/X sky130_fd_sc_hd__buf_2
XFILLER_141_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15087_ _14917_/X _15083_/X _15086_/X _14803_/A vssd1 vssd1 vccd1 vccd1 _15087_/X
+ sky130_fd_sc_hd__a211o_1
X_19964_ _19954_/Y _19955_/X _19962_/X _19963_/X _19651_/X vssd1 vssd1 vccd1 vccd1
+ _19964_/X sky130_fd_sc_hd__a221o_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14038_ _13911_/A _14489_/A _17545_/C _12902_/X _25907_/Q vssd1 vssd1 vccd1 vccd1
+ _14038_/X sky130_fd_sc_hd__o32a_1
X_18915_ _27084_/Q _19058_/A _19059_/A _27182_/Q _19060_/A vssd1 vssd1 vccd1 vccd1
+ _18915_/X sky130_fd_sc_hd__a221o_1
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19895_ _19896_/A _19896_/B vssd1 vssd1 vccd1 vccd1 _19895_/X sky130_fd_sc_hd__or2_1
XFILLER_68_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18846_ _18723_/X _18842_/X _18845_/X _18782_/X vssd1 vssd1 vccd1 vccd1 _18847_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_267_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18777_ _19076_/A vssd1 vssd1 vccd1 vccd1 _18777_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15989_ _26108_/Q _26009_/Q _15989_/S vssd1 vssd1 vccd1 vccd1 _15989_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17728_ _17750_/A _17728_/B vssd1 vssd1 vccd1 vccd1 _17730_/B sky130_fd_sc_hd__nor2_4
XFILLER_82_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17659_ _17553_/X _17658_/Y _22535_/B vssd1 vssd1 vccd1 vccd1 _25597_/D sky130_fd_sc_hd__a21o_1
XFILLER_24_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20670_ _20670_/A _20670_/B vssd1 vssd1 vccd1 vccd1 _20670_/X sky130_fd_sc_hd__or2_1
XFILLER_149_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19329_ _19323_/X _19324_/X _19328_/X _18636_/X vssd1 vssd1 vccd1 vccd1 _19329_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_259_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22340_ _17087_/C _26225_/Q _22340_/S vssd1 vssd1 vccd1 vccd1 _22340_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22271_ _22271_/A vssd1 vssd1 vccd1 vccd1 _22271_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24010_ _24010_/A vssd1 vssd1 vccd1 vccd1 _26877_/D sky130_fd_sc_hd__clkbuf_1
X_21222_ _21217_/X _21220_/X _21289_/A vssd1 vssd1 vccd1 vccd1 _21222_/X sky130_fd_sc_hd__a21o_1
XFILLER_145_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21153_ _25923_/Q _21148_/X _21149_/X input23/X vssd1 vssd1 vccd1 vccd1 _21154_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_105_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20104_ _27149_/Q _27083_/Q vssd1 vssd1 vccd1 vccd1 _20131_/A sky130_fd_sc_hd__and2_1
X_25961_ _26995_/CLK _25961_/D vssd1 vssd1 vccd1 vccd1 _25961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21084_ _21138_/A vssd1 vssd1 vccd1 vccd1 _21100_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_259_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24912_ _24941_/A vssd1 vssd1 vccd1 vccd1 _24957_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_20035_ _20194_/B _18883_/Y _19911_/A _20034_/X vssd1 vssd1 vccd1 vccd1 _20035_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_246_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25892_ _27287_/CLK _25892_/D vssd1 vssd1 vccd1 vccd1 _25892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24843_ _24841_/Y _24842_/X _24835_/X vssd1 vssd1 vccd1 vccd1 _27116_/D sky130_fd_sc_hd__a21oi_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24774_ _24771_/X _24636_/A _24772_/Y _24773_/X vssd1 vssd1 vccd1 vccd1 _24774_/X
+ sky130_fd_sc_hd__a31o_1
X_21986_ _26106_/Q _20903_/X _21994_/S vssd1 vssd1 vccd1 vccd1 _21987_/A sky130_fd_sc_hd__mux2_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23725_ _23725_/A vssd1 vssd1 vccd1 vccd1 _23725_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_242_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26513_ _27288_/CLK _26513_/D vssd1 vssd1 vccd1 vccd1 _26513_/Q sky130_fd_sc_hd__dfxtp_1
X_20937_ _25849_/Q _20935_/X _20949_/S vssd1 vssd1 vccd1 vccd1 _20938_/A sky130_fd_sc_hd__mux2_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26444_ _27283_/CLK _26444_/D vssd1 vssd1 vccd1 vccd1 _26444_/Q sky130_fd_sc_hd__dfxtp_1
X_23656_ _26735_/Q _23571_/X _23656_/S vssd1 vssd1 vccd1 vccd1 _23657_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20868_ _20868_/A _20868_/B _21888_/C vssd1 vssd1 vccd1 vccd1 _25321_/A sky130_fd_sc_hd__or3_4
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22607_ _22607_/A vssd1 vssd1 vccd1 vccd1 _22618_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_230_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26375_ _27278_/CLK _26375_/D vssd1 vssd1 vccd1 vccd1 _26375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23587_ _23587_/A vssd1 vssd1 vccd1 vccd1 _23587_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20799_ _21709_/A _20799_/B vssd1 vssd1 vccd1 vccd1 _25795_/D sky130_fd_sc_hd__nor2_1
X_25326_ _27264_/Q _23690_/A _25332_/S vssd1 vssd1 vccd1 vccd1 _25327_/A sky130_fd_sc_hd__mux2_1
X_13340_ _13340_/A vssd1 vssd1 vccd1 vccd1 _14751_/A sky130_fd_sc_hd__buf_4
XFILLER_183_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22538_ _22567_/A vssd1 vssd1 vccd1 vccd1 _22538_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25257_ _25257_/A vssd1 vssd1 vccd1 vccd1 _27233_/D sky130_fd_sc_hd__clkbuf_1
X_13271_ _13976_/A vssd1 vssd1 vccd1 vccd1 _14228_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_154_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22469_ _26211_/Q _22459_/X _22467_/X _22468_/X vssd1 vssd1 vccd1 vccd1 _26259_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_129_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27154_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15010_ _14987_/Y _14994_/Y _14790_/X _15009_/Y vssd1 vssd1 vccd1 vccd1 _15010_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24208_ _24208_/A vssd1 vssd1 vccd1 vccd1 _24938_/A sky130_fd_sc_hd__buf_4
XFILLER_154_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25188_ _24664_/B _25172_/X _25187_/X _27204_/Q _25179_/X vssd1 vssd1 vccd1 vccd1
+ _27204_/D sky130_fd_sc_hd__o221a_1
XFILLER_118_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24139_ _24139_/A vssd1 vssd1 vccd1 vccd1 _26935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16961_ _16414_/Y _16952_/X _16834_/A vssd1 vssd1 vccd1 vccd1 _16965_/B sky130_fd_sc_hd__o21ai_2
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18700_ _17375_/X _18459_/X _18699_/X _18154_/A _18466_/X vssd1 vssd1 vccd1 vccd1
+ _18700_/X sky130_fd_sc_hd__a221o_1
XFILLER_77_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15912_ _25578_/Q _15948_/B _15243_/A _15911_/X vssd1 vssd1 vccd1 vccd1 _17829_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_1_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19680_ _19642_/X _19645_/X _19649_/Y _19651_/X _19679_/X vssd1 vssd1 vccd1 vccd1
+ _19680_/X sky130_fd_sc_hd__a311o_2
X_16892_ _16887_/X _16889_/X _16891_/X vssd1 vssd1 vccd1 vccd1 _16893_/B sky130_fd_sc_hd__a21boi_4
XFILLER_204_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18631_ _18631_/A vssd1 vssd1 vccd1 vccd1 _25607_/D sky130_fd_sc_hd__clkbuf_1
X_15843_ _15843_/A _15843_/B vssd1 vssd1 vccd1 vccd1 _15843_/X sky130_fd_sc_hd__or2_1
XFILLER_209_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18562_ _27109_/Q _18504_/X _18560_/X _18561_/X vssd1 vssd1 vccd1 vccd1 _18562_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_218_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15774_ _27310_/Q _26567_/Q _15931_/S vssd1 vssd1 vccd1 vccd1 _15774_/X sky130_fd_sc_hd__mux2_1
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _13993_/A vssd1 vssd1 vccd1 vccd1 _14518_/S sky130_fd_sc_hd__buf_4
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17513_ _12803_/X _17662_/B _17503_/X _18027_/A _17512_/X vssd1 vssd1 vccd1 vccd1
+ _17513_/X sky130_fd_sc_hd__o311a_1
XFILLER_233_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ _14725_/A vssd1 vssd1 vccd1 vccd1 _16439_/A sky130_fd_sc_hd__buf_8
XFILLER_73_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ _18492_/A _18489_/X _18492_/Y _18799_/A vssd1 vssd1 vccd1 vccd1 _18493_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17444_ _17444_/A _17697_/B _17444_/C _17444_/D vssd1 vssd1 vccd1 vccd1 _19570_/D
+ sky130_fd_sc_hd__or4_2
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14656_ _15026_/B vssd1 vssd1 vccd1 vccd1 _16501_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13607_ _13164_/A _13588_/X _13595_/X _13606_/X vssd1 vssd1 vccd1 vccd1 _13607_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_177_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17375_ _25544_/Q vssd1 vssd1 vccd1 vccd1 _17375_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_220_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14587_ _15659_/A vssd1 vssd1 vccd1 vccd1 _16170_/A sky130_fd_sc_hd__buf_2
XFILLER_159_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19114_ _18841_/X _19088_/Y _19103_/X _19113_/Y _18375_/X vssd1 vssd1 vccd1 vccd1
+ _19114_/X sky130_fd_sc_hd__a32o_1
X_16326_ _15065_/A _26709_/Q _26837_/Q _16399_/S _15048_/A vssd1 vssd1 vccd1 vccd1
+ _16326_/X sky130_fd_sc_hd__a221o_1
X_13538_ _15488_/A _26598_/Q _15841_/S _26338_/Q _13834_/A vssd1 vssd1 vccd1 vccd1
+ _13538_/X sky130_fd_sc_hd__o221a_1
XFILLER_229_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19045_ _19045_/A _19045_/B vssd1 vssd1 vccd1 vccd1 _19045_/Y sky130_fd_sc_hd__xnor2_4
X_13469_ _14535_/A vssd1 vssd1 vccd1 vccd1 _14725_/A sky130_fd_sc_hd__buf_6
X_16257_ _14742_/A _26415_/Q _15308_/S _16256_/X vssd1 vssd1 vccd1 vccd1 _16257_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15208_ _15203_/X _15204_/X _16442_/S vssd1 vssd1 vccd1 vccd1 _15208_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16188_ _13242_/X _16186_/X _16187_/X _14801_/A vssd1 vssd1 vccd1 vccd1 _16188_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15139_ _23587_/A vssd1 vssd1 vccd1 vccd1 _15139_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19947_ _19947_/A _20055_/B vssd1 vssd1 vccd1 vccd1 _19947_/X sky130_fd_sc_hd__or2_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19878_ _25669_/Q _19906_/C vssd1 vssd1 vccd1 vccd1 _19878_/X sky130_fd_sc_hd__xor2_1
XFILLER_229_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18829_ _18829_/A vssd1 vssd1 vccd1 vccd1 _18829_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21840_ _21851_/A vssd1 vssd1 vccd1 vccd1 _21849_/S sky130_fd_sc_hd__buf_4
XFILLER_208_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21771_ _21771_/A vssd1 vssd1 vccd1 vccd1 _26018_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_270_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23510_ _23591_/A vssd1 vssd1 vccd1 vccd1 _23610_/S sky130_fd_sc_hd__buf_4
X_20722_ _20496_/X _25759_/Q _20728_/S vssd1 vssd1 vccd1 vccd1 _20723_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24490_ _26315_/Q _24393_/X _24394_/X input229/X _24457_/X vssd1 vssd1 vccd1 vccd1
+ _24490_/X sky130_fd_sc_hd__a221o_1
XFILLER_223_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23441_ _26653_/Q _23041_/X _23447_/S vssd1 vssd1 vccd1 vccd1 _23442_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20653_ _26272_/Q _20646_/X _20652_/X _20644_/X vssd1 vssd1 vccd1 vccd1 _25735_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26160_ _27264_/CLK _26160_/D vssd1 vssd1 vccd1 vccd1 _26160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23372_ _23372_/A vssd1 vssd1 vccd1 vccd1 _26622_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20584_ _23757_/A vssd1 vssd1 vccd1 vccd1 _20584_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25111_ _27186_/Q _25085_/X _25110_/X vssd1 vssd1 vccd1 vccd1 _27186_/D sky130_fd_sc_hd__o21ba_1
X_22323_ _26219_/Q _22310_/X _22316_/X _26320_/Q _22317_/X vssd1 vssd1 vccd1 vccd1
+ _22323_/X sky130_fd_sc_hd__a221o_1
XFILLER_99_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26091_ _27257_/CLK _26091_/D vssd1 vssd1 vccd1 vccd1 _26091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25042_ _27173_/Q _25030_/X _25041_/X vssd1 vssd1 vccd1 vccd1 _27173_/D sky130_fd_sc_hd__o21ba_1
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22254_ _22269_/A vssd1 vssd1 vccd1 vccd1 _22254_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21205_ _24501_/A vssd1 vssd1 vccd1 vccd1 _21885_/A sky130_fd_sc_hd__buf_2
XFILLER_145_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22185_ _22200_/A vssd1 vssd1 vccd1 vccd1 _22185_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21136_ _21136_/A _21136_/B vssd1 vssd1 vccd1 vccd1 _21137_/A sky130_fd_sc_hd__or2_1
XFILLER_278_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26993_ _27001_/CLK _26993_/D vssd1 vssd1 vccd1 vccd1 _26993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25944_ _27022_/CLK _25944_/D vssd1 vssd1 vccd1 vccd1 _25944_/Q sky130_fd_sc_hd__dfxtp_1
X_21067_ input42/X _21195_/A _20487_/B vssd1 vssd1 vccd1 vccd1 _21174_/A sky130_fd_sc_hd__a21o_4
XFILLER_246_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20018_ _25672_/Q _20017_/C _22498_/A vssd1 vssd1 vccd1 vccd1 _20018_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_219_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25875_ _26465_/CLK _25875_/D vssd1 vssd1 vccd1 vccd1 _25875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12840_ _25868_/Q vssd1 vssd1 vccd1 vccd1 _13741_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_62_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24826_ _20652_/A _24810_/X _24690_/Y _24811_/X vssd1 vssd1 vccd1 vccd1 _24826_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12771_/A vssd1 vssd1 vccd1 vccd1 _12772_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21969_ _21969_/A vssd1 vssd1 vccd1 vccd1 _26098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24757_ _24764_/A _24757_/B vssd1 vssd1 vccd1 vccd1 _27095_/D sky130_fd_sc_hd__nor2_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14510_ _26780_/Q _26424_/Q _14518_/S vssd1 vssd1 vccd1 vccd1 _14510_/X sky130_fd_sc_hd__mux2_1
XFILLER_215_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15490_/A vssd1 vssd1 vccd1 vccd1 _15491_/A sky130_fd_sc_hd__clkbuf_2
X_23708_ _23708_/A vssd1 vssd1 vccd1 vccd1 _26754_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24688_ _24699_/A _24688_/B vssd1 vssd1 vccd1 vccd1 _27079_/D sky130_fd_sc_hd__nor2_1
XFILLER_214_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26427_ _27267_/CLK _26427_/D vssd1 vssd1 vccd1 vccd1 _26427_/Q sky130_fd_sc_hd__dfxtp_2
X_14441_ _14424_/X _14427_/X _14440_/X _14523_/A vssd1 vssd1 vccd1 vccd1 _14441_/X
+ sky130_fd_sc_hd__a22o_1
X_23639_ _26727_/Q _23546_/X _23645_/S vssd1 vssd1 vccd1 vccd1 _23640_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14372_ _27297_/Q _26554_/Q _14391_/S vssd1 vssd1 vccd1 vccd1 _14372_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17160_ _25465_/S vssd1 vssd1 vccd1 vccd1 _20707_/C sky130_fd_sc_hd__buf_6
XFILLER_128_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26358_ _27293_/CLK _26358_/D vssd1 vssd1 vccd1 vccd1 _26358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16111_ _16111_/A _16111_/B vssd1 vssd1 vccd1 vccd1 _16111_/X sky130_fd_sc_hd__or2_1
XFILLER_10_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ _15322_/A vssd1 vssd1 vccd1 vccd1 _16189_/S sky130_fd_sc_hd__buf_6
X_25309_ _23770_/X _27257_/Q _25315_/S vssd1 vssd1 vccd1 vccd1 _25310_/A sky130_fd_sc_hd__mux2_1
X_17091_ _26236_/Q _17091_/B _17091_/C vssd1 vssd1 vccd1 vccd1 _22210_/A sky130_fd_sc_hd__or3_2
X_26289_ _26292_/CLK _26289_/D vssd1 vssd1 vccd1 vccd1 _26289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13254_ _13254_/A vssd1 vssd1 vccd1 vccd1 _13255_/A sky130_fd_sc_hd__buf_2
X_16042_ _18906_/A _16627_/B _18901_/S vssd1 vssd1 vccd1 vccd1 _16626_/B sky130_fd_sc_hd__a21oi_4
XFILLER_143_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13185_ _13185_/A _25584_/Q vssd1 vssd1 vccd1 vccd1 _13209_/A sky130_fd_sc_hd__nand2_1
XFILLER_135_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_123_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19801_ _19824_/B _18434_/Y _19663_/X _19800_/X vssd1 vssd1 vccd1 vccd1 _19801_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_124_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17993_ _18214_/A vssd1 vssd1 vccd1 vccd1 _18861_/A sky130_fd_sc_hd__buf_2
XFILLER_123_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19732_ _19776_/A _19776_/B vssd1 vssd1 vccd1 vccd1 _19853_/A sky130_fd_sc_hd__xnor2_1
X_16944_ _16944_/A vssd1 vssd1 vccd1 vccd1 _16944_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_97_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27297_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19663_ _19670_/A vssd1 vssd1 vccd1 vccd1 _19663_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_26_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27326_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16875_ _16893_/A _16875_/B vssd1 vssd1 vccd1 vccd1 _16876_/A sky130_fd_sc_hd__and2_1
XFILLER_92_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18614_ _27142_/Q vssd1 vssd1 vccd1 vccd1 _19896_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15826_ _15824_/X _15825_/X _15826_/S vssd1 vssd1 vccd1 vccd1 _15826_/X sky130_fd_sc_hd__mux2_1
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19594_ _19594_/A _19911_/A vssd1 vssd1 vccd1 vccd1 _20189_/B sky130_fd_sc_hd__nand2_2
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18545_ _17961_/B _17915_/X _18729_/A vssd1 vssd1 vccd1 vccd1 _18546_/A sky130_fd_sc_hd__mux2_1
XFILLER_252_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15757_ _15606_/X _15755_/X _15756_/X _14228_/X vssd1 vssd1 vccd1 vccd1 _15757_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12969_ _12866_/A _12866_/B _12961_/A _21429_/A _21630_/A vssd1 vssd1 vccd1 vccd1
+ _12969_/Y sky130_fd_sc_hd__a221oi_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14708_ _14708_/A vssd1 vssd1 vccd1 vccd1 _14709_/A sky130_fd_sc_hd__clkbuf_4
X_18476_ _18891_/A _18434_/Y _18473_/X _18475_/X _18005_/A vssd1 vssd1 vccd1 vccd1
+ _18476_/X sky130_fd_sc_hd__a221o_1
XFILLER_233_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15688_ _25813_/Q _27247_/Q _15914_/S vssd1 vssd1 vccd1 vccd1 _15689_/B sky130_fd_sc_hd__mux2_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17427_ _17427_/A _25560_/Q _17427_/C vssd1 vssd1 vccd1 vccd1 _17434_/C sky130_fd_sc_hd__and3_1
XFILLER_178_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14639_ _14870_/A vssd1 vssd1 vccd1 vccd1 _16324_/S sky130_fd_sc_hd__buf_4
XFILLER_14_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17358_ _17356_/X _17360_/C _17357_/Y vssd1 vssd1 vccd1 vccd1 _25538_/D sky130_fd_sc_hd__o21a_1
XFILLER_158_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16309_ _27288_/Q _26481_/Q _16315_/S vssd1 vssd1 vccd1 vccd1 _16309_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17289_ _17287_/X _17293_/C _17288_/Y vssd1 vssd1 vccd1 vccd1 _25517_/D sky130_fd_sc_hd__o21a_1
XFILLER_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19028_ _25551_/Q _18825_/X _19027_/X _18829_/X _18830_/X vssd1 vssd1 vccd1 vccd1
+ _19028_/X sky130_fd_sc_hd__a221o_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23990_ _26869_/Q _23590_/X _23998_/S vssd1 vssd1 vccd1 vccd1 _23991_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22941_ _26446_/Q _22714_/X _22945_/S vssd1 vssd1 vccd1 vccd1 _22942_/A sky130_fd_sc_hd__mux2_1
XFILLER_284_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25660_ _25660_/CLK _25660_/D vssd1 vssd1 vccd1 vccd1 _25660_/Q sky130_fd_sc_hd__dfxtp_1
X_22872_ _22872_/A vssd1 vssd1 vccd1 vccd1 _26415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_283_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21823_ _26041_/Q _20910_/X _21827_/S vssd1 vssd1 vccd1 vccd1 _21824_/A sky130_fd_sc_hd__mux2_1
X_24611_ _24611_/A _24621_/B vssd1 vssd1 vccd1 vccd1 _24611_/Y sky130_fd_sc_hd__nand2_1
XFILLER_243_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25591_ _25596_/CLK _25591_/D vssd1 vssd1 vccd1 vccd1 _25591_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27330_ _27330_/A vssd1 vssd1 vccd1 vccd1 _27330_/X sky130_fd_sc_hd__buf_2
X_24542_ _24542_/A _24542_/B vssd1 vssd1 vccd1 vccd1 _24543_/B sky130_fd_sc_hd__or2_1
X_21754_ _20550_/X _26011_/Q _21754_/S vssd1 vssd1 vccd1 vccd1 _21755_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20705_ _25756_/Q _22130_/A vssd1 vssd1 vccd1 vccd1 _20706_/A sky130_fd_sc_hd__and2_1
XFILLER_212_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24473_ _24473_/A vssd1 vssd1 vccd1 vccd1 _24473_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27261_ _27326_/CLK _27261_/D vssd1 vssd1 vccd1 vccd1 _27261_/Q sky130_fd_sc_hd__dfxtp_1
X_21685_ _25982_/Q input194/X _21685_/S vssd1 vssd1 vccd1 vccd1 _21686_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26212_ _26322_/CLK _26212_/D vssd1 vssd1 vccd1 vccd1 _26212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23424_ _26646_/Q _23121_/X _23430_/S vssd1 vssd1 vccd1 vccd1 _23425_/A sky130_fd_sc_hd__mux2_1
X_20636_ _26265_/Q _20633_/X _20635_/X _20631_/X vssd1 vssd1 vccd1 vccd1 _25728_/D
+ sky130_fd_sc_hd__o211a_1
X_27192_ _27198_/CLK _27192_/D vssd1 vssd1 vccd1 vccd1 _27192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26143_ _26531_/CLK _26143_/D vssd1 vssd1 vccd1 vccd1 _26143_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_165_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23355_ _20609_/X _26616_/Q _23357_/S vssd1 vssd1 vccd1 vccd1 _23356_/A sky130_fd_sc_hd__mux2_1
X_20567_ _23744_/A vssd1 vssd1 vccd1 vccd1 _20567_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_166_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22306_ _26213_/Q _22294_/X _22300_/X _26314_/Q _22301_/X vssd1 vssd1 vccd1 vccd1
+ _22306_/X sky130_fd_sc_hd__a221o_1
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26074_ _27277_/CLK _26074_/D vssd1 vssd1 vccd1 vccd1 _26074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23286_ _23286_/A vssd1 vssd1 vccd1 vccd1 _26585_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20498_ _20498_/A vssd1 vssd1 vccd1 vccd1 _25693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25025_ _22478_/A _25015_/X _25004_/X _18329_/A _25024_/X vssd1 vssd1 vccd1 vccd1
+ _25025_/X sky130_fd_sc_hd__a221o_1
X_22237_ _22630_/B vssd1 vssd1 vccd1 vccd1 _22270_/A sky130_fd_sc_hd__buf_2
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22168_ _26174_/Q _22152_/X _22167_/X _22164_/X vssd1 vssd1 vccd1 vccd1 _26174_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21119_ _21119_/A vssd1 vssd1 vccd1 vccd1 _25913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26976_ _26980_/CLK _26976_/D vssd1 vssd1 vccd1 vccd1 _26976_/Q sky130_fd_sc_hd__dfxtp_1
X_22099_ _26157_/Q _20964_/X _22099_/S vssd1 vssd1 vccd1 vccd1 _22100_/A sky130_fd_sc_hd__mux2_1
X_14990_ _14766_/A _14988_/X _14989_/X _12757_/A vssd1 vssd1 vccd1 vccd1 _14990_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_75_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13941_ _13941_/A vssd1 vssd1 vccd1 vccd1 _13941_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25927_ _27213_/CLK _25927_/D vssd1 vssd1 vccd1 vccd1 _25927_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16660_ _16660_/A _20973_/B vssd1 vssd1 vccd1 vccd1 _16661_/A sky130_fd_sc_hd__or2b_2
X_13872_ _25876_/Q _14273_/B vssd1 vssd1 vccd1 vccd1 _13872_/X sky130_fd_sc_hd__or2_1
X_25858_ _26453_/CLK _25858_/D vssd1 vssd1 vccd1 vccd1 _25858_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_262_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15611_ _15598_/X _15601_/X _15610_/Y vssd1 vssd1 vccd1 vccd1 _15611_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_62_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12823_ _12953_/A _25480_/Q vssd1 vssd1 vccd1 vccd1 _12866_/A sky130_fd_sc_hd__or2b_1
X_24809_ _27108_/Q _24818_/B vssd1 vssd1 vccd1 vccd1 _24809_/Y sky130_fd_sc_hd__nand2_1
X_16591_ _16591_/A _17162_/A vssd1 vssd1 vccd1 vccd1 _17971_/D sky130_fd_sc_hd__or2_4
X_25789_ _27326_/CLK _25789_/D vssd1 vssd1 vccd1 vccd1 _25789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18330_ _18942_/B _18328_/X _18329_/Y _18358_/A vssd1 vssd1 vccd1 vccd1 _18330_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15542_ _25814_/Q _15255_/A _16059_/S _15541_/X vssd1 vssd1 vccd1 vccd1 _15542_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12754_ _12754_/A vssd1 vssd1 vccd1 vccd1 _12755_/A sky130_fd_sc_hd__buf_6
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18261_ _18063_/X _18059_/C _18262_/S vssd1 vssd1 vccd1 vccd1 _18261_/X sky130_fd_sc_hd__mux2_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15473_ _15471_/X _15472_/X _15473_/S vssd1 vssd1 vccd1 vccd1 _15473_/X sky130_fd_sc_hd__mux2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _25568_/Q _17500_/B _18028_/B vssd1 vssd1 vccd1 vccd1 _12810_/A sky130_fd_sc_hd__or3b_4
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_144_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25796_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17212_ _25496_/Q _17529_/A _17146_/A _17443_/B vssd1 vssd1 vccd1 vccd1 _17213_/B
+ sky130_fd_sc_hd__a22o_1
X_14424_ _25798_/Q _14713_/D _14423_/X _15727_/S vssd1 vssd1 vccd1 vccd1 _14424_/X
+ sky130_fd_sc_hd__a211o_1
X_18192_ _18898_/A _18799_/B _18191_/X vssd1 vssd1 vccd1 vccd1 _18193_/B sky130_fd_sc_hd__a21bo_1
XFILLER_128_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17143_ _17143_/A vssd1 vssd1 vccd1 vccd1 _25476_/D sky130_fd_sc_hd__clkbuf_1
X_14355_ _14355_/A _14355_/B vssd1 vssd1 vccd1 vccd1 _14355_/X sky130_fd_sc_hd__and2_1
XFILLER_156_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13306_ _16342_/S _13300_/X _13301_/X _13467_/A vssd1 vssd1 vccd1 vccd1 _13306_/X
+ sky130_fd_sc_hd__a31o_1
X_17074_ _26239_/Q vssd1 vssd1 vccd1 vccd1 _22361_/B sky130_fd_sc_hd__clkbuf_1
X_14286_ _26783_/Q _26427_/Q _14296_/S vssd1 vssd1 vccd1 vccd1 _14286_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16025_ _13835_/A _26856_/Q _25770_/Q _15515_/S _16022_/A vssd1 vssd1 vccd1 vccd1
+ _16025_/X sky130_fd_sc_hd__a221o_1
X_13237_ _13336_/A vssd1 vssd1 vccd1 vccd1 _13644_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13168_ _13168_/A vssd1 vssd1 vccd1 vccd1 _14681_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_170_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13099_ _14107_/A vssd1 vssd1 vccd1 vccd1 _14010_/S sky130_fd_sc_hd__buf_2
X_17976_ _18254_/A vssd1 vssd1 vccd1 vccd1 _18209_/S sky130_fd_sc_hd__buf_2
XFILLER_85_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19715_ _20236_/A vssd1 vssd1 vccd1 vccd1 _24986_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_66_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16927_ _16927_/A _16927_/B vssd1 vssd1 vccd1 vccd1 _16978_/C sky130_fd_sc_hd__nor2_1
XFILLER_226_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19646_ _19646_/A vssd1 vssd1 vccd1 vccd1 _20461_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_281_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16858_ _16858_/A vssd1 vssd1 vccd1 vccd1 _16858_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15809_ _26078_/Q _15797_/B _13134_/A _15808_/X vssd1 vssd1 vccd1 vccd1 _15809_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19577_ _19577_/A _19577_/B _19577_/C _19576_/X vssd1 vssd1 vccd1 vccd1 _19581_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_81_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16789_ _18035_/A vssd1 vssd1 vccd1 vccd1 _16938_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18528_ _18474_/A _18526_/X _18382_/X vssd1 vssd1 vccd1 vccd1 _18528_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18459_ _18459_/A vssd1 vssd1 vccd1 vccd1 _18459_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_222_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21470_ _21430_/X _18995_/X _21431_/X _25814_/Q _21403_/X vssd1 vssd1 vccd1 vccd1
+ _21470_/X sky130_fd_sc_hd__a221o_1
XFILLER_14_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20421_ _22531_/A _20396_/X _19780_/X vssd1 vssd1 vccd1 vccd1 _20421_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23140_ _23196_/A vssd1 vssd1 vccd1 vccd1 _23209_/S sky130_fd_sc_hd__buf_6
X_20352_ _20352_/A _20352_/B vssd1 vssd1 vccd1 vccd1 _20352_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23071_ _26498_/Q _23069_/X _23083_/S vssd1 vssd1 vccd1 vccd1 _23072_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20283_ _20299_/A _20283_/B vssd1 vssd1 vccd1 vccd1 _20300_/D sky130_fd_sc_hd__xnor2_1
XFILLER_115_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22022_ _22022_/A vssd1 vssd1 vccd1 vccd1 _26122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_276_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26830_ _27249_/CLK _26830_/D vssd1 vssd1 vccd1 vccd1 _26830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_275_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26761_ _27304_/CLK _26761_/D vssd1 vssd1 vccd1 vccd1 _26761_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23973_ _23973_/A vssd1 vssd1 vccd1 vccd1 _26861_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25712_ _27283_/CLK _25712_/D vssd1 vssd1 vccd1 vccd1 _25712_/Q sky130_fd_sc_hd__dfxtp_1
X_22924_ _22924_/A vssd1 vssd1 vccd1 vccd1 _26438_/D sky130_fd_sc_hd__clkbuf_1
X_26692_ _26916_/CLK _26692_/D vssd1 vssd1 vccd1 vccd1 _26692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25643_ _26813_/CLK _25643_/D vssd1 vssd1 vccd1 vccd1 _25643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22855_ _22855_/A vssd1 vssd1 vccd1 vccd1 _26407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21806_ _21806_/A vssd1 vssd1 vccd1 vccd1 _26033_/D sky130_fd_sc_hd__clkbuf_1
X_22786_ _22786_/A vssd1 vssd1 vccd1 vccd1 _26377_/D sky130_fd_sc_hd__clkbuf_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25574_ _25590_/CLK _25574_/D vssd1 vssd1 vccd1 vccd1 _25574_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27313_ _27313_/CLK _27313_/D vssd1 vssd1 vccd1 vccd1 _27313_/Q sky130_fd_sc_hd__dfxtp_1
X_21737_ _20517_/X _26003_/Q _21743_/S vssd1 vssd1 vccd1 vccd1 _21738_/A sky130_fd_sc_hd__mux2_1
X_24525_ _26322_/Q _21881_/X _21883_/X input236/X _24501_/X vssd1 vssd1 vccd1 vccd1
+ _24525_/X sky130_fd_sc_hd__a221o_2
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27244_ _27308_/CLK _27244_/D vssd1 vssd1 vccd1 vccd1 _27244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24456_ _24456_/A vssd1 vssd1 vccd1 vccd1 _24456_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_21668_ _25974_/Q input209/X _21674_/S vssd1 vssd1 vccd1 vccd1 _21669_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23407_ _23407_/A vssd1 vssd1 vccd1 vccd1 _26638_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20619_ _20619_/A vssd1 vssd1 vccd1 vccd1 _25722_/D sky130_fd_sc_hd__clkbuf_1
X_24387_ _24659_/B vssd1 vssd1 vccd1 vccd1 _24559_/A sky130_fd_sc_hd__inv_2
X_27175_ _27198_/CLK _27175_/D vssd1 vssd1 vccd1 vccd1 _27175_/Q sky130_fd_sc_hd__dfxtp_1
X_21599_ _25495_/Q _21620_/B vssd1 vssd1 vccd1 vccd1 _21599_/X sky130_fd_sc_hd__or2_1
X_14140_ _13911_/A _13561_/A _14139_/X _14029_/B _25930_/Q vssd1 vssd1 vccd1 vccd1
+ _14936_/C sky130_fd_sc_hd__o32a_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23338_ _20575_/X _26608_/Q _23346_/S vssd1 vssd1 vccd1 vccd1 _23339_/A sky130_fd_sc_hd__mux2_1
X_26126_ _27259_/CLK _26126_/D vssd1 vssd1 vccd1 vccd1 _26126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14071_ _14453_/A _26881_/Q _26753_/Q _13657_/A _14384_/A vssd1 vssd1 vccd1 vccd1
+ _14071_/X sky130_fd_sc_hd__a221o_1
X_26057_ _26453_/CLK _26057_/D vssd1 vssd1 vccd1 vccd1 _26057_/Q sky130_fd_sc_hd__dfxtp_2
X_23269_ _26577_/Q _23117_/X _23277_/S vssd1 vssd1 vccd1 vccd1 _23270_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13022_ _13022_/A vssd1 vssd1 vccd1 vccd1 _13862_/A sky130_fd_sc_hd__clkbuf_4
X_25008_ _24781_/Y _25137_/A _25007_/Y _24773_/X vssd1 vssd1 vccd1 vccd1 _25008_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_279_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17830_ _18838_/A _18794_/A _18855_/B vssd1 vssd1 vccd1 vccd1 _17830_/X sky130_fd_sc_hd__o21a_1
XFILLER_117_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17761_ _17742_/Y _17744_/X _17760_/X vssd1 vssd1 vccd1 vccd1 _17761_/X sky130_fd_sc_hd__o21a_2
X_26959_ _26992_/CLK _26959_/D vssd1 vssd1 vccd1 vccd1 _26959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_282_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14973_ _14693_/S _14970_/X _14972_/X _14662_/A vssd1 vssd1 vccd1 vccd1 _14973_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_282_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19500_ _19568_/B vssd1 vssd1 vccd1 vccd1 _19510_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_75_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16712_ _18324_/A _18324_/B vssd1 vssd1 vccd1 vccd1 _16714_/A sky130_fd_sc_hd__or2_2
XFILLER_235_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13924_ _13928_/A _13921_/Y _13922_/Y _13923_/X vssd1 vssd1 vccd1 vccd1 _13925_/B
+ sky130_fd_sc_hd__a211o_2
X_17692_ _17704_/S _25590_/Q _16481_/A _17691_/X vssd1 vssd1 vccd1 vccd1 _17722_/B
+ sky130_fd_sc_hd__o31ai_4
XFILLER_212_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19431_ _25531_/Q _18743_/X _18744_/X _25563_/Q vssd1 vssd1 vccd1 vccd1 _19431_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16643_ _25794_/Q vssd1 vssd1 vccd1 vccd1 _17533_/A sky130_fd_sc_hd__inv_2
XFILLER_263_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13855_ _26915_/Q _14001_/B vssd1 vssd1 vccd1 vccd1 _13855_/X sky130_fd_sc_hd__or2_1
XINSDIODE2_404 _17043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_415 _17009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_426 _12781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_437 _25729_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19362_ _19354_/Y _19357_/X _19358_/Y _19361_/X vssd1 vssd1 vccd1 vccd1 _19362_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12806_ _14358_/B vssd1 vssd1 vccd1 vccd1 _18076_/B sky130_fd_sc_hd__buf_2
X_16574_ _16776_/A _16773_/A vssd1 vssd1 vccd1 vccd1 _16575_/D sky130_fd_sc_hd__or2_2
XINSDIODE2_448 _26940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13786_ _13485_/X _13784_/X _13785_/X _12754_/A vssd1 vssd1 vccd1 vccd1 _13787_/C
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_459 _25984_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18313_ _18602_/A vssd1 vssd1 vccd1 vccd1 _18936_/A sky130_fd_sc_hd__clkbuf_2
X_15525_ _19031_/A vssd1 vssd1 vccd1 vccd1 _20141_/A sky130_fd_sc_hd__inv_2
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _13664_/A vssd1 vssd1 vccd1 vccd1 _12738_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19293_ _19423_/B _19577_/B _18183_/X vssd1 vssd1 vccd1 vccd1 _19293_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_163_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _25536_/Q _18825_/A _18243_/X _18829_/A _18830_/A vssd1 vssd1 vccd1 vccd1
+ _18244_/X sky130_fd_sc_hd__a221o_1
XFILLER_124_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15456_ _13694_/A _26894_/Q _26766_/Q _15630_/A vssd1 vssd1 vccd1 vccd1 _15456_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14407_ _14407_/A vssd1 vssd1 vccd1 vccd1 _14407_/X sky130_fd_sc_hd__buf_6
X_18175_ _18468_/A vssd1 vssd1 vccd1 vccd1 _18832_/A sky130_fd_sc_hd__clkbuf_2
X_15387_ _15370_/X _15386_/X _14591_/A vssd1 vssd1 vccd1 vccd1 _15387_/X sky130_fd_sc_hd__a21o_2
XFILLER_129_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17126_ _17137_/A _17126_/B vssd1 vssd1 vccd1 vccd1 _17127_/A sky130_fd_sc_hd__and2_1
X_14338_ _25585_/Q _26490_/Q _26362_/Q _14109_/B _13139_/A vssd1 vssd1 vccd1 vccd1
+ _14338_/X sky130_fd_sc_hd__o221a_1
XFILLER_156_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17057_ _26586_/Q _17003_/X _20794_/C _17051_/X vssd1 vssd1 vccd1 vccd1 _17057_/X
+ sky130_fd_sc_hd__a22o_4
X_14269_ _26523_/Q _26131_/Q _14269_/S vssd1 vssd1 vccd1 vccd1 _14269_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16008_ _15490_/A _26340_/Q _26600_/Q _15858_/S _16006_/A vssd1 vssd1 vccd1 vccd1
+ _16008_/X sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27312_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ _17955_/X _17958_/X _18050_/S vssd1 vssd1 vccd1 vccd1 _17959_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20970_ _23785_/A vssd1 vssd1 vccd1 vccd1 _20970_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19629_ _25173_/A vssd1 vssd1 vccd1 vccd1 _25218_/A sky130_fd_sc_hd__clkinv_4
XFILLER_53_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22640_ _23684_/A vssd1 vssd1 vccd1 vccd1 _22640_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_198_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22571_ _26304_/Q _22578_/B vssd1 vssd1 vccd1 vccd1 _22571_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24310_ _24327_/A _24310_/B _24311_/B vssd1 vssd1 vccd1 vccd1 _26994_/D sky130_fd_sc_hd__nor3_1
X_21522_ _25489_/Q _21574_/B vssd1 vssd1 vccd1 vccd1 _21522_/X sky130_fd_sc_hd__or2_1
X_25290_ _25290_/A vssd1 vssd1 vccd1 vccd1 _27248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24241_ _24269_/A _24243_/B vssd1 vssd1 vccd1 vccd1 _24241_/Y sky130_fd_sc_hd__nor2_1
XFILLER_210_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21453_ _21448_/Y _21452_/X _21425_/X vssd1 vssd1 vccd1 vccd1 _21453_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_108_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20404_ _20426_/A _20405_/B vssd1 vssd1 vccd1 vccd1 _20406_/A sky130_fd_sc_hd__or2_1
X_24172_ _26948_/Q _24175_/C vssd1 vssd1 vccd1 vccd1 _24178_/C sky130_fd_sc_hd__and2_1
X_21384_ input44/X input79/X _21422_/S vssd1 vssd1 vccd1 vccd1 _21385_/A sky130_fd_sc_hd__mux2_8
X_23123_ _23123_/A vssd1 vssd1 vccd1 vccd1 _26514_/D sky130_fd_sc_hd__clkbuf_1
X_20335_ _25684_/Q _20334_/C _22524_/A vssd1 vssd1 vccd1 vccd1 _20335_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23054_ _23137_/S vssd1 vssd1 vccd1 vccd1 _23067_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_122_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20266_ _19740_/X _20262_/Y _20265_/X _20067_/A vssd1 vssd1 vccd1 vccd1 _20266_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_115_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22005_ _26115_/Q _20932_/X _22005_/S vssd1 vssd1 vccd1 vccd1 _22006_/A sky130_fd_sc_hd__mux2_1
XFILLER_277_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput104 dout0[7] vssd1 vssd1 vccd1 vccd1 input104/X sky130_fd_sc_hd__clkbuf_2
XTAP_5326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20197_ _20426_/A _20299_/B vssd1 vssd1 vccd1 vccd1 _20199_/A sky130_fd_sc_hd__nor2_1
XFILLER_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput115 dout1[17] vssd1 vssd1 vccd1 vccd1 input115/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput126 dout1[27] vssd1 vssd1 vccd1 vccd1 input126/X sky130_fd_sc_hd__clkbuf_1
XFILLER_277_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput137 dout1[37] vssd1 vssd1 vccd1 vccd1 input137/X sky130_fd_sc_hd__clkbuf_2
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26813_ _26813_/CLK _26813_/D vssd1 vssd1 vccd1 vccd1 _26813_/Q sky130_fd_sc_hd__dfxtp_1
Xinput148 dout1[47] vssd1 vssd1 vccd1 vccd1 input148/X sky130_fd_sc_hd__clkbuf_2
XTAP_5359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput159 dout1[57] vssd1 vssd1 vccd1 vccd1 input159/X sky130_fd_sc_hd__clkbuf_2
XFILLER_276_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26744_ _26744_/CLK _26744_/D vssd1 vssd1 vccd1 vccd1 _26744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23956_ _24002_/S vssd1 vssd1 vccd1 vccd1 _23965_/S sky130_fd_sc_hd__buf_6
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22907_ _22907_/A vssd1 vssd1 vccd1 vccd1 _26430_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_272_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26675_ _27329_/A _26675_/D vssd1 vssd1 vccd1 vccd1 _26675_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23887_ _23722_/X _26823_/Q _23893_/S vssd1 vssd1 vccd1 vccd1 _23888_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13640_ _25580_/Q vssd1 vssd1 vccd1 vccd1 _13641_/B sky130_fd_sc_hd__buf_8
XFILLER_72_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25626_ _27327_/CLK _25626_/D vssd1 vssd1 vccd1 vccd1 _25626_/Q sky130_fd_sc_hd__dfxtp_4
X_22838_ _26400_/Q _22669_/X _22840_/S vssd1 vssd1 vccd1 vccd1 _22839_/A sky130_fd_sc_hd__mux2_1
XFILLER_260_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25557_ _25992_/CLK _25557_/D vssd1 vssd1 vccd1 vccd1 _25557_/Q sky130_fd_sc_hd__dfxtp_1
X_13571_ input170/X input142/X _14402_/S vssd1 vssd1 vccd1 vccd1 _13572_/B sky130_fd_sc_hd__mux2_8
XFILLER_25_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22769_ _22815_/S vssd1 vssd1 vccd1 vccd1 _22778_/S sky130_fd_sc_hd__buf_2
XFILLER_188_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15310_ _16185_/A _15310_/B vssd1 vssd1 vccd1 vccd1 _15310_/X sky130_fd_sc_hd__or2_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24508_ _24454_/X _25623_/Q _24507_/X vssd1 vssd1 vccd1 vccd1 _24972_/A sky130_fd_sc_hd__o21ai_4
XFILLER_158_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16290_ _16288_/A _19158_/S _16288_/B vssd1 vssd1 vccd1 vccd1 _16290_/X sky130_fd_sc_hd__o21ba_1
XFILLER_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25488_ _26683_/CLK _25488_/D vssd1 vssd1 vccd1 vccd1 _25488_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27227_ _27227_/CLK _27227_/D vssd1 vssd1 vccd1 vccd1 _27227_/Q sky130_fd_sc_hd__dfxtp_1
X_15241_ _17846_/B vssd1 vssd1 vccd1 vccd1 _19237_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_24439_ _24696_/B vssd1 vssd1 vccd1 vccd1 _24585_/A sky130_fd_sc_hd__clkinv_2
XFILLER_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27158_ _27160_/CLK _27158_/D vssd1 vssd1 vccd1 vccd1 _27158_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_138_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15172_ _26544_/Q _26152_/Q _16396_/S vssd1 vssd1 vccd1 vccd1 _15172_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26109_ _26468_/CLK _26109_/D vssd1 vssd1 vccd1 vccd1 _26109_/Q sky130_fd_sc_hd__dfxtp_4
X_14123_ _13008_/A _23526_/A _14122_/X _13026_/A vssd1 vssd1 vccd1 vccd1 _16827_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_67_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19980_ _19980_/A _19980_/B _19980_/C _19951_/C vssd1 vssd1 vccd1 vccd1 _20081_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_125_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27089_ _27213_/CLK _27089_/D vssd1 vssd1 vccd1 vccd1 _27089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18931_ _18967_/A _18931_/B vssd1 vssd1 vccd1 vccd1 _18931_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14054_ _14054_/A vssd1 vssd1 vccd1 vccd1 _14553_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_4_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13005_ _13005_/A _13005_/B _13005_/C vssd1 vssd1 vccd1 vccd1 _13006_/B sky130_fd_sc_hd__or3_1
XFILLER_239_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18862_ _18368_/A _18371_/A _18862_/S vssd1 vssd1 vccd1 vccd1 _18862_/X sky130_fd_sc_hd__mux2_1
XFILLER_234_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17813_ _17813_/A _17813_/B vssd1 vssd1 vccd1 vccd1 _17813_/X sky130_fd_sc_hd__and2_1
XFILLER_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18793_ _18724_/A _18724_/B _18726_/A vssd1 vssd1 vccd1 vccd1 _18794_/B sky130_fd_sc_hd__o21bai_1
XTAP_5860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17744_ _27133_/Q _27037_/Q _18952_/B vssd1 vssd1 vccd1 vccd1 _17744_/X sky130_fd_sc_hd__mux2_1
XTAP_5893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14956_ _14956_/A _14956_/B vssd1 vssd1 vccd1 vccd1 _14956_/Y sky130_fd_sc_hd__nand2_1
XFILLER_235_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13907_ _17797_/B _13908_/B vssd1 vssd1 vccd1 vccd1 _18498_/S sky130_fd_sc_hd__and2_1
X_17675_ _17708_/A vssd1 vssd1 vccd1 vccd1 _17691_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14887_ _19887_/A _18785_/A _14718_/X _14886_/X vssd1 vssd1 vccd1 vccd1 _17852_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_236_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_201 _14480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19414_ _25753_/Q _19414_/B vssd1 vssd1 vccd1 vccd1 _19415_/B sky130_fd_sc_hd__or2_1
XFILLER_62_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_212 _16916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16626_ _18941_/A _16626_/B vssd1 vssd1 vccd1 vccd1 _16751_/A sky130_fd_sc_hd__xnor2_4
XINSDIODE2_223 _20034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13838_ _15205_/A _13836_/X _13837_/X _13366_/A vssd1 vssd1 vccd1 vccd1 _13839_/B
+ sky130_fd_sc_hd__a31o_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_234 _16517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_245 _18541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_256 _16914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19345_ _18895_/X _19329_/X _19344_/X _19078_/X vssd1 vssd1 vccd1 vccd1 _19345_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_267 _24277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16557_ _16557_/A vssd1 vssd1 vccd1 vccd1 _19392_/B sky130_fd_sc_hd__buf_2
XINSDIODE2_278 _27327_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13769_ _25805_/Q _27239_/Q _13829_/S vssd1 vssd1 vccd1 vccd1 _13769_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_289 _25819_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15508_ _26538_/Q _26146_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15509_/B sky130_fd_sc_hd__mux2_1
XFILLER_241_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19276_ _19276_/A _19276_/B vssd1 vssd1 vccd1 vccd1 _19277_/B sky130_fd_sc_hd__nand2_1
X_16488_ _12722_/B _16476_/X _16481_/X _16487_/Y _17195_/A vssd1 vssd1 vccd1 vccd1
+ _16488_/X sky130_fd_sc_hd__a221o_1
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18227_ _25727_/Q _19709_/A _18227_/C vssd1 vssd1 vccd1 vccd1 _18287_/B sky130_fd_sc_hd__and3_1
X_15439_ _15439_/A _15439_/B vssd1 vssd1 vccd1 vccd1 _19109_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18158_ _18443_/A vssd1 vssd1 vccd1 vccd1 _18810_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17109_ _17137_/A _17109_/B vssd1 vssd1 vccd1 vccd1 _17110_/A sky130_fd_sc_hd__and2_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18089_ _20034_/B vssd1 vssd1 vccd1 vccd1 _20280_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20120_ _20120_/A _20227_/B vssd1 vssd1 vccd1 vccd1 _20120_/X sky130_fd_sc_hd__or2_1
XFILLER_259_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20051_ _19993_/X _20048_/X _20049_/Y _20050_/Y vssd1 vssd1 vccd1 vccd1 _20051_/X
+ sky130_fd_sc_hd__o31a_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23810_ _23715_/X _26789_/Q _23810_/S vssd1 vssd1 vccd1 vccd1 _23811_/A sky130_fd_sc_hd__mux2_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24790_ _24801_/A vssd1 vssd1 vccd1 vccd1 _24874_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23741_ _23741_/A vssd1 vssd1 vccd1 vccd1 _23741_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20953_ _25854_/Q _20951_/X _20965_/S vssd1 vssd1 vccd1 vccd1 _20954_/A sky130_fd_sc_hd__mux2_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26460_ _27267_/CLK _26460_/D vssd1 vssd1 vccd1 vccd1 _26460_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ _23699_/A vssd1 vssd1 vccd1 vccd1 _20884_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_23672_ _26742_/Q _23594_/X _23678_/S vssd1 vssd1 vccd1 vccd1 _23673_/A sky130_fd_sc_hd__mux2_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25411_ _23709_/X _27302_/Q _25415_/S vssd1 vssd1 vccd1 vccd1 _25412_/A sky130_fd_sc_hd__mux2_1
X_22623_ _22567_/A _22622_/Y _22614_/X vssd1 vssd1 vccd1 vccd1 _26324_/D sky130_fd_sc_hd__a21oi_1
X_26391_ _26917_/CLK _26391_/D vssd1 vssd1 vccd1 vccd1 _26391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22554_ _22554_/A vssd1 vssd1 vccd1 vccd1 _22607_/A sky130_fd_sc_hd__clkbuf_2
X_25342_ _25342_/A vssd1 vssd1 vccd1 vccd1 _27271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21505_ _25955_/Q _21443_/X _21504_/Y _21467_/X vssd1 vssd1 vccd1 vccd1 _25955_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_10_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25273_ _25319_/S vssd1 vssd1 vccd1 vccd1 _25282_/S sky130_fd_sc_hd__buf_6
X_22485_ _22485_/A _22491_/B vssd1 vssd1 vccd1 vccd1 _22486_/A sky130_fd_sc_hd__and2_1
XFILLER_148_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27012_ _27044_/CLK _27012_/D vssd1 vssd1 vccd1 vccd1 _27012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24224_ _26965_/Q _24227_/C vssd1 vssd1 vccd1 vccd1 _24225_/B sky130_fd_sc_hd__and2_1
XFILLER_194_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21436_ _21414_/X _21435_/X _21407_/X vssd1 vssd1 vccd1 vccd1 _21436_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_181_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24155_ _24164_/A _24160_/C vssd1 vssd1 vccd1 vccd1 _24155_/Y sky130_fd_sc_hd__nor2_1
XFILLER_181_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21367_ _21589_/A vssd1 vssd1 vccd1 vccd1 _21367_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_257_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20318_ _27125_/Q _20248_/X _20276_/X _20317_/X vssd1 vssd1 vccd1 vccd1 _20318_/X
+ sky130_fd_sc_hd__o211a_1
X_23106_ _26509_/Q _23105_/X _23115_/S vssd1 vssd1 vccd1 vccd1 _23107_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24086_ _24086_/A vssd1 vssd1 vccd1 vccd1 _26911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21298_ _21293_/Y _21295_/Y _21297_/X vssd1 vssd1 vccd1 vccd1 _21298_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_122_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23037_ _23118_/A vssd1 vssd1 vccd1 vccd1 _23137_/S sky130_fd_sc_hd__clkbuf_8
X_20249_ _20249_/A _20249_/B vssd1 vssd1 vccd1 vccd1 _20277_/A sky130_fd_sc_hd__nand2_2
XFILLER_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14810_ _26094_/Q _25899_/Q _14813_/S vssd1 vssd1 vccd1 vccd1 _14810_/X sky130_fd_sc_hd__mux2_1
XTAP_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _12913_/A _13925_/B _12929_/X vssd1 vssd1 vccd1 vccd1 _15790_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24988_ _25208_/A vssd1 vssd1 vccd1 vccd1 _24988_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_218_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26727_ _27306_/CLK _26727_/D vssd1 vssd1 vccd1 vccd1 _26727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14741_ _14741_/A vssd1 vssd1 vccd1 vccd1 _14742_/A sky130_fd_sc_hd__buf_2
X_23939_ _26846_/Q _23517_/X _23943_/S vssd1 vssd1 vccd1 vccd1 _23940_/A sky130_fd_sc_hd__mux2_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ _17460_/A vssd1 vssd1 vccd1 vccd1 _17461_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26658_ _27301_/CLK _26658_/D vssd1 vssd1 vccd1 vccd1 _26658_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14672_ _14670_/X _14671_/X _14700_/S vssd1 vssd1 vccd1 vccd1 _14672_/X sky130_fd_sc_hd__mux2_1
XFILLER_260_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16411_ _14601_/X _16409_/Y _16410_/X vssd1 vssd1 vccd1 vccd1 _16411_/X sky130_fd_sc_hd__o21a_1
XFILLER_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13623_ _15826_/S _13623_/B vssd1 vssd1 vccd1 vccd1 _13623_/X sky130_fd_sc_hd__or2_1
XFILLER_26_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25609_ _25725_/CLK _25609_/D vssd1 vssd1 vccd1 vccd1 _25609_/Q sky130_fd_sc_hd__dfxtp_4
X_17391_ _24966_/A vssd1 vssd1 vccd1 vccd1 _17430_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_260_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26589_ _26909_/CLK _26589_/D vssd1 vssd1 vccd1 vccd1 _26589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19130_ _27220_/Q _19331_/B vssd1 vssd1 vccd1 vccd1 _19130_/X sky130_fd_sc_hd__and2_1
XFILLER_9_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16342_ _16340_/X _16341_/X _16342_/S vssd1 vssd1 vccd1 vccd1 _16342_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13554_ _13554_/A vssd1 vssd1 vccd1 vccd1 _16735_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19061_ _27088_/Q _19058_/X _19059_/X _27186_/Q _19060_/X vssd1 vssd1 vccd1 vccd1
+ _19061_/X sky130_fd_sc_hd__a221o_1
X_16273_ _26643_/Q _26739_/Q _16273_/S vssd1 vssd1 vccd1 vccd1 _16273_/X sky130_fd_sc_hd__mux2_1
X_13485_ _13791_/A vssd1 vssd1 vccd1 vccd1 _13485_/X sky130_fd_sc_hd__buf_2
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18012_ _19218_/A _19253_/A vssd1 vssd1 vccd1 vccd1 _18285_/A sky130_fd_sc_hd__nor2_1
X_15224_ _15085_/X _15221_/X _15223_/X _14793_/A vssd1 vssd1 vccd1 vccd1 _15224_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_166_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput408 _17099_/X vssd1 vssd1 vccd1 vccd1 jtag_tdo sky130_fd_sc_hd__buf_2
X_15155_ _26352_/Q _26612_/Q _16395_/S vssd1 vssd1 vccd1 vccd1 _15155_/X sky130_fd_sc_hd__mux2_1
Xoutput419 _25954_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[18] sky130_fd_sc_hd__buf_2
XFILLER_126_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14106_ _13409_/A _14102_/X _14105_/X _13862_/A vssd1 vssd1 vccd1 vccd1 _14106_/X
+ sky130_fd_sc_hd__a211o_1
X_15086_ _26090_/Q _14891_/A _15084_/X _15085_/X vssd1 vssd1 vccd1 vccd1 _15086_/X
+ sky130_fd_sc_hd__o211a_1
X_19963_ _24848_/A vssd1 vssd1 vccd1 vccd1 _19963_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14037_ input162/X input137/X _14488_/S vssd1 vssd1 vccd1 vccd1 _17545_/C sky130_fd_sc_hd__mux2_8
X_18914_ _27214_/Q _18949_/B vssd1 vssd1 vccd1 vccd1 _18914_/X sky130_fd_sc_hd__and2_1
X_19894_ _20712_/A vssd1 vssd1 vccd1 vccd1 _19894_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18845_ _18892_/C _18844_/X vssd1 vssd1 vccd1 vccd1 _18845_/X sky130_fd_sc_hd__or2b_2
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18776_ _18775_/X _18773_/X _18705_/X vssd1 vssd1 vccd1 vccd1 _18776_/X sky130_fd_sc_hd__o21ba_1
XTAP_5690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15988_ _26532_/Q _26140_/Q _15988_/S vssd1 vssd1 vccd1 vccd1 _15988_/X sky130_fd_sc_hd__mux2_1
XFILLER_227_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17727_ _17730_/A _17732_/B vssd1 vssd1 vccd1 vccd1 _18458_/A sky130_fd_sc_hd__and2_1
XFILLER_36_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14939_ _14601_/X _14937_/Y _14938_/X vssd1 vssd1 vccd1 vccd1 _14939_/X sky130_fd_sc_hd__o21a_1
XFILLER_209_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17658_ _17658_/A _20687_/B vssd1 vssd1 vccd1 vccd1 _17658_/Y sky130_fd_sc_hd__nand2_2
XFILLER_235_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16609_ _16612_/A _16612_/B vssd1 vssd1 vccd1 vccd1 _16613_/A sky130_fd_sc_hd__or2_1
XFILLER_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17589_ _25916_/Q _17568_/X _13928_/B _17577_/X vssd1 vssd1 vccd1 vccd1 _17589_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_189_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19328_ _19327_/X _16566_/A _19328_/S vssd1 vssd1 vccd1 vccd1 _19328_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19259_ _27094_/Q _18508_/X _18509_/X _27192_/Q _18510_/X vssd1 vssd1 vccd1 vccd1
+ _19259_/X sky130_fd_sc_hd__a221o_1
XFILLER_192_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22270_ _22270_/A vssd1 vssd1 vccd1 vccd1 _22270_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21221_ _21221_/A _21221_/B vssd1 vssd1 vccd1 vccd1 _21289_/A sky130_fd_sc_hd__nor2_1
XFILLER_172_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21152_ _21152_/A vssd1 vssd1 vccd1 vccd1 _25922_/D sky130_fd_sc_hd__clkbuf_1
X_20103_ _27117_/Q _20079_/X _19967_/X _20102_/Y vssd1 vssd1 vccd1 vccd1 _20103_/X
+ sky130_fd_sc_hd__o211a_1
X_25960_ _26995_/CLK _25960_/D vssd1 vssd1 vccd1 vccd1 _25960_/Q sky130_fd_sc_hd__dfxtp_1
X_21083_ _21083_/A vssd1 vssd1 vccd1 vccd1 _25903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24911_ _27135_/Q _24902_/X _24910_/Y vssd1 vssd1 vccd1 vccd1 _27135_/D sky130_fd_sc_hd__o21a_1
X_20034_ _20034_/A _20034_/B vssd1 vssd1 vccd1 vccd1 _20034_/X sky130_fd_sc_hd__and2_1
X_25891_ _26611_/CLK _25891_/D vssd1 vssd1 vccd1 vccd1 _25891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24842_ _20664_/A _24829_/X _24707_/Y _24830_/X vssd1 vssd1 vccd1 vccd1 _24842_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_58_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24773_ _25027_/A vssd1 vssd1 vccd1 vccd1 _24773_/X sky130_fd_sc_hd__clkbuf_2
X_21985_ _22031_/S vssd1 vssd1 vccd1 vccd1 _21994_/S sky130_fd_sc_hd__buf_2
XFILLER_268_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26512_ _26739_/CLK _26512_/D vssd1 vssd1 vccd1 vccd1 _26512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23724_ _23724_/A vssd1 vssd1 vccd1 vccd1 _26759_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ _20952_/A vssd1 vssd1 vccd1 vccd1 _20949_/S sky130_fd_sc_hd__buf_4
XFILLER_270_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_8_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_8_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26443_ _26796_/CLK _26443_/D vssd1 vssd1 vccd1 vccd1 _26443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23655_ _23655_/A vssd1 vssd1 vccd1 vccd1 _26734_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20867_ _22817_/A _23363_/A _23363_/B vssd1 vssd1 vccd1 vccd1 _23788_/A sky130_fd_sc_hd__or3_4
XFILLER_41_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22606_ _22606_/A vssd1 vssd1 vccd1 vccd1 _22606_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26374_ _26467_/CLK _26374_/D vssd1 vssd1 vccd1 vccd1 _26374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23586_ _23586_/A vssd1 vssd1 vccd1 vccd1 _26707_/D sky130_fd_sc_hd__clkbuf_1
X_20798_ _21709_/A _20798_/B vssd1 vssd1 vccd1 vccd1 _25794_/D sky130_fd_sc_hd__nor2_1
XFILLER_139_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25325_ _25325_/A vssd1 vssd1 vccd1 vccd1 _27263_/D sky130_fd_sc_hd__clkbuf_1
X_22537_ _22606_/A vssd1 vssd1 vccd1 vccd1 _22567_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25256_ _23693_/X _27233_/Q _25260_/S vssd1 vssd1 vccd1 vccd1 _25257_/A sky130_fd_sc_hd__mux2_1
X_13270_ _17658_/A _25583_/Q vssd1 vssd1 vccd1 vccd1 _13976_/A sky130_fd_sc_hd__nand2_4
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22468_ _24415_/A vssd1 vssd1 vccd1 vccd1 _22468_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_185_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24207_ _26959_/Q _24205_/B _24206_/Y vssd1 vssd1 vccd1 vccd1 _26959_/D sky130_fd_sc_hd__o21a_1
X_21419_ _20656_/A _21415_/X _21350_/A _21418_/X vssd1 vssd1 vccd1 vccd1 _21419_/X
+ sky130_fd_sc_hd__o211a_1
X_22399_ _22394_/A _22381_/X _22389_/X _22405_/A vssd1 vssd1 vccd1 vccd1 _22400_/B
+ sky130_fd_sc_hd__o211a_1
X_25187_ _25217_/A vssd1 vssd1 vccd1 vccd1 _25187_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24138_ _26935_/Q _23597_/X _24142_/S vssd1 vssd1 vccd1 vccd1 _24139_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_169_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25737_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_123_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16960_ _16960_/A vssd1 vssd1 vccd1 vccd1 _16960_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24069_ _24069_/A vssd1 vssd1 vccd1 vccd1 _26904_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15911_ _13009_/A _15913_/A _15910_/X _14124_/B vssd1 vssd1 vccd1 vccd1 _15911_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_277_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16891_ _16955_/B _16841_/B _16840_/Y _16868_/A _16939_/B vssd1 vssd1 vccd1 vccd1
+ _16891_/X sky130_fd_sc_hd__o221a_1
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18630_ _18630_/A _18630_/B vssd1 vssd1 vccd1 vccd1 _18631_/A sky130_fd_sc_hd__and2_1
X_15842_ _26502_/Q _26374_/Q _15842_/S vssd1 vssd1 vccd1 vccd1 _15843_/B sky130_fd_sc_hd__mux2_1
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ _27077_/Q _18508_/X _18509_/X _27175_/Q _18510_/X vssd1 vssd1 vccd1 vccd1
+ _18561_/X sky130_fd_sc_hd__a221o_1
XFILLER_246_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _13347_/A _15771_/X _15772_/X _14228_/X vssd1 vssd1 vccd1 vccd1 _15773_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12985_ _14348_/S vssd1 vssd1 vccd1 vccd1 _13993_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ _19455_/B _18077_/A _17662_/A _17971_/A vssd1 vssd1 vccd1 vccd1 _17512_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_261_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _14724_/A vssd1 vssd1 vccd1 vccd1 _14724_/X sky130_fd_sc_hd__buf_2
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18492_ _18492_/A _18492_/B vssd1 vssd1 vccd1 vccd1 _18492_/Y sky130_fd_sc_hd__nor2_1
XFILLER_206_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17443_ _17443_/A _17443_/B vssd1 vssd1 vccd1 vccd1 _19570_/C sky130_fd_sc_hd__nand2_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14655_ _16243_/B vssd1 vssd1 vccd1 vccd1 _15026_/B sky130_fd_sc_hd__buf_2
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13606_ _13433_/X _13598_/X _13605_/X _13112_/A vssd1 vssd1 vccd1 vccd1 _13606_/X
+ sky130_fd_sc_hd__o211a_1
X_17374_ _25543_/Q _17372_/B _17373_/Y vssd1 vssd1 vccd1 vccd1 _25543_/D sky130_fd_sc_hd__o21a_1
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14586_ _15012_/S vssd1 vssd1 vccd1 vccd1 _18059_/A sky130_fd_sc_hd__buf_4
XFILLER_220_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19113_ _19104_/X _19107_/X _19112_/X vssd1 vssd1 vccd1 vccd1 _19113_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16325_ _26645_/Q _26741_/Q _16325_/S vssd1 vssd1 vccd1 vccd1 _16325_/X sky130_fd_sc_hd__mux2_1
X_13537_ _26498_/Q _26370_/Q _15857_/S vssd1 vssd1 vccd1 vccd1 _13537_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19044_ _25616_/Q _18971_/X _19043_/X _19007_/X vssd1 vssd1 vccd1 vccd1 _25616_/D
+ sky130_fd_sc_hd__o211a_1
X_16256_ _26931_/Q _16256_/B vssd1 vssd1 vccd1 vccd1 _16256_/X sky130_fd_sc_hd__or2_1
X_13468_ _25582_/Q vssd1 vssd1 vccd1 vccd1 _14535_/A sky130_fd_sc_hd__clkbuf_2
X_15207_ _16278_/S vssd1 vssd1 vccd1 vccd1 _16442_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_145_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16187_ _14742_/A _25779_/Q _16255_/S _26865_/Q _15301_/S vssd1 vssd1 vccd1 vccd1
+ _16187_/X sky130_fd_sc_hd__o221a_1
X_13399_ _15532_/B vssd1 vssd1 vccd1 vccd1 _16130_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15138_ _25622_/Q _14597_/A _15137_/X _14618_/A vssd1 vssd1 vccd1 vccd1 _23587_/A
+ sky130_fd_sc_hd__o22a_4
X_15069_ _14881_/A _15060_/X _15068_/Y _14706_/X vssd1 vssd1 vccd1 vccd1 _15069_/X
+ sky130_fd_sc_hd__o211a_1
X_19946_ _19946_/A vssd1 vssd1 vccd1 vccd1 _20652_/A sky130_fd_sc_hd__buf_8
XFILLER_87_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19877_ _20079_/A vssd1 vssd1 vccd1 vccd1 _19877_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18828_ _26954_/Q _18826_/X _18827_/X _26986_/Q vssd1 vssd1 vccd1 vccd1 _18828_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_83_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18759_ _18821_/A vssd1 vssd1 vccd1 vccd1 _18759_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21770_ _20580_/X _26018_/Q _21776_/S vssd1 vssd1 vccd1 vccd1 _21771_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20721_ _20721_/A vssd1 vssd1 vccd1 vccd1 _25758_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23440_ _23440_/A vssd1 vssd1 vccd1 vccd1 _26652_/D sky130_fd_sc_hd__clkbuf_1
X_20652_ _20652_/A _20656_/B vssd1 vssd1 vccd1 vccd1 _20652_/X sky130_fd_sc_hd__or2_1
X_23371_ _26622_/Q _23044_/X _23375_/S vssd1 vssd1 vccd1 vccd1 _23372_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20583_ _23581_/A vssd1 vssd1 vccd1 vccd1 _23757_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25110_ _24725_/Y _25097_/X _25108_/Y _25109_/X vssd1 vssd1 vccd1 vccd1 _25110_/X
+ sky130_fd_sc_hd__a31o_1
X_22322_ _26219_/Q _22315_/X _22321_/X _22319_/X vssd1 vssd1 vccd1 vccd1 _26219_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26090_ _27257_/CLK _26090_/D vssd1 vssd1 vccd1 vccd1 _26090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22253_ _26197_/Q _22235_/X _22252_/X _22243_/X vssd1 vssd1 vccd1 vccd1 _26197_/D
+ sky130_fd_sc_hd__o211a_1
X_25041_ _24668_/Y _25014_/X _25040_/Y _25027_/X vssd1 vssd1 vccd1 vccd1 _25041_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_118_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_3_0_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_21204_ _24457_/A vssd1 vssd1 vccd1 vccd1 _24501_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22184_ _26179_/Q _22169_/X _22183_/X _22181_/X vssd1 vssd1 vccd1 vccd1 _26179_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21135_ _25918_/Q _21130_/X _21131_/X input17/X vssd1 vssd1 vccd1 vccd1 _21136_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_105_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26992_ _26992_/CLK _26992_/D vssd1 vssd1 vccd1 vccd1 _26992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25943_ _27058_/CLK _25943_/D vssd1 vssd1 vccd1 vccd1 _25943_/Q sky130_fd_sc_hd__dfxtp_1
X_21066_ _25935_/Q _21065_/Y _25901_/Q vssd1 vssd1 vccd1 vccd1 _21070_/B sky130_fd_sc_hd__o21ba_1
XFILLER_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20017_ _25673_/Q _25672_/Q _20017_/C vssd1 vssd1 vccd1 vccd1 _20030_/B sky130_fd_sc_hd__and3_1
XFILLER_274_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25874_ _27267_/CLK _25874_/D vssd1 vssd1 vccd1 vccd1 _25874_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_246_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24825_ _27112_/Q _24837_/B vssd1 vssd1 vccd1 vccd1 _24825_/Y sky130_fd_sc_hd__nand2_1
XFILLER_246_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12770_ _12770_/A vssd1 vssd1 vccd1 vccd1 _12771_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_215_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24756_ _27095_/Q _24744_/X _25147_/A _24740_/X vssd1 vssd1 vccd1 vccd1 _24757_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_21968_ _26098_/Q _20878_/X _21972_/S vssd1 vssd1 vccd1 vccd1 _21969_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23707_ _23706_/X _26754_/Q _23716_/S vssd1 vssd1 vccd1 vccd1 _23708_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20919_ _23734_/A vssd1 vssd1 vccd1 vccd1 _20919_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24687_ _27079_/Q _24680_/X _24686_/Y _24676_/X vssd1 vssd1 vccd1 vccd1 _24688_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_21899_ _21899_/A vssd1 vssd1 vccd1 vccd1 _26067_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26426_ _27264_/CLK _26426_/D vssd1 vssd1 vccd1 vccd1 _26426_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_230_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14440_ _14432_/X _14439_/X _14440_/S vssd1 vssd1 vccd1 vccd1 _14440_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23638_ _23638_/A vssd1 vssd1 vccd1 vccd1 _26726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14371_ _13644_/X _14369_/X _14370_/X _13358_/A vssd1 vssd1 vccd1 vccd1 _14371_/X
+ sky130_fd_sc_hd__a211o_1
X_26357_ _27292_/CLK _26357_/D vssd1 vssd1 vccd1 vccd1 _26357_/Q sky130_fd_sc_hd__dfxtp_2
X_23569_ _26702_/Q _23568_/X _23572_/S vssd1 vssd1 vccd1 vccd1 _23570_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16110_ _25816_/Q _27250_/Q _16110_/S vssd1 vssd1 vccd1 vccd1 _16111_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13322_ _15394_/A _13316_/X _13321_/X _13291_/X vssd1 vssd1 vccd1 vccd1 _13322_/X
+ sky130_fd_sc_hd__o211a_1
X_25308_ _25308_/A vssd1 vssd1 vccd1 vccd1 _27256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17090_ _26233_/Q _26232_/Q vssd1 vssd1 vccd1 vccd1 _17091_/B sky130_fd_sc_hd__nand2_1
XFILLER_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26288_ _26292_/CLK _26288_/D vssd1 vssd1 vccd1 vccd1 _26288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16041_ _16628_/B _18851_/B _18862_/S vssd1 vssd1 vccd1 vccd1 _16627_/B sky130_fd_sc_hd__o21bai_4
X_13253_ _13472_/A vssd1 vssd1 vccd1 vccd1 _13254_/A sky130_fd_sc_hd__clkbuf_4
X_25239_ _25208_/A _19620_/X _24771_/X _24758_/B _25219_/X vssd1 vssd1 vccd1 vccd1
+ _25239_/X sky130_fd_sc_hd__a221o_1
XFILLER_182_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13184_ _13641_/A _25583_/Q vssd1 vssd1 vccd1 vccd1 _13365_/A sky130_fd_sc_hd__and2_4
XFILLER_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19800_ _19800_/A _20055_/B vssd1 vssd1 vccd1 vccd1 _19800_/X sky130_fd_sc_hd__or2_1
XFILLER_2_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17992_ _17992_/A _17992_/B _17669_/A vssd1 vssd1 vccd1 vccd1 _18214_/A sky130_fd_sc_hd__or3b_4
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19731_ _17669_/B _19589_/B _18027_/A _16476_/S vssd1 vssd1 vccd1 vccd1 _19776_/B
+ sky130_fd_sc_hd__o2bb2a_2
X_16943_ _16986_/A _16943_/B vssd1 vssd1 vccd1 vccd1 _16944_/A sky130_fd_sc_hd__and2_1
XFILLER_278_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19662_ _20034_/B vssd1 vssd1 vccd1 vccd1 _19882_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16874_ _16855_/A _16872_/X _16873_/X _16842_/A vssd1 vssd1 vccd1 vccd1 _16875_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_77_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15825_ _26110_/Q _26011_/Q _15825_/S vssd1 vssd1 vccd1 vccd1 _15825_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18613_ _27110_/Q _18504_/A _18610_/X _18612_/X vssd1 vssd1 vccd1 vccd1 _18613_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_219_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19593_ _19583_/Y _19586_/X _17512_/X vssd1 vssd1 vccd1 vccd1 _19911_/A sky130_fd_sc_hd__a21o_4
XFILLER_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15756_ _13351_/A _26891_/Q _26763_/Q _15197_/A _13359_/A vssd1 vssd1 vccd1 vccd1
+ _15756_/X sky130_fd_sc_hd__a221o_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18544_ _18544_/A _18544_/B vssd1 vssd1 vccd1 vccd1 _18544_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12968_ _25498_/Q vssd1 vssd1 vccd1 vccd1 _21630_/A sky130_fd_sc_hd__clkinv_4
Xclkbuf_leaf_66_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27269_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14707_ _14956_/A _14700_/X _14704_/Y _14706_/X vssd1 vssd1 vccd1 vccd1 _14707_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_221_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18475_ _18382_/X _18474_/Y _17671_/X vssd1 vssd1 vccd1 vccd1 _18475_/X sky130_fd_sc_hd__o21a_1
XFILLER_206_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15687_ _27311_/Q _26568_/Q _16178_/S vssd1 vssd1 vccd1 vccd1 _15687_/X sky130_fd_sc_hd__mux2_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _12899_/A vssd1 vssd1 vccd1 vccd1 _13737_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_21_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _17427_/A _17427_/C _25560_/Q vssd1 vssd1 vccd1 vccd1 _17428_/B sky130_fd_sc_hd__a21oi_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14638_ _27325_/Q _26582_/Q _14652_/S vssd1 vssd1 vccd1 vccd1 _14638_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17357_ _17356_/X _17360_/C _17318_/X vssd1 vssd1 vccd1 vccd1 _17357_/Y sky130_fd_sc_hd__a21oi_1
X_14569_ _16706_/A _16706_/B _16707_/B vssd1 vssd1 vccd1 vccd1 _16713_/B sky130_fd_sc_hd__a21oi_1
XFILLER_174_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16308_ _16306_/X _16307_/X _16308_/S vssd1 vssd1 vccd1 vccd1 _16308_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17288_ _17287_/X _17293_/C _17269_/X vssd1 vssd1 vccd1 vccd1 _17288_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19027_ _26959_/Q _18826_/X _18827_/X _26991_/Q vssd1 vssd1 vccd1 vccd1 _19027_/X
+ sky130_fd_sc_hd__a22o_1
X_16239_ _26351_/Q _26611_/Q _16240_/S vssd1 vssd1 vccd1 vccd1 _16239_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19929_ _19930_/A _27077_/Q vssd1 vssd1 vccd1 vccd1 _19933_/A sky130_fd_sc_hd__or2_1
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22940_ _22940_/A vssd1 vssd1 vccd1 vccd1 _26445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22871_ _26415_/Q _22717_/X _22873_/S vssd1 vssd1 vccd1 vccd1 _22872_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24610_ _24610_/A vssd1 vssd1 vccd1 vccd1 _24621_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21822_ _21822_/A vssd1 vssd1 vccd1 vccd1 _26040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25590_ _25590_/CLK _25590_/D vssd1 vssd1 vccd1 vccd1 _25590_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_37_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24541_ _24989_/A _24541_/B vssd1 vssd1 vccd1 vccd1 _25206_/D sky130_fd_sc_hd__nand2_2
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21753_ _21753_/A vssd1 vssd1 vccd1 vccd1 _26010_/D sky130_fd_sc_hd__clkbuf_1
XPHY_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20704_ _26292_/Q _20687_/B _20703_/Y _20697_/X vssd1 vssd1 vccd1 vccd1 _25755_/D
+ sky130_fd_sc_hd__o211a_1
X_27260_ _27324_/CLK _27260_/D vssd1 vssd1 vccd1 vccd1 _27260_/Q sky130_fd_sc_hd__dfxtp_1
X_24472_ _24472_/A vssd1 vssd1 vccd1 vccd1 _24472_/X sky130_fd_sc_hd__buf_2
X_21684_ _21684_/A vssd1 vssd1 vccd1 vccd1 _25981_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26211_ _26974_/CLK _26211_/D vssd1 vssd1 vccd1 vccd1 _26211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23423_ _23423_/A vssd1 vssd1 vccd1 vccd1 _26645_/D sky130_fd_sc_hd__clkbuf_1
X_20635_ _20635_/A _20643_/B vssd1 vssd1 vccd1 vccd1 _20635_/X sky130_fd_sc_hd__or2_1
X_27191_ _27196_/CLK _27191_/D vssd1 vssd1 vccd1 vccd1 _27191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26142_ _26599_/CLK _26142_/D vssd1 vssd1 vccd1 vccd1 _26142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20566_ _23568_/A vssd1 vssd1 vccd1 vccd1 _23744_/A sky130_fd_sc_hd__clkbuf_2
X_23354_ _23354_/A vssd1 vssd1 vccd1 vccd1 _26615_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22305_ _26213_/Q _22299_/X _22302_/X _22304_/X vssd1 vssd1 vccd1 vccd1 _26213_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26073_ _26595_/CLK _26073_/D vssd1 vssd1 vccd1 vccd1 _26073_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_164_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20497_ _20496_/X _25693_/Q _20509_/S vssd1 vssd1 vccd1 vccd1 _20498_/A sky130_fd_sc_hd__mux2_1
X_23285_ _26585_/Q input248/X _23289_/S vssd1 vssd1 vccd1 vccd1 _23286_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25024_ _25024_/A vssd1 vssd1 vccd1 vccd1 _25024_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22236_ _26230_/Q _22416_/B _22236_/C vssd1 vssd1 vccd1 vccd1 _22630_/B sky130_fd_sc_hd__and3_2
X_22167_ _26173_/Q _22154_/X _22115_/X _22166_/X _22155_/X vssd1 vssd1 vccd1 vccd1
+ _22167_/X sky130_fd_sc_hd__a221o_1
XFILLER_106_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21118_ _21118_/A _21118_/B vssd1 vssd1 vccd1 vccd1 _21119_/A sky130_fd_sc_hd__or2_1
XFILLER_8_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26975_ _26980_/CLK _26975_/D vssd1 vssd1 vccd1 vccd1 _26975_/Q sky130_fd_sc_hd__dfxtp_1
X_22098_ _22098_/A vssd1 vssd1 vccd1 vccd1 _26156_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13940_ _13512_/A _13936_/X _13938_/X _13939_/X vssd1 vssd1 vccd1 vccd1 _13947_/B
+ sky130_fd_sc_hd__o211a_1
X_21049_ _21049_/A vssd1 vssd1 vccd1 vccd1 _25893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25926_ _27213_/CLK _25926_/D vssd1 vssd1 vccd1 vccd1 _25926_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13871_ _14109_/B vssd1 vssd1 vccd1 vccd1 _14273_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25857_ _26453_/CLK _25857_/D vssd1 vssd1 vccd1 vccd1 _25857_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_207_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15610_ _15610_/A _15610_/B vssd1 vssd1 vccd1 vccd1 _15610_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12822_ _12822_/A vssd1 vssd1 vccd1 vccd1 _12953_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_24808_ _24806_/Y _24807_/X _24796_/X vssd1 vssd1 vccd1 vccd1 _27107_/D sky130_fd_sc_hd__a21oi_1
X_16590_ _16962_/A _19571_/B vssd1 vssd1 vccd1 vccd1 _16957_/A sky130_fd_sc_hd__nand2_1
XFILLER_90_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25788_ _27293_/CLK _25788_/D vssd1 vssd1 vccd1 vccd1 _25788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15541_ _27248_/Q _15635_/B vssd1 vssd1 vccd1 vccd1 _15541_/X sky130_fd_sc_hd__or2_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ _13945_/A vssd1 vssd1 vccd1 vccd1 _12754_/A sky130_fd_sc_hd__clkbuf_4
X_24739_ _24739_/A _24739_/B vssd1 vssd1 vccd1 vccd1 _24739_/Y sky130_fd_sc_hd__nand2_4
XFILLER_203_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _18256_/X _18259_/X _18487_/A vssd1 vssd1 vccd1 vccd1 _18260_/X sky130_fd_sc_hd__mux2_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15472_ _26506_/Q _26378_/Q _15796_/S vssd1 vssd1 vccd1 vccd1 _15472_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12684_ _13641_/A _25566_/Q _25565_/Q vssd1 vssd1 vccd1 vccd1 _18028_/B sky130_fd_sc_hd__and3_2
XFILLER_187_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _19847_/A vssd1 vssd1 vccd1 vccd1 _17443_/B sky130_fd_sc_hd__buf_6
XFILLER_230_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14423_ _27232_/Q _15725_/S _13124_/A _14422_/X vssd1 vssd1 vccd1 vccd1 _14423_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_187_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26409_ _27280_/CLK _26409_/D vssd1 vssd1 vccd1 vccd1 _26409_/Q sky130_fd_sc_hd__dfxtp_1
X_18191_ _18364_/A vssd1 vssd1 vccd1 vccd1 _18191_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17142_ _17200_/A _17142_/B vssd1 vssd1 vccd1 vccd1 _17143_/A sky130_fd_sc_hd__and2_1
X_14354_ _14346_/X _14353_/X _14354_/S vssd1 vssd1 vccd1 vccd1 _14355_/B sky130_fd_sc_hd__mux2_1
XFILLER_168_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_184_wb_clk_i _26681_/CLK vssd1 vssd1 vccd1 vccd1 _26905_/CLK sky130_fd_sc_hd__clkbuf_16
X_13305_ _13305_/A vssd1 vssd1 vccd1 vccd1 _13467_/A sky130_fd_sc_hd__buf_4
XFILLER_6_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17073_ _22350_/S vssd1 vssd1 vccd1 vccd1 _22340_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_156_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14285_ _14566_/A _14566_/B vssd1 vssd1 vccd1 vccd1 _18317_/S sky130_fd_sc_hd__nor2_4
XFILLER_109_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_113_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26987_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16024_ _13835_/A _26920_/Q _26404_/Q _15515_/S _13827_/A vssd1 vssd1 vccd1 vccd1
+ _16024_/X sky130_fd_sc_hd__a221o_1
XFILLER_6_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13236_ _15424_/A _13236_/B vssd1 vssd1 vccd1 vccd1 _13236_/X sky130_fd_sc_hd__or2_1
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13167_ _14523_/A vssd1 vssd1 vccd1 vccd1 _13168_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_152_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13098_ _14352_/S vssd1 vssd1 vccd1 vccd1 _14107_/A sky130_fd_sc_hd__clkbuf_2
X_17975_ _17975_/A vssd1 vssd1 vccd1 vccd1 _18254_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19714_ _19766_/A _19712_/Y _19926_/A vssd1 vssd1 vccd1 vccd1 _19714_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_238_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16926_ _16951_/A vssd1 vssd1 vccd1 vccd1 _16986_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_272_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19645_ _27069_/Q _19870_/B _27135_/Q vssd1 vssd1 vccd1 vccd1 _19645_/X sky130_fd_sc_hd__a21o_1
XFILLER_253_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16857_ _16864_/A _16857_/B vssd1 vssd1 vccd1 vccd1 _16858_/A sky130_fd_sc_hd__and2_1
XFILLER_92_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15808_ _25883_/Q _15808_/B vssd1 vssd1 vccd1 vccd1 _15808_/X sky130_fd_sc_hd__or2_1
X_16788_ _16788_/A vssd1 vssd1 vccd1 vccd1 _16794_/B sky130_fd_sc_hd__clkbuf_4
X_19576_ _19574_/X _19576_/B _19576_/C _19576_/D vssd1 vssd1 vccd1 vccd1 _19576_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_92_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15739_ _26503_/Q _26375_/Q _15989_/S vssd1 vssd1 vccd1 vccd1 _15739_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18527_ _18435_/X _18524_/X _18526_/X vssd1 vssd1 vccd1 vccd1 _18527_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18458_ _18458_/A vssd1 vssd1 vccd1 vccd1 _18459_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17409_ _17428_/A _17409_/B _17410_/B vssd1 vssd1 vccd1 vccd1 _25554_/D sky130_fd_sc_hd__nor3_1
X_18389_ _18812_/A vssd1 vssd1 vccd1 vccd1 _18504_/A sky130_fd_sc_hd__clkbuf_2
X_20420_ _22531_/A _20420_/B _20420_/C vssd1 vssd1 vccd1 vccd1 _20467_/C sky130_fd_sc_hd__and3_2
XFILLER_267_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20351_ _20351_/A _20351_/B vssd1 vssd1 vccd1 vccd1 _20352_/B sky130_fd_sc_hd__nand2_1
XFILLER_146_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23070_ _23137_/S vssd1 vssd1 vccd1 vccd1 _23083_/S sky130_fd_sc_hd__buf_6
X_20282_ _25747_/Q _19727_/X _20281_/X _19920_/A vssd1 vssd1 vccd1 vccd1 _20283_/B
+ sky130_fd_sc_hd__o22a_1
X_22021_ _26122_/Q _20955_/X _22027_/S vssd1 vssd1 vccd1 vccd1 _22022_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26760_ _27307_/CLK _26760_/D vssd1 vssd1 vccd1 vccd1 _26760_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23972_ _26861_/Q _23565_/X _23976_/S vssd1 vssd1 vccd1 vccd1 _23973_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25711_ _26673_/CLK _25711_/D vssd1 vssd1 vccd1 vccd1 _25711_/Q sky130_fd_sc_hd__dfxtp_1
X_22923_ _26438_/Q _22688_/X _22923_/S vssd1 vssd1 vccd1 vccd1 _22924_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26691_ _26916_/CLK _26691_/D vssd1 vssd1 vccd1 vccd1 _26691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25642_ _25661_/CLK _25642_/D vssd1 vssd1 vccd1 vccd1 _25642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22854_ _26407_/Q _22691_/X _22862_/S vssd1 vssd1 vccd1 vccd1 _22855_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21805_ _26033_/Q _20884_/X _21805_/S vssd1 vssd1 vccd1 vccd1 _21806_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25573_ _25590_/CLK _25573_/D vssd1 vssd1 vccd1 vccd1 _25573_/Q sky130_fd_sc_hd__dfxtp_4
X_22785_ _26377_/Q _22698_/X _22789_/S vssd1 vssd1 vccd1 vccd1 _22786_/A sky130_fd_sc_hd__mux2_1
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27312_ _27312_/CLK _27312_/D vssd1 vssd1 vccd1 vccd1 _27312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24524_ _27033_/Q _24506_/X _24522_/Y _24523_/X vssd1 vssd1 vccd1 vccd1 _27033_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21736_ _21736_/A vssd1 vssd1 vccd1 vccd1 _26002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27243_ _27307_/CLK _27243_/D vssd1 vssd1 vccd1 vccd1 _27243_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24455_ _24455_/A vssd1 vssd1 vccd1 vccd1 _24455_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21667_ _21667_/A vssd1 vssd1 vccd1 vccd1 _25973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23406_ _26638_/Q _23095_/X _23408_/S vssd1 vssd1 vccd1 vccd1 _23407_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27174_ _27198_/CLK _27174_/D vssd1 vssd1 vccd1 vccd1 _27174_/Q sky130_fd_sc_hd__dfxtp_1
X_20618_ _20617_/X _25722_/Q _20622_/S vssd1 vssd1 vccd1 vccd1 _20619_/A sky130_fd_sc_hd__mux2_1
X_24386_ _24381_/X _25602_/Q _24385_/X vssd1 vssd1 vccd1 vccd1 _24659_/B sky130_fd_sc_hd__o21a_4
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21598_ _25962_/Q _21573_/X _21596_/Y _21597_/X vssd1 vssd1 vccd1 vccd1 _25962_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_193_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26125_ _27292_/CLK _26125_/D vssd1 vssd1 vccd1 vccd1 _26125_/Q sky130_fd_sc_hd__dfxtp_1
X_23337_ _23348_/A vssd1 vssd1 vccd1 vccd1 _23346_/S sky130_fd_sc_hd__clkbuf_4
X_20549_ _23555_/A vssd1 vssd1 vccd1 vccd1 _23731_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_137_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14070_ _26657_/Q _25697_/Q _14474_/S vssd1 vssd1 vccd1 vccd1 _14070_/X sky130_fd_sc_hd__mux2_1
X_26056_ _26900_/CLK _26056_/D vssd1 vssd1 vccd1 vccd1 _26056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23268_ _23268_/A vssd1 vssd1 vccd1 vccd1 _23277_/S sky130_fd_sc_hd__buf_4
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13021_ _13139_/A vssd1 vssd1 vccd1 vccd1 _13022_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_152_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25007_ _20624_/A _25003_/X _25006_/X vssd1 vssd1 vccd1 vccd1 _25007_/Y sky130_fd_sc_hd__o21ai_1
X_22219_ input6/X input281/X _22226_/S vssd1 vssd1 vccd1 vccd1 _22219_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23199_ _26546_/Q _23121_/X _23205_/S vssd1 vssd1 vccd1 vccd1 _23200_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17760_ _17752_/X _17755_/X _18756_/A _27005_/Q _18821_/A vssd1 vssd1 vccd1 vccd1
+ _17760_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14972_ _26092_/Q _14960_/B _14969_/S _14971_/X vssd1 vssd1 vccd1 vccd1 _14972_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26958_ _26992_/CLK _26958_/D vssd1 vssd1 vccd1 vccd1 _26958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_266_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13923_ _14025_/A _13923_/B _14025_/B vssd1 vssd1 vccd1 vccd1 _13923_/X sky130_fd_sc_hd__or3_1
X_16711_ _16711_/A _17800_/C vssd1 vssd1 vccd1 vccd1 _18324_/A sky130_fd_sc_hd__and2_1
X_17691_ _17691_/A _17691_/B vssd1 vssd1 vccd1 vccd1 _17691_/X sky130_fd_sc_hd__or2_2
X_25909_ _27122_/CLK _25909_/D vssd1 vssd1 vccd1 vccd1 _25909_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_267_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26889_ _26889_/CLK _26889_/D vssd1 vssd1 vccd1 vccd1 _26889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19430_ _19423_/X _19426_/Y _19429_/X _18738_/X vssd1 vssd1 vccd1 vccd1 _19430_/X
+ sky130_fd_sc_hd__a22o_1
X_16642_ _25796_/Q _21070_/A vssd1 vssd1 vccd1 vccd1 _16642_/Y sky130_fd_sc_hd__nor2_1
XFILLER_262_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13854_ _27302_/Q _26559_/Q _15807_/S vssd1 vssd1 vccd1 vccd1 _13854_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_405 _17043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_416 _17009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12805_ _13215_/A _25578_/Q _25577_/Q vssd1 vssd1 vccd1 vccd1 _14358_/B sky130_fd_sc_hd__and3_1
XFILLER_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16573_ _16573_/A _16573_/B vssd1 vssd1 vccd1 vccd1 _16773_/A sky130_fd_sc_hd__nor2_1
XINSDIODE2_427 _12781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19361_ _18682_/X _18269_/B _19360_/X _19018_/A vssd1 vssd1 vccd1 vccd1 _19361_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_250_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13785_ _13266_/A _26692_/Q _26820_/Q _13262_/A _14768_/A vssd1 vssd1 vccd1 vccd1
+ _13785_/X sky130_fd_sc_hd__a221o_1
XFILLER_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_438 _25729_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_449 _26940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15524_ _13207_/A _23568_/A _15523_/Y _13214_/A vssd1 vssd1 vccd1 vccd1 _19031_/A
+ sky130_fd_sc_hd__o211ai_4
X_18312_ _18040_/X _18311_/X _17988_/A vssd1 vssd1 vccd1 vccd1 _18312_/Y sky130_fd_sc_hd__o21ai_1
X_12736_ _12736_/A vssd1 vssd1 vccd1 vccd1 _13664_/A sky130_fd_sc_hd__buf_2
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19292_ _19325_/A _19292_/B vssd1 vssd1 vccd1 vccd1 _19577_/B sky130_fd_sc_hd__xnor2_2
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18243_ _26944_/Q _18826_/A _18827_/A _26976_/Q vssd1 vssd1 vccd1 vccd1 _18243_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15455_ _26670_/Q _16069_/S _15454_/X _13051_/A vssd1 vssd1 vccd1 vccd1 _15455_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_188_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14406_ _14237_/B _13574_/X _14405_/X _14610_/A vssd1 vssd1 vccd1 vccd1 _14406_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18174_ _17347_/X _18825_/A _18171_/X _18829_/A _18830_/A vssd1 vssd1 vccd1 vccd1
+ _18174_/X sky130_fd_sc_hd__a221o_1
X_15386_ _15187_/X _15377_/X _15385_/X _14709_/A vssd1 vssd1 vccd1 vccd1 _15386_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_156_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17125_ _25471_/Q _17105_/X _17107_/X _25568_/Q vssd1 vssd1 vccd1 vccd1 _17126_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14337_ _26066_/Q _25871_/Q _14513_/S vssd1 vssd1 vccd1 vccd1 _14337_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17056_ _20798_/B _17056_/B vssd1 vssd1 vccd1 vccd1 _20794_/C sky130_fd_sc_hd__nand2_2
X_14268_ _14264_/X _14267_/X _14268_/S vssd1 vssd1 vccd1 vccd1 _14268_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16007_ _15516_/A _16004_/X _16006_/X _13832_/A vssd1 vssd1 vccd1 vccd1 _16007_/X
+ sky130_fd_sc_hd__o211a_1
X_13219_ _15916_/A vssd1 vssd1 vccd1 vccd1 _13284_/A sky130_fd_sc_hd__buf_2
X_14199_ _15588_/A _25833_/Q _26033_/Q _13675_/S _13644_/X vssd1 vssd1 vccd1 vccd1
+ _14199_/X sky130_fd_sc_hd__a221o_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_10_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_10_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _17956_/X _17957_/X _17958_/S vssd1 vssd1 vccd1 vccd1 _17958_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_81_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27299_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_238_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16909_ _16938_/B vssd1 vssd1 vccd1 vccd1 _16909_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17889_ _17881_/X _17886_/Y _18044_/S vssd1 vssd1 vccd1 vccd1 _17889_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_opt_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26609_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19628_ _19628_/A _19628_/B _19628_/C vssd1 vssd1 vccd1 vccd1 _25173_/A sky130_fd_sc_hd__nor3_4
XFILLER_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19559_ _25657_/Q _19563_/B vssd1 vssd1 vccd1 vccd1 _19559_/X sky130_fd_sc_hd__or2_1
XFILLER_15_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22570_ _22567_/X _22569_/Y _22561_/X vssd1 vssd1 vccd1 vccd1 _26303_/D sky130_fd_sc_hd__a21oi_1
XFILLER_210_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21521_ _25956_/Q _21506_/X _21520_/Y _21467_/X vssd1 vssd1 vccd1 vccd1 _25956_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_278_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24240_ _26970_/Q _26969_/Q _24240_/C vssd1 vssd1 vccd1 vccd1 _24243_/B sky130_fd_sc_hd__and3_1
X_21452_ _21421_/X _25863_/Q _21450_/Y _21451_/X vssd1 vssd1 vccd1 vccd1 _21452_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20403_ _19381_/A _20355_/X _20402_/Y _20357_/X vssd1 vssd1 vccd1 vccd1 _20405_/B
+ sky130_fd_sc_hd__o22a_1
X_24171_ _24239_/A vssd1 vssd1 vccd1 vccd1 _24188_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21383_ _21342_/X _21382_/X _21336_/X vssd1 vssd1 vccd1 vccd1 _21383_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_162_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23122_ _26514_/Q _23121_/X _23131_/S vssd1 vssd1 vccd1 vccd1 _23123_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20334_ _25685_/Q _25684_/Q _20334_/C vssd1 vssd1 vccd1 vccd1 _20382_/C sky130_fd_sc_hd__and3_1
XFILLER_116_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23053_ _23526_/A vssd1 vssd1 vccd1 vccd1 _23053_/X sky130_fd_sc_hd__buf_2
X_20265_ _20452_/A _20265_/B _20265_/C vssd1 vssd1 vccd1 vccd1 _20265_/X sky130_fd_sc_hd__and3_1
XFILLER_162_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22004_ _22004_/A vssd1 vssd1 vccd1 vccd1 _26114_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20196_ _20677_/A _20091_/A _20195_/Y _20115_/A vssd1 vssd1 vccd1 vccd1 _20299_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput105 dout0[8] vssd1 vssd1 vccd1 vccd1 input105/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput116 dout1[18] vssd1 vssd1 vccd1 vccd1 input116/X sky130_fd_sc_hd__clkbuf_1
XTAP_5338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput127 dout1[28] vssd1 vssd1 vccd1 vccd1 input127/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26812_ _26813_/CLK _26812_/D vssd1 vssd1 vccd1 vccd1 _26812_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput138 dout1[38] vssd1 vssd1 vccd1 vccd1 input138/X sky130_fd_sc_hd__clkbuf_2
XFILLER_248_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput149 dout1[48] vssd1 vssd1 vccd1 vccd1 input149/X sky130_fd_sc_hd__clkbuf_2
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26743_ _26903_/CLK _26743_/D vssd1 vssd1 vccd1 vccd1 _26743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23955_ _23955_/A vssd1 vssd1 vccd1 vccd1 _26853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22906_ _26430_/Q _22663_/X _22912_/S vssd1 vssd1 vccd1 vccd1 _22907_/A sky130_fd_sc_hd__mux2_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26674_ _27317_/CLK _26674_/D vssd1 vssd1 vccd1 vccd1 _26674_/Q sky130_fd_sc_hd__dfxtp_1
X_23886_ _23886_/A vssd1 vssd1 vccd1 vccd1 _26822_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25625_ _27327_/CLK _25625_/D vssd1 vssd1 vccd1 vccd1 _25625_/Q sky130_fd_sc_hd__dfxtp_2
X_22837_ _22837_/A vssd1 vssd1 vccd1 vccd1 _26399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25556_ _25992_/CLK _25556_/D vssd1 vssd1 vccd1 vccd1 _25556_/Q sky130_fd_sc_hd__dfxtp_1
X_13570_ _13570_/A vssd1 vssd1 vccd1 vccd1 _15874_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22768_ _22768_/A vssd1 vssd1 vccd1 vccd1 _26369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24507_ _26318_/Q _24455_/X _24456_/X input232/X _24501_/X vssd1 vssd1 vccd1 vccd1
+ _24507_/X sky130_fd_sc_hd__a221o_1
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21719_ _21719_/A vssd1 vssd1 vccd1 vccd1 _25996_/D sky130_fd_sc_hd__clkbuf_1
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25487_ _26843_/CLK _25487_/D vssd1 vssd1 vccd1 vccd1 _25487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22699_ _26345_/Q _22698_/X _22705_/S vssd1 vssd1 vccd1 vccd1 _22700_/A sky130_fd_sc_hd__mux2_1
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27226_ _27227_/CLK _27226_/D vssd1 vssd1 vccd1 vccd1 _27226_/Q sky130_fd_sc_hd__dfxtp_1
X_15240_ _19240_/S _15240_/B vssd1 vssd1 vccd1 vccd1 _17846_/B sky130_fd_sc_hd__nor2_1
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24438_ _24381_/X _25611_/Q _24437_/X vssd1 vssd1 vccd1 vccd1 _24696_/B sky130_fd_sc_hd__o21a_4
XFILLER_157_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27157_ _27160_/CLK _27157_/D vssd1 vssd1 vccd1 vccd1 _27157_/Q sky130_fd_sc_hd__dfxtp_4
X_15171_ _15165_/X _15166_/X _15170_/X vssd1 vssd1 vccd1 vccd1 _15171_/X sky130_fd_sc_hd__o21a_1
X_24369_ _27006_/Q _24357_/X _24368_/Y _22468_/X vssd1 vssd1 vccd1 vccd1 _27006_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26108_ _27275_/CLK _26108_/D vssd1 vssd1 vccd1 vccd1 _26108_/Q sky130_fd_sc_hd__dfxtp_1
X_14122_ _14101_/X _14121_/X _13172_/A vssd1 vssd1 vccd1 vccd1 _14122_/X sky130_fd_sc_hd__a21o_1
XFILLER_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27088_ _27213_/CLK _27088_/D vssd1 vssd1 vccd1 vccd1 _27088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26039_ _26601_/CLK _26039_/D vssd1 vssd1 vccd1 vccd1 _26039_/Q sky130_fd_sc_hd__dfxtp_2
X_14053_ _14051_/X _14052_/X _14473_/S vssd1 vssd1 vccd1 vccd1 _14053_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18930_ _18891_/X _18894_/X _18928_/X _18929_/X vssd1 vssd1 vccd1 vccd1 _18931_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13004_ _20485_/A _14354_/S _13015_/A _23363_/B _13003_/Y vssd1 vssd1 vccd1 vccd1
+ _13005_/C sky130_fd_sc_hd__a221o_1
XFILLER_234_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18861_ _18861_/A vssd1 vssd1 vccd1 vccd1 _18861_/X sky130_fd_sc_hd__buf_2
XFILLER_267_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17812_ _18251_/B _18251_/C _18251_/A vssd1 vssd1 vccd1 vccd1 _18325_/B sky130_fd_sc_hd__a21oi_2
XFILLER_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18792_ _18792_/A vssd1 vssd1 vccd1 vccd1 _18792_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17743_ _18615_/A vssd1 vssd1 vccd1 vccd1 _18952_/B sky130_fd_sc_hd__clkbuf_2
X_14955_ _12751_/A _14953_/X _14954_/X vssd1 vssd1 vccd1 vccd1 _14956_/B sky130_fd_sc_hd__o21ai_1
XFILLER_208_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13906_ _13636_/B _16833_/B _13904_/X _15948_/B vssd1 vssd1 vccd1 vccd1 _13908_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_263_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17674_ _26063_/Q vssd1 vssd1 vccd1 vccd1 _17708_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14886_ _16250_/A _14886_/B vssd1 vssd1 vccd1 vccd1 _14886_/X sky130_fd_sc_hd__or2_1
XFILLER_263_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19413_ _25753_/Q _19414_/B vssd1 vssd1 vccd1 vccd1 _19421_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_202 _14480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13837_ _13835_/X _26851_/Q _25765_/Q _15514_/S _13775_/A vssd1 vssd1 vccd1 vccd1
+ _13837_/X sky130_fd_sc_hd__a221o_1
X_16625_ _16625_/A vssd1 vssd1 vccd1 vccd1 _18941_/A sky130_fd_sc_hd__inv_2
XINSDIODE2_213 _16901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_224 _23549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_235 _19046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_246 _16735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_257 _24630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16556_ _16556_/A _19393_/A vssd1 vssd1 vccd1 vccd1 _16557_/A sky130_fd_sc_hd__nor2_1
X_19344_ _19196_/X _19342_/Y _19343_/X _16566_/A _19076_/X vssd1 vssd1 vccd1 vccd1
+ _19344_/X sky130_fd_sc_hd__o32a_2
X_13768_ _13766_/X _13767_/X _13779_/A vssd1 vssd1 vccd1 vccd1 _13768_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_268 _24277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_279 _27327_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15507_ _26798_/Q _26442_/Q _16113_/A vssd1 vssd1 vccd1 vccd1 _15507_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12719_ _25579_/Q vssd1 vssd1 vccd1 vccd1 _18076_/A sky130_fd_sc_hd__buf_2
XFILLER_30_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19275_ _18544_/A _18421_/B _18427_/X _18495_/A vssd1 vssd1 vccd1 vccd1 _19275_/X
+ sky130_fd_sc_hd__o22a_1
X_16487_ _16481_/A _16486_/Y _12706_/A vssd1 vssd1 vccd1 vccd1 _16487_/Y sky130_fd_sc_hd__a21oi_1
X_13699_ _15547_/A vssd1 vssd1 vccd1 vccd1 _15141_/A sky130_fd_sc_hd__buf_2
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15438_ _17790_/A _15438_/B vssd1 vssd1 vccd1 vccd1 _15439_/B sky130_fd_sc_hd__nor2_1
X_18226_ _18226_/A vssd1 vssd1 vccd1 vccd1 _25600_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18157_ _25503_/Q _18807_/A _18808_/A _17347_/X vssd1 vssd1 vccd1 vccd1 _18157_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15369_ _15019_/A _15364_/X _15368_/X _14678_/A vssd1 vssd1 vccd1 vccd1 _15369_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17108_ _25468_/Q _17105_/X _17107_/X _25565_/Q vssd1 vssd1 vccd1 vccd1 _17109_/B
+ sky130_fd_sc_hd__a22o_1
X_18088_ _18088_/A vssd1 vssd1 vccd1 vccd1 _20034_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17039_ _17039_/A vssd1 vssd1 vccd1 vccd1 _17039_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20050_ _27147_/Q _20219_/B vssd1 vssd1 vccd1 vccd1 _20050_/Y sky130_fd_sc_hd__nand2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23740_ _23740_/A vssd1 vssd1 vccd1 vccd1 _26764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_254_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20952_ _20952_/A vssd1 vssd1 vccd1 vccd1 _20965_/S sky130_fd_sc_hd__buf_6
XFILLER_260_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23671_ _23671_/A vssd1 vssd1 vccd1 vccd1 _26741_/D sky130_fd_sc_hd__clkbuf_1
X_20883_ _20883_/A vssd1 vssd1 vccd1 vccd1 _25832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25410_ _25410_/A vssd1 vssd1 vccd1 vccd1 _27301_/D sky130_fd_sc_hd__clkbuf_1
X_22622_ _26324_/Q _22632_/B vssd1 vssd1 vccd1 vccd1 _22622_/Y sky130_fd_sc_hd__nand2_1
X_26390_ _27293_/CLK _26390_/D vssd1 vssd1 vccd1 vccd1 _26390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25341_ _27271_/Q _23712_/A _25343_/S vssd1 vssd1 vccd1 vccd1 _25342_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22553_ _22567_/A vssd1 vssd1 vccd1 vccd1 _22553_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21504_ _21499_/Y _21503_/X _21492_/X vssd1 vssd1 vccd1 vccd1 _21504_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_194_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25272_ _25272_/A vssd1 vssd1 vccd1 vccd1 _27240_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22484_ _22484_/A vssd1 vssd1 vccd1 vccd1 _26267_/D sky130_fd_sc_hd__clkbuf_1
X_27011_ _27044_/CLK _27011_/D vssd1 vssd1 vccd1 vccd1 _27011_/Q sky130_fd_sc_hd__dfxtp_1
X_24223_ _24239_/A vssd1 vssd1 vccd1 vccd1 _24237_/A sky130_fd_sc_hd__clkbuf_2
X_21435_ _20662_/A _21415_/X _21350_/A _21434_/X vssd1 vssd1 vccd1 vccd1 _21435_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24154_ _26942_/Q _24157_/C vssd1 vssd1 vccd1 vccd1 _24160_/C sky130_fd_sc_hd__and2_1
XFILLER_163_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21366_ _21364_/X _18622_/X _21365_/X _25806_/Q _21322_/X vssd1 vssd1 vccd1 vccd1
+ _21366_/X sky130_fd_sc_hd__a221o_1
XFILLER_162_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23105_ _23578_/A vssd1 vssd1 vccd1 vccd1 _23105_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_218_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20317_ _24986_/B _20317_/B _20317_/C vssd1 vssd1 vccd1 vccd1 _20317_/X sky130_fd_sc_hd__or3_1
XFILLER_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24085_ _26911_/Q _23520_/X _24087_/S vssd1 vssd1 vccd1 vccd1 _24086_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21297_ _21556_/A vssd1 vssd1 vccd1 vccd1 _21297_/X sky130_fd_sc_hd__buf_4
XFILLER_27_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23036_ _25393_/A _23291_/B vssd1 vssd1 vccd1 vccd1 _23118_/A sky130_fd_sc_hd__nor2_8
XFILLER_122_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20248_ _20248_/A vssd1 vssd1 vccd1 vccd1 _20248_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20179_ _24810_/A vssd1 vssd1 vccd1 vccd1 _20179_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_276_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24987_ _27165_/Q vssd1 vssd1 vccd1 vccd1 _25208_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_218_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ _26810_/Q _26454_/Q _16510_/A vssd1 vssd1 vccd1 vccd1 _14740_/X sky130_fd_sc_hd__mux2_1
X_23938_ _23938_/A vssd1 vssd1 vccd1 vccd1 _26845_/D sky130_fd_sc_hd__clkbuf_1
X_26726_ _27278_/CLK _26726_/D vssd1 vssd1 vccd1 vccd1 _26726_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26657_ _26657_/CLK _26657_/D vssd1 vssd1 vccd1 vccd1 _26657_/Q sky130_fd_sc_hd__dfxtp_1
X_14671_ _26518_/Q _26390_/Q _14699_/S vssd1 vssd1 vccd1 vccd1 _14671_/X sky130_fd_sc_hd__mux2_1
X_23869_ _23696_/X _26815_/Q _23871_/S vssd1 vssd1 vccd1 vccd1 _23870_/A sky130_fd_sc_hd__mux2_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16410_ _25657_/Q _14609_/A _14613_/X vssd1 vssd1 vccd1 vccd1 _16410_/X sky130_fd_sc_hd__a21o_1
XFILLER_83_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13622_ _26789_/Q _26433_/Q _15725_/S vssd1 vssd1 vccd1 vccd1 _13623_/B sky130_fd_sc_hd__mux2_1
X_25608_ _25725_/CLK _25608_/D vssd1 vssd1 vccd1 vccd1 _25608_/Q sky130_fd_sc_hd__dfxtp_4
X_17390_ _17428_/A _17390_/B _17392_/B vssd1 vssd1 vccd1 vccd1 _25548_/D sky130_fd_sc_hd__nor3_1
XFILLER_220_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26588_ _26909_/CLK _26588_/D vssd1 vssd1 vccd1 vccd1 _26588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16341_ _26121_/Q _26022_/Q _16341_/S vssd1 vssd1 vccd1 vccd1 _16341_/X sky130_fd_sc_hd__mux2_1
X_25539_ _26974_/CLK _25539_/D vssd1 vssd1 vccd1 vccd1 _25539_/Q sky130_fd_sc_hd__dfxtp_1
X_13553_ _18645_/S _13553_/B vssd1 vssd1 vccd1 vccd1 _13554_/A sky130_fd_sc_hd__nor2_1
XFILLER_73_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19060_ _19060_/A vssd1 vssd1 vccd1 vccd1 _19060_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16272_ _16270_/X _16271_/X _16278_/S vssd1 vssd1 vccd1 vccd1 _16272_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13484_ _13484_/A vssd1 vssd1 vccd1 vccd1 _13791_/A sky130_fd_sc_hd__buf_2
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27209_ _27230_/CLK _27209_/D vssd1 vssd1 vccd1 vccd1 _27209_/Q sky130_fd_sc_hd__dfxtp_1
X_15223_ _14744_/A _26416_/Q _15120_/S _15222_/X vssd1 vssd1 vccd1 vccd1 _15223_/X
+ sky130_fd_sc_hd__o211a_1
X_18011_ _18377_/A _18895_/A _18010_/X _24986_/A vssd1 vssd1 vccd1 vccd1 _19253_/A
+ sky130_fd_sc_hd__o31ai_4
XFILLER_157_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15154_ _16161_/S vssd1 vssd1 vccd1 vccd1 _16395_/S sky130_fd_sc_hd__buf_4
Xoutput409 _25968_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_ack_o sky130_fd_sc_hd__buf_2
XFILLER_181_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14105_ _26069_/Q _14103_/X _14107_/A _14104_/X vssd1 vssd1 vccd1 vccd1 _14105_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15085_ _15085_/A vssd1 vssd1 vccd1 vccd1 _15085_/X sky130_fd_sc_hd__clkbuf_2
X_19962_ _19960_/Y _19961_/X _19957_/A _20323_/B vssd1 vssd1 vccd1 vccd1 _19962_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_268_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18913_ _25516_/Q _18556_/A _18557_/A _25548_/Q vssd1 vssd1 vccd1 vccd1 _18913_/X
+ sky130_fd_sc_hd__a22o_1
X_14036_ _15874_/A _15874_/B _15874_/C _14035_/X vssd1 vssd1 vccd1 vccd1 _14036_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_268_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19893_ _27110_/Q _19877_/X _19761_/X _19892_/X vssd1 vssd1 vccd1 vccd1 _19893_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_267_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18844_ _25736_/Q _19946_/A _18843_/D _25737_/Q vssd1 vssd1 vccd1 vccd1 _18844_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_110_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18775_ _18945_/A vssd1 vssd1 vccd1 vccd1 _18775_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15987_ _15818_/S _15986_/X _13998_/S vssd1 vssd1 vccd1 vccd1 _15987_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17726_ _17732_/A _17732_/B vssd1 vssd1 vccd1 vccd1 _18443_/A sky130_fd_sc_hd__nand2_1
XFILLER_270_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14938_ _25658_/Q _24351_/B _14613_/X vssd1 vssd1 vccd1 vccd1 _14938_/X sky130_fd_sc_hd__a21o_1
XFILLER_250_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17657_ _20689_/A vssd1 vssd1 vccd1 vccd1 _20687_/B sky130_fd_sc_hd__buf_6
X_14869_ _26125_/Q _26026_/Q _14876_/S vssd1 vssd1 vccd1 vccd1 _14869_/X sky130_fd_sc_hd__mux2_1
X_16608_ _19155_/A _19156_/B vssd1 vssd1 vccd1 vccd1 _16638_/A sky130_fd_sc_hd__xnor2_4
XFILLER_17_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17588_ _17995_/A vssd1 vssd1 vccd1 vccd1 _19455_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_250_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19327_ _19327_/A _19327_/B vssd1 vssd1 vccd1 vccd1 _19327_/X sky130_fd_sc_hd__xor2_1
XFILLER_204_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_16539_ _27294_/Q _26487_/Q _16541_/S vssd1 vssd1 vccd1 vccd1 _16539_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19258_ _27224_/Q _19258_/B vssd1 vssd1 vccd1 vccd1 _19258_/X sky130_fd_sc_hd__and2_1
XFILLER_192_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18209_ _17878_/X _17908_/X _18209_/S vssd1 vssd1 vccd1 vccd1 _18209_/X sky130_fd_sc_hd__mux2_1
X_19189_ _19191_/B _19189_/B vssd1 vssd1 vccd1 vccd1 _19189_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_157_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21220_ _21283_/A _17764_/X _21285_/A _25797_/Q _21251_/A vssd1 vssd1 vccd1 vccd1
+ _21220_/X sky130_fd_sc_hd__a221o_1
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21151_ _21154_/A _21151_/B vssd1 vssd1 vccd1 vccd1 _21152_/A sky130_fd_sc_hd__or2_1
X_20102_ _20102_/A _20102_/B vssd1 vssd1 vccd1 vccd1 _20102_/Y sky130_fd_sc_hd__nand2_1
XFILLER_160_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21082_ _21197_/A _21082_/B vssd1 vssd1 vccd1 vccd1 _21083_/A sky130_fd_sc_hd__or2_1
X_24910_ _24553_/A _24978_/B _24909_/X vssd1 vssd1 vccd1 vccd1 _24910_/Y sky130_fd_sc_hd__a21oi_1
X_20033_ _25738_/Q vssd1 vssd1 vccd1 vccd1 _20662_/A sky130_fd_sc_hd__buf_8
XFILLER_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25890_ _26609_/CLK _25890_/D vssd1 vssd1 vccd1 vccd1 _25890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24841_ _27116_/Q _24856_/B vssd1 vssd1 vccd1 vccd1 _24841_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24772_ _24781_/A _24772_/B vssd1 vssd1 vccd1 vccd1 _24772_/Y sky130_fd_sc_hd__nand2_4
X_21984_ _21984_/A vssd1 vssd1 vccd1 vccd1 _26105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26511_ _27287_/CLK _26511_/D vssd1 vssd1 vccd1 vccd1 _26511_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23723_ _23722_/X _26759_/Q _23732_/S vssd1 vssd1 vccd1 vccd1 _23724_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20935_ _23750_/A vssd1 vssd1 vccd1 vccd1 _20935_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26442_ _27281_/CLK _26442_/D vssd1 vssd1 vccd1 vccd1 _26442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23654_ _26734_/Q _23568_/X _23656_/S vssd1 vssd1 vccd1 vccd1 _23655_/A sky130_fd_sc_hd__mux2_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20866_ _23684_/A vssd1 vssd1 vccd1 vccd1 _20866_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22605_ _22593_/X _22604_/Y _22600_/X vssd1 vssd1 vccd1 vccd1 _26317_/D sky130_fd_sc_hd__a21oi_1
XFILLER_223_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26373_ _26468_/CLK _26373_/D vssd1 vssd1 vccd1 vccd1 _26373_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23585_ _26707_/Q _23584_/X _23588_/S vssd1 vssd1 vccd1 vccd1 _23586_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20797_ _20797_/A vssd1 vssd1 vccd1 vccd1 _25793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25324_ _27263_/Q _23684_/A _25332_/S vssd1 vssd1 vccd1 vccd1 _25325_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22536_ _22536_/A _22536_/B vssd1 vssd1 vccd1 vccd1 _22606_/A sky130_fd_sc_hd__nand2_2
XFILLER_210_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25255_ _25255_/A vssd1 vssd1 vccd1 vccd1 _27232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22467_ _26259_/Q _22470_/B vssd1 vssd1 vccd1 vccd1 _22467_/X sky130_fd_sc_hd__or2_1
X_24206_ _24216_/A _24213_/C vssd1 vssd1 vccd1 vccd1 _24206_/Y sky130_fd_sc_hd__nor2_1
XFILLER_185_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21418_ _21416_/X _21417_/X _21367_/X vssd1 vssd1 vccd1 vccd1 _21418_/X sky130_fd_sc_hd__a21o_1
XFILLER_182_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25186_ _24659_/B _25172_/X _25175_/X _27203_/Q _25179_/X vssd1 vssd1 vccd1 vccd1
+ _27203_/D sky130_fd_sc_hd__o221a_1
X_22398_ _22395_/A _22360_/C _22385_/X _22390_/Y _22395_/Y vssd1 vssd1 vccd1 vccd1
+ _22400_/A sky130_fd_sc_hd__o311a_1
XFILLER_191_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24137_ _24137_/A vssd1 vssd1 vccd1 vccd1 _26934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21349_ _26585_/Q _21349_/B _21562_/C _21562_/D vssd1 vssd1 vccd1 vccd1 _21350_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_162_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24068_ _26904_/Q _23600_/X _24070_/S vssd1 vssd1 vccd1 vccd1 _24069_/A sky130_fd_sc_hd__mux2_1
X_15910_ _13173_/A _15909_/X _13027_/A vssd1 vssd1 vccd1 vccd1 _15910_/X sky130_fd_sc_hd__o21a_1
XFILLER_2_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23019_ _23019_/A vssd1 vssd1 vccd1 vccd1 _23028_/S sky130_fd_sc_hd__buf_4
XFILLER_89_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16890_ _16890_/A vssd1 vssd1 vccd1 vccd1 _16939_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_265_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15841_ _26078_/Q _25883_/Q _15841_/S vssd1 vssd1 vccd1 vccd1 _15841_/X sky130_fd_sc_hd__mux2_1
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _27207_/Q _19258_/B vssd1 vssd1 vccd1 vccd1 _18560_/X sky130_fd_sc_hd__and2_1
XFILLER_18_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _25597_/Q _25585_/Q vssd1 vssd1 vccd1 vccd1 _14348_/S sky130_fd_sc_hd__and2b_2
X_15772_ _13351_/A _26111_/Q _26012_/Q _15197_/A _13359_/A vssd1 vssd1 vccd1 vccd1
+ _15772_/X sky130_fd_sc_hd__a221o_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ _19594_/A vssd1 vssd1 vccd1 vccd1 _18027_/A sky130_fd_sc_hd__clkbuf_4
X_26709_ _27253_/CLK _26709_/D vssd1 vssd1 vccd1 vccd1 _26709_/Q sky130_fd_sc_hd__dfxtp_1
X_14723_ _14723_/A vssd1 vssd1 vccd1 vccd1 _14724_/A sky130_fd_sc_hd__buf_4
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18491_ _18489_/S _18257_/X _18490_/X vssd1 vssd1 vccd1 vccd1 _18492_/B sky130_fd_sc_hd__a21oi_2
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _16310_/B vssd1 vssd1 vccd1 vccd1 _16243_/B sky130_fd_sc_hd__clkbuf_4
X_17442_ _17529_/A vssd1 vssd1 vccd1 vccd1 _20686_/A sky130_fd_sc_hd__buf_6
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _13065_/A _13601_/X _13604_/X _13142_/A vssd1 vssd1 vccd1 vccd1 _13605_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_177_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17373_ _17382_/A _17379_/C vssd1 vssd1 vccd1 vccd1 _17373_/Y sky130_fd_sc_hd__nor2_1
XFILLER_232_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14585_ _16451_/S vssd1 vssd1 vccd1 vccd1 _15012_/S sky130_fd_sc_hd__buf_2
XFILLER_158_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19112_ _19118_/B _19328_/S _18183_/X _19111_/Y vssd1 vssd1 vccd1 vccd1 _19112_/X
+ sky130_fd_sc_hd__a211o_1
X_13536_ _13534_/X _13535_/X _15606_/A vssd1 vssd1 vccd1 vccd1 _13536_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16324_ _16322_/X _16323_/X _16324_/S vssd1 vssd1 vccd1 vccd1 _16324_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16255_ _27318_/Q _26575_/Q _16255_/S vssd1 vssd1 vccd1 vccd1 _16255_/X sky130_fd_sc_hd__mux2_1
X_19043_ _15441_/X _18890_/X _19041_/Y _19042_/Y _18933_/X vssd1 vssd1 vccd1 vccd1
+ _19043_/X sky130_fd_sc_hd__a221o_2
X_13467_ _13467_/A vssd1 vssd1 vccd1 vccd1 _14786_/A sky130_fd_sc_hd__buf_6
XFILLER_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15206_ _16183_/S vssd1 vssd1 vccd1 vccd1 _16278_/S sky130_fd_sc_hd__buf_4
XFILLER_173_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16186_ _25818_/Q _27252_/Q _16186_/S vssd1 vssd1 vccd1 vccd1 _16186_/X sky130_fd_sc_hd__mux2_1
X_13398_ _12871_/Y _13393_/X _13397_/X _12943_/Y _12951_/X vssd1 vssd1 vccd1 vccd1
+ _13398_/Y sky130_fd_sc_hd__a221oi_2
X_15137_ _14601_/A _15134_/Y _15136_/X vssd1 vssd1 vccd1 vccd1 _15137_/X sky130_fd_sc_hd__o21a_1
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15068_ _16405_/A _15068_/B vssd1 vssd1 vccd1 vccd1 _15068_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19945_ _12674_/A _19914_/X _19944_/X vssd1 vssd1 vccd1 vccd1 _19950_/A sky130_fd_sc_hd__o21a_1
XFILLER_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14019_ _19798_/A _14124_/B vssd1 vssd1 vccd1 vccd1 _14019_/X sky130_fd_sc_hd__or2_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19876_ _20225_/A vssd1 vssd1 vccd1 vccd1 _19876_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18827_ _18827_/A vssd1 vssd1 vccd1 vccd1 _18827_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_283_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18758_ _27145_/Q _19465_/B vssd1 vssd1 vccd1 vccd1 _18758_/X sky130_fd_sc_hd__or2_1
XFILLER_271_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17709_ _17704_/S _19916_/A _17708_/X vssd1 vssd1 vccd1 vccd1 _17735_/B sky130_fd_sc_hd__o21ai_1
XFILLER_224_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18689_ _18679_/X _18680_/Y _18688_/X _18220_/X vssd1 vssd1 vccd1 vccd1 _18712_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20720_ _20484_/X _25758_/Q _20728_/S vssd1 vssd1 vccd1 vccd1 _20721_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20651_ _26271_/Q _20646_/X _20650_/X _20644_/X vssd1 vssd1 vccd1 vccd1 _25734_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23370_ _23370_/A vssd1 vssd1 vccd1 vccd1 _26621_/D sky130_fd_sc_hd__clkbuf_1
X_20582_ _20582_/A vssd1 vssd1 vccd1 vccd1 _25713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22321_ _26218_/Q _22310_/X _22316_/X _26319_/Q _22317_/X vssd1 vssd1 vccd1 vccd1
+ _22321_/X sky130_fd_sc_hd__a221o_1
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25040_ _20639_/A _25031_/X _25039_/X vssd1 vssd1 vccd1 vccd1 _25040_/Y sky130_fd_sc_hd__o21ai_1
X_22252_ _26196_/Q _22249_/X _22238_/X _26297_/Q _22241_/X vssd1 vssd1 vccd1 vccd1
+ _22252_/X sky130_fd_sc_hd__a221o_1
XFILLER_118_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21203_ _21203_/A vssd1 vssd1 vccd1 vccd1 _24457_/A sky130_fd_sc_hd__clkbuf_4
X_22183_ _26178_/Q _22171_/X _22179_/X input277/X _22172_/X vssd1 vssd1 vccd1 vccd1
+ _22183_/X sky130_fd_sc_hd__a221o_1
XFILLER_160_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21134_ _21134_/A vssd1 vssd1 vccd1 vccd1 _25917_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26991_ _26996_/CLK _26991_/D vssd1 vssd1 vccd1 vccd1 _26991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25942_ _27058_/CLK _25942_/D vssd1 vssd1 vccd1 vccd1 _25942_/Q sky130_fd_sc_hd__dfxtp_1
X_21065_ _25465_/S _21190_/A _16826_/A vssd1 vssd1 vccd1 vccd1 _21065_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_87_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20016_ _19725_/X _20014_/Y _20015_/X vssd1 vssd1 vccd1 vccd1 _20020_/A sky130_fd_sc_hd__a21o_1
XFILLER_280_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25873_ _27267_/CLK _25873_/D vssd1 vssd1 vccd1 vccd1 _25873_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_247_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24824_ _24822_/Y _24823_/X _24816_/X vssd1 vssd1 vccd1 vccd1 _27111_/D sky130_fd_sc_hd__a21oi_1
XFILLER_274_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24755_ _24781_/A _24755_/B vssd1 vssd1 vccd1 vccd1 _25147_/A sky130_fd_sc_hd__nand2_4
X_21967_ _21967_/A vssd1 vssd1 vccd1 vccd1 _26097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23706_ _23706_/A vssd1 vssd1 vccd1 vccd1 _23706_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20918_ _20918_/A vssd1 vssd1 vccd1 vccd1 _25843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24686_ _24703_/A _24686_/B vssd1 vssd1 vccd1 vccd1 _24686_/Y sky130_fd_sc_hd__nand2_1
X_21898_ _20504_/X _26067_/Q _21900_/S vssd1 vssd1 vccd1 vccd1 _21899_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26425_ _27264_/CLK _26425_/D vssd1 vssd1 vccd1 vccd1 _26425_/Q sky130_fd_sc_hd__dfxtp_2
X_23637_ _26726_/Q _23542_/X _23645_/S vssd1 vssd1 vccd1 vccd1 _23638_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20849_ _20849_/A vssd1 vssd1 vccd1 vccd1 _25820_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14370_ _13664_/A _26590_/Q _14296_/S _26330_/Q _13244_/A vssd1 vssd1 vccd1 vccd1
+ _14370_/X sky130_fd_sc_hd__o221a_1
X_26356_ _27291_/CLK _26356_/D vssd1 vssd1 vccd1 vccd1 _26356_/Q sky130_fd_sc_hd__dfxtp_2
X_23568_ _23568_/A vssd1 vssd1 vccd1 vccd1 _23568_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13321_ _13321_/A _13321_/B vssd1 vssd1 vccd1 vccd1 _13321_/X sky130_fd_sc_hd__or2_1
XFILLER_10_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25307_ _23766_/X _27256_/Q _25315_/S vssd1 vssd1 vccd1 vccd1 _25308_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22519_ _22519_/A vssd1 vssd1 vccd1 vccd1 _26283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26287_ _26292_/CLK _26287_/D vssd1 vssd1 vccd1 vccd1 _26287_/Q sky130_fd_sc_hd__dfxtp_1
X_23499_ _23499_/A vssd1 vssd1 vccd1 vccd1 _26679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ _17831_/A _16040_/B vssd1 vssd1 vccd1 vccd1 _18862_/S sky130_fd_sc_hd__and2_1
X_13252_ _13252_/A vssd1 vssd1 vccd1 vccd1 _13472_/A sky130_fd_sc_hd__buf_2
XFILLER_183_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25238_ _27225_/Q _25217_/X _25237_/X _25221_/X vssd1 vssd1 vccd1 vccd1 _27225_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25169_ _24772_/Y _25124_/X _25168_/Y _17339_/A vssd1 vssd1 vccd1 vccd1 _25169_/X
+ sky130_fd_sc_hd__a31o_1
X_13183_ _25596_/Q _15659_/A _16860_/A _16508_/S vssd1 vssd1 vccd1 vccd1 _17824_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_123_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17991_ _18602_/A vssd1 vssd1 vccd1 vccd1 _19454_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19730_ _20635_/A _19727_/X _19729_/X _19604_/X vssd1 vssd1 vccd1 vccd1 _19776_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_284_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16942_ _16942_/A _16942_/B vssd1 vssd1 vccd1 vccd1 _16943_/B sky130_fd_sc_hd__nor2_4
XFILLER_1_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19661_ _19943_/B vssd1 vssd1 vccd1 vccd1 _19661_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16873_ _16910_/A _16873_/B vssd1 vssd1 vccd1 vccd1 _16873_/X sky130_fd_sc_hd__or2_1
XFILLER_237_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18612_ _19957_/B _18508_/A _18509_/A _27176_/Q _18510_/A vssd1 vssd1 vccd1 vccd1
+ _18612_/X sky130_fd_sc_hd__a221o_1
XFILLER_253_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15824_ _26534_/Q _26142_/Q _15825_/S vssd1 vssd1 vccd1 vccd1 _15824_/X sky130_fd_sc_hd__mux2_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19592_ _19633_/C vssd1 vssd1 vccd1 vccd1 _25119_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ _17967_/X _18488_/Y _17988_/X vssd1 vssd1 vccd1 vccd1 _18544_/B sky130_fd_sc_hd__o21ai_1
X_12967_ _15532_/B vssd1 vssd1 vccd1 vccd1 _16212_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15755_ _13351_/A _26699_/Q _26827_/Q _13492_/X _13363_/A vssd1 vssd1 vccd1 vccd1
+ _15755_/X sky130_fd_sc_hd__a221o_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ _14706_/A vssd1 vssd1 vccd1 vccd1 _14706_/X sky130_fd_sc_hd__buf_6
X_18474_ _18474_/A _18474_/B vssd1 vssd1 vccd1 vccd1 _18474_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12898_ input126/X input161/X _14488_/S vssd1 vssd1 vccd1 vccd1 _12898_/X sky130_fd_sc_hd__mux2_8
XFILLER_205_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15686_ _16342_/S _15684_/X _15685_/X _14820_/A vssd1 vssd1 vccd1 vccd1 _15686_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17425_ _17427_/A _17427_/C _17424_/Y vssd1 vssd1 vccd1 vccd1 _25559_/D sky130_fd_sc_hd__o21a_1
XFILLER_178_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14637_ _14692_/S vssd1 vssd1 vccd1 vccd1 _14652_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17356_ _25538_/Q vssd1 vssd1 vccd1 vccd1 _17356_/X sky130_fd_sc_hd__buf_2
XFILLER_193_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14568_ _17983_/A _17805_/B vssd1 vssd1 vccd1 vccd1 _16707_/B sky130_fd_sc_hd__nor2_2
XFILLER_186_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27301_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_159_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16307_ _26513_/Q _26385_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _16307_/X sky130_fd_sc_hd__mux2_1
X_13519_ _14453_/A vssd1 vssd1 vccd1 vccd1 _13520_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_147_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14499_ _25797_/Q _27231_/Q _15895_/S vssd1 vssd1 vccd1 vccd1 _14499_/X sky130_fd_sc_hd__mux2_1
X_17287_ _25517_/Q vssd1 vssd1 vccd1 vccd1 _17287_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19026_ _27055_/Q _18811_/X _19023_/X _19025_/X _18823_/X vssd1 vssd1 vccd1 vccd1
+ _19026_/X sky130_fd_sc_hd__o221a_2
XFILLER_174_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16238_ _14877_/S _16235_/X _16237_/X _14661_/A vssd1 vssd1 vccd1 vccd1 _16238_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_173_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16169_ _15071_/A _16133_/Y _16168_/Y _15830_/A vssd1 vssd1 vccd1 vccd1 _16921_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_88_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19928_ _19908_/X _19927_/X _20079_/A _27111_/Q vssd1 vssd1 vccd1 vccd1 _19928_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_141_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19859_ _19980_/A _19981_/A vssd1 vssd1 vccd1 vccd1 _19860_/B sky130_fd_sc_hd__nor2_1
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22870_ _22870_/A vssd1 vssd1 vccd1 vccd1 _26414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_283_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21821_ _26040_/Q _20907_/X _21827_/S vssd1 vssd1 vccd1 vccd1 _21822_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24540_ _24457_/A _25491_/Q _17703_/X _24352_/X vssd1 vssd1 vccd1 vccd1 _24541_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_24_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21752_ _20546_/X _26010_/Q _21754_/S vssd1 vssd1 vccd1 vccd1 _21753_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20703_ _20703_/A _20703_/B vssd1 vssd1 vccd1 vccd1 _20703_/Y sky130_fd_sc_hd__nand2_1
X_24471_ _27023_/Q _24448_/X _24469_/Y _24470_/X vssd1 vssd1 vccd1 vccd1 _27023_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21683_ _25981_/Q input193/X _21685_/S vssd1 vssd1 vccd1 vccd1 _21684_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26210_ _26322_/CLK _26210_/D vssd1 vssd1 vccd1 vccd1 _26210_/Q sky130_fd_sc_hd__dfxtp_1
X_23422_ _26645_/Q _23117_/X _23430_/S vssd1 vssd1 vccd1 vccd1 _23423_/A sky130_fd_sc_hd__mux2_1
X_20634_ _20674_/A vssd1 vssd1 vccd1 vccd1 _20643_/B sky130_fd_sc_hd__clkbuf_1
X_27190_ _27196_/CLK _27190_/D vssd1 vssd1 vccd1 vccd1 _27190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26141_ _26468_/CLK _26141_/D vssd1 vssd1 vccd1 vccd1 _26141_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_138_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23353_ _20605_/X _26615_/Q _23357_/S vssd1 vssd1 vccd1 vccd1 _23354_/A sky130_fd_sc_hd__mux2_1
X_20565_ _20565_/A vssd1 vssd1 vccd1 vccd1 _25709_/D sky130_fd_sc_hd__clkbuf_1
X_22304_ _22428_/A vssd1 vssd1 vccd1 vccd1 _22304_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26072_ _26601_/CLK _26072_/D vssd1 vssd1 vccd1 vccd1 _26072_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_153_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23284_ _23284_/A vssd1 vssd1 vccd1 vccd1 _26584_/D sky130_fd_sc_hd__clkbuf_1
X_20496_ _23690_/A vssd1 vssd1 vccd1 vccd1 _20496_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25023_ _27170_/Q _25000_/X _25022_/X vssd1 vssd1 vccd1 vccd1 _27170_/D sky130_fd_sc_hd__o21ba_1
XFILLER_118_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22235_ _22269_/A vssd1 vssd1 vccd1 vccd1 _22235_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22166_ _22166_/A _22207_/S vssd1 vssd1 vccd1 vccd1 _22166_/X sky130_fd_sc_hd__or2b_1
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21117_ _25913_/Q _21112_/X _21113_/X input12/X vssd1 vssd1 vccd1 vccd1 _21118_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_278_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26974_ _26974_/CLK _26974_/D vssd1 vssd1 vccd1 vccd1 _26974_/Q sky130_fd_sc_hd__dfxtp_1
X_22097_ _26156_/Q _20961_/X _22099_/S vssd1 vssd1 vccd1 vccd1 _22098_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21048_ _25893_/Q _20948_/X _21048_/S vssd1 vssd1 vccd1 vccd1 _21049_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25925_ _27213_/CLK _25925_/D vssd1 vssd1 vccd1 vccd1 _25925_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_75_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13870_ _27270_/Q _26463_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _13870_/X sky130_fd_sc_hd__mux2_1
XFILLER_235_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25856_ _26900_/CLK _25856_/D vssd1 vssd1 vccd1 vccd1 _25856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12821_ _17224_/A _21320_/A _21300_/A vssd1 vssd1 vccd1 vccd1 _12973_/A sky130_fd_sc_hd__or3b_1
XFILLER_234_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24807_ _20639_/A _24789_/X _24668_/Y _24791_/X vssd1 vssd1 vccd1 vccd1 _24807_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_234_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22999_ _22999_/A vssd1 vssd1 vccd1 vccd1 _26471_/D sky130_fd_sc_hd__clkbuf_1
X_25787_ _27324_/CLK _25787_/D vssd1 vssd1 vccd1 vccd1 _25787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12752_ _25584_/Q vssd1 vssd1 vccd1 vccd1 _13945_/A sky130_fd_sc_hd__buf_2
X_15540_ _26861_/Q _25775_/Q _15540_/S vssd1 vssd1 vccd1 vccd1 _15540_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24738_ _24742_/A _24738_/B vssd1 vssd1 vccd1 vccd1 _27091_/D sky130_fd_sc_hd__nor2_1
XFILLER_131_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15471_ _26346_/Q _26606_/Q _15471_/S vssd1 vssd1 vccd1 vccd1 _15471_/X sky130_fd_sc_hd__mux2_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _13001_/A vssd1 vssd1 vccd1 vccd1 _13641_/A sky130_fd_sc_hd__buf_4
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24669_ _27075_/Q _24657_/X _24668_/Y _24660_/X vssd1 vssd1 vccd1 vccd1 _24670_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _12673_/A _27296_/Q _26553_/Q _14273_/B _13022_/A vssd1 vssd1 vccd1 vccd1
+ _14422_/X sky130_fd_sc_hd__o221a_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _17210_/A vssd1 vssd1 vccd1 vccd1 _17529_/A sky130_fd_sc_hd__buf_2
XFILLER_202_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26408_ _26604_/CLK _26408_/D vssd1 vssd1 vccd1 vccd1 _26408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18190_ _18684_/S _18344_/A _17984_/Y vssd1 vssd1 vccd1 vccd1 _18799_/B sky130_fd_sc_hd__a21o_1
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14353_ _13630_/A _14349_/X _14352_/X _14331_/A vssd1 vssd1 vccd1 vccd1 _14353_/X
+ sky130_fd_sc_hd__o22a_1
X_17141_ _25476_/Q _17105_/X _17107_/X _25573_/Q vssd1 vssd1 vccd1 vccd1 _17142_/B
+ sky130_fd_sc_hd__a22o_1
X_26339_ _26467_/CLK _26339_/D vssd1 vssd1 vccd1 vccd1 _26339_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13304_ _13304_/A vssd1 vssd1 vccd1 vccd1 _13305_/A sky130_fd_sc_hd__buf_4
XFILLER_144_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17072_ _26237_/Q vssd1 vssd1 vccd1 vccd1 _22350_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_183_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14284_ _13105_/B _14362_/B _14283_/Y vssd1 vssd1 vccd1 vccd1 _14566_/B sky130_fd_sc_hd__a21oi_4
XFILLER_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16023_ _13814_/X _16020_/X _16022_/X _13475_/A vssd1 vssd1 vccd1 vccd1 _16023_/X
+ sky130_fd_sc_hd__o211a_1
X_13235_ _26631_/Q _26727_/Q _15662_/S vssd1 vssd1 vccd1 vccd1 _13236_/B sky130_fd_sc_hd__mux2_1
XFILLER_7_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13166_ _14355_/A vssd1 vssd1 vccd1 vccd1 _14523_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_153_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27093_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_269_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13097_ _13185_/A _25586_/Q vssd1 vssd1 vccd1 vccd1 _14352_/S sky130_fd_sc_hd__nand2_4
X_17974_ _18042_/S _18186_/A _17886_/Y vssd1 vssd1 vccd1 vccd1 _17974_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19713_ _19779_/A vssd1 vssd1 vccd1 vccd1 _19926_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16925_ _16925_/A vssd1 vssd1 vccd1 vccd1 _16925_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19644_ _19646_/A vssd1 vssd1 vccd1 vccd1 _19870_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_66_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16856_ _16836_/X _16852_/X _16855_/Y _16842_/X vssd1 vssd1 vccd1 vccd1 _16857_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_253_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15807_ _27277_/Q _26470_/Q _15807_/S vssd1 vssd1 vccd1 vccd1 _15807_/X sky130_fd_sc_hd__mux2_1
X_19575_ _19575_/A _19575_/B vssd1 vssd1 vccd1 vccd1 _19576_/B sky130_fd_sc_hd__nor2_1
XFILLER_65_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16787_ _16853_/A vssd1 vssd1 vccd1 vccd1 _16973_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_206_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13999_ _13985_/X _13989_/X _13998_/X _13608_/X _13107_/A vssd1 vssd1 vccd1 vccd1
+ _13999_/X sky130_fd_sc_hd__a221o_1
XFILLER_92_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18526_ _19268_/B _19824_/A vssd1 vssd1 vccd1 vccd1 _18526_/X sky130_fd_sc_hd__and2b_1
X_15738_ _26343_/Q _26603_/Q _15989_/S vssd1 vssd1 vccd1 vccd1 _15738_/X sky130_fd_sc_hd__mux2_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18457_ _27166_/Q _18121_/A _18121_/B _18456_/X vssd1 vssd1 vccd1 vccd1 _18457_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15669_ _26080_/Q _25885_/Q _16277_/S vssd1 vssd1 vccd1 vccd1 _15669_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17408_ _17408_/A _25554_/Q _17408_/C vssd1 vssd1 vccd1 vccd1 _17410_/B sky130_fd_sc_hd__and3_1
XFILLER_194_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18388_ _18811_/A vssd1 vssd1 vccd1 vccd1 _18503_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17339_ _17339_/A vssd1 vssd1 vccd1 vccd1 _17380_/A sky130_fd_sc_hd__buf_2
XFILLER_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20350_ _19763_/X _20348_/Y _20349_/X _20707_/D vssd1 vssd1 vccd1 vccd1 _20350_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19009_ _19252_/A vssd1 vssd1 vccd1 vccd1 _19317_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20281_ _20280_/B _20279_/Y _19589_/B _20280_/Y vssd1 vssd1 vccd1 vccd1 _20281_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22020_ _22020_/A vssd1 vssd1 vccd1 vccd1 _26121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_283_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23971_ _23971_/A vssd1 vssd1 vccd1 vccd1 _26860_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22922_ _22922_/A vssd1 vssd1 vccd1 vccd1 _26437_/D sky130_fd_sc_hd__clkbuf_1
X_25710_ _26531_/CLK _25710_/D vssd1 vssd1 vccd1 vccd1 _25710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26690_ _26880_/CLK _26690_/D vssd1 vssd1 vccd1 vccd1 _26690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25641_ _25660_/CLK _25641_/D vssd1 vssd1 vccd1 vccd1 _25641_/Q sky130_fd_sc_hd__dfxtp_1
X_22853_ _22875_/A vssd1 vssd1 vccd1 vccd1 _22862_/S sky130_fd_sc_hd__buf_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21804_ _21804_/A vssd1 vssd1 vccd1 vccd1 _26032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25572_ _25590_/CLK _25572_/D vssd1 vssd1 vccd1 vccd1 _25572_/Q sky130_fd_sc_hd__dfxtp_4
X_22784_ _22784_/A vssd1 vssd1 vccd1 vccd1 _26376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24523_ _24551_/A vssd1 vssd1 vccd1 vccd1 _24523_/X sky130_fd_sc_hd__clkbuf_2
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27311_ _27311_/CLK _27311_/D vssd1 vssd1 vccd1 vccd1 _27311_/Q sky130_fd_sc_hd__dfxtp_1
X_21735_ _20512_/X _26002_/Q _21743_/S vssd1 vssd1 vccd1 vccd1 _21736_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24454_ _24454_/A vssd1 vssd1 vccd1 vccd1 _24454_/X sky130_fd_sc_hd__buf_4
X_27242_ _27306_/CLK _27242_/D vssd1 vssd1 vccd1 vccd1 _27242_/Q sky130_fd_sc_hd__dfxtp_1
X_21666_ _25973_/Q input208/X _21674_/S vssd1 vssd1 vccd1 vccd1 _21667_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23405_ _23405_/A vssd1 vssd1 vccd1 vccd1 _26637_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20617_ _23782_/A vssd1 vssd1 vccd1 vccd1 _20617_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_27173_ _27173_/CLK _27173_/D vssd1 vssd1 vccd1 vccd1 _27173_/Q sky130_fd_sc_hd__dfxtp_1
X_24385_ _26297_/Q _24382_/X _24383_/X input241/X _24384_/X vssd1 vssd1 vccd1 vccd1
+ _24385_/X sky130_fd_sc_hd__a221o_1
X_21597_ _21597_/A vssd1 vssd1 vccd1 vccd1 _21597_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26124_ _27291_/CLK _26124_/D vssd1 vssd1 vccd1 vccd1 _26124_/Q sky130_fd_sc_hd__dfxtp_2
X_23336_ _23336_/A vssd1 vssd1 vccd1 vccd1 _26607_/D sky130_fd_sc_hd__clkbuf_1
X_20548_ _20548_/A vssd1 vssd1 vccd1 vccd1 _25705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26055_ _26483_/CLK _26055_/D vssd1 vssd1 vccd1 vccd1 _26055_/Q sky130_fd_sc_hd__dfxtp_1
X_23267_ _23267_/A vssd1 vssd1 vccd1 vccd1 _26576_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20479_ _20478_/A _20478_/B _20478_/Y _19787_/A vssd1 vssd1 vccd1 vccd1 _20480_/B
+ sky130_fd_sc_hd__a211o_1
X_13020_ _14253_/S vssd1 vssd1 vccd1 vccd1 _15825_/S sky130_fd_sc_hd__clkbuf_4
X_25006_ _16855_/A _25004_/X _25756_/Q _25005_/X vssd1 vssd1 vccd1 vccd1 _25006_/X
+ sky130_fd_sc_hd__a211o_1
X_22218_ _26188_/Q _22200_/X _22215_/X _22217_/X vssd1 vssd1 vccd1 vccd1 _26188_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23198_ _23198_/A vssd1 vssd1 vccd1 vccd1 _26545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22149_ _26168_/Q _22136_/X _22147_/X _22148_/X vssd1 vssd1 vccd1 vccd1 _26168_/D
+ sky130_fd_sc_hd__o211a_1
X_26957_ _26992_/CLK _26957_/D vssd1 vssd1 vccd1 vccd1 _26957_/Q sky130_fd_sc_hd__dfxtp_1
X_14971_ _25897_/Q _15026_/B vssd1 vssd1 vccd1 vccd1 _14971_/X sky130_fd_sc_hd__or2_1
XFILLER_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16710_ _25664_/Q vssd1 vssd1 vccd1 vccd1 _22478_/A sky130_fd_sc_hd__buf_2
XFILLER_120_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13922_ _25924_/Q _13922_/B vssd1 vssd1 vccd1 vccd1 _13922_/Y sky130_fd_sc_hd__nor2_1
X_25908_ _27122_/CLK _25908_/D vssd1 vssd1 vccd1 vccd1 _25908_/Q sky130_fd_sc_hd__dfxtp_4
X_17690_ _17691_/A _17470_/A _17689_/X vssd1 vssd1 vccd1 vccd1 _17747_/B sky130_fd_sc_hd__o21ai_1
X_26888_ _27310_/CLK _26888_/D vssd1 vssd1 vccd1 vccd1 _26888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16641_ _16641_/A _21075_/B vssd1 vssd1 vccd1 vccd1 _21070_/A sky130_fd_sc_hd__nand2_8
XFILLER_274_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25839_ _26601_/CLK _25839_/D vssd1 vssd1 vccd1 vccd1 _25839_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_263_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13853_ _13180_/A _19824_/A _13852_/X vssd1 vssd1 vccd1 vccd1 _17797_/B sky130_fd_sc_hd__o21a_2
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_406 _17044_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_417 _17009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19360_ _16561_/B _17997_/A _19359_/Y _16560_/A vssd1 vssd1 vccd1 vccd1 _19360_/X
+ sky130_fd_sc_hd__a22o_1
X_12804_ _14188_/A _14189_/A _12803_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _19076_/A
+ sky130_fd_sc_hd__a211o_4
X_16572_ _19237_/A _16572_/B vssd1 vssd1 vccd1 vccd1 _16573_/B sky130_fd_sc_hd__nor2_1
XINSDIODE2_428 _12781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13784_ _26628_/Q _26724_/Q _15914_/S vssd1 vssd1 vccd1 vccd1 _13784_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_439 _25729_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18311_ _18858_/S _18256_/X _18271_/X vssd1 vssd1 vccd1 vccd1 _18311_/X sky130_fd_sc_hd__o21a_1
XFILLER_231_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15523_ _15495_/Y _15505_/Y _15522_/Y _13314_/A _13638_/X vssd1 vssd1 vccd1 vccd1
+ _15523_/Y sky130_fd_sc_hd__o221ai_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12735_ _14453_/A vssd1 vssd1 vccd1 vccd1 _12736_/A sky130_fd_sc_hd__buf_2
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19291_ _19277_/A _19276_/B _17785_/X vssd1 vssd1 vccd1 vccd1 _19292_/B sky130_fd_sc_hd__o21ai_2
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _27040_/Q _19055_/A _18237_/X _18241_/X _19066_/A vssd1 vssd1 vccd1 vccd1
+ _18242_/X sky130_fd_sc_hd__o221a_2
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _25710_/Q _15468_/B vssd1 vssd1 vccd1 vccd1 _15454_/X sky130_fd_sc_hd__or2_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14405_ _25903_/Q _12902_/A _14404_/Y _14486_/A vssd1 vssd1 vccd1 vccd1 _14405_/X
+ sky130_fd_sc_hd__o211a_1
X_18173_ _18465_/A vssd1 vssd1 vccd1 vccd1 _18830_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15385_ _15379_/X _15381_/X _15384_/X _16328_/A _12704_/A vssd1 vssd1 vccd1 vccd1
+ _15385_/X sky130_fd_sc_hd__o221a_1
XFILLER_128_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17124_ _25470_/Q _17114_/X _17123_/X _17120_/X vssd1 vssd1 vccd1 vccd1 _25470_/D
+ sky130_fd_sc_hd__o211a_1
X_14336_ _13083_/A _26458_/Q _14265_/S _27265_/Q _14331_/A vssd1 vssd1 vccd1 vccd1
+ _14336_/X sky130_fd_sc_hd__o221a_1
XFILLER_190_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14267_ _13889_/A _14265_/X _14266_/X vssd1 vssd1 vccd1 vccd1 _14267_/X sky130_fd_sc_hd__o21a_1
X_17055_ _17055_/A _17055_/B _17055_/C _17055_/D vssd1 vssd1 vccd1 vccd1 _17056_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_100_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16006_ _16006_/A _16006_/B vssd1 vssd1 vccd1 vccd1 _16006_/X sky130_fd_sc_hd__or2_1
X_13218_ _13358_/A vssd1 vssd1 vccd1 vccd1 _15916_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_171_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14198_ _26784_/Q _26428_/Q _15858_/S vssd1 vssd1 vccd1 vccd1 _14198_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13149_ _14004_/S vssd1 vssd1 vccd1 vccd1 _15796_/S sky130_fd_sc_hd__clkbuf_4
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _15528_/B _16038_/B _17957_/S vssd1 vssd1 vccd1 vccd1 _17957_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16908_ _16908_/A _16927_/B vssd1 vssd1 vccd1 vccd1 _16963_/C sky130_fd_sc_hd__nor2_1
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17888_ _18063_/S vssd1 vssd1 vccd1 vccd1 _18044_/S sky130_fd_sc_hd__buf_2
XFILLER_266_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19627_ _27054_/Q _21264_/A input178/X _19622_/X _19626_/X vssd1 vssd1 vccd1 vccd1
+ _19628_/C sky130_fd_sc_hd__a311o_1
XFILLER_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16839_ _16839_/A _16859_/A vssd1 vssd1 vccd1 vccd1 _16840_/A sky130_fd_sc_hd__nand2_2
XFILLER_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19558_ _19551_/X _19308_/X _19557_/X _19555_/X vssd1 vssd1 vccd1 vccd1 _25656_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_241_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_50_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27249_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18509_ _18509_/A vssd1 vssd1 vccd1 vccd1 _18509_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19489_ _19541_/A vssd1 vssd1 vccd1 vccd1 _19489_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21520_ _21515_/Y _21519_/X _21492_/X vssd1 vssd1 vccd1 vccd1 _21520_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_33_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21451_ _21581_/A vssd1 vssd1 vccd1 vccd1 _21451_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20402_ _19374_/A _18092_/A _19382_/X _20328_/X vssd1 vssd1 vccd1 vccd1 _20402_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_119_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24170_ _24222_/A _24170_/B _24175_/C vssd1 vssd1 vccd1 vccd1 _26947_/D sky130_fd_sc_hd__nor3_1
XFILLER_175_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21382_ _20650_/A _21343_/X _21350_/X _21381_/X vssd1 vssd1 vccd1 vccd1 _21382_/X
+ sky130_fd_sc_hd__o211a_1
X_23121_ _23594_/A vssd1 vssd1 vccd1 vccd1 _23121_/X sky130_fd_sc_hd__clkbuf_2
X_20333_ _19766_/X _20332_/Y _20015_/X vssd1 vssd1 vccd1 vccd1 _20337_/A sky130_fd_sc_hd__a21o_1
X_23052_ _23052_/A vssd1 vssd1 vccd1 vccd1 _26492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20264_ _25682_/Q _20286_/C vssd1 vssd1 vccd1 vccd1 _20265_/C sky130_fd_sc_hd__or2_1
XFILLER_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22003_ _26114_/Q _20929_/X _22005_/S vssd1 vssd1 vccd1 vccd1 _22004_/A sky130_fd_sc_hd__mux2_1
XTAP_5306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20195_ _20141_/B _19115_/Y _19911_/X _20194_/Y vssd1 vssd1 vccd1 vccd1 _20195_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput106 dout0[9] vssd1 vssd1 vccd1 vccd1 input106/X sky130_fd_sc_hd__clkbuf_2
XTAP_5328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput117 dout1[19] vssd1 vssd1 vccd1 vccd1 input117/X sky130_fd_sc_hd__clkbuf_1
X_26811_ _26843_/CLK _26811_/D vssd1 vssd1 vccd1 vccd1 _26811_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput128 dout1[29] vssd1 vssd1 vccd1 vccd1 input128/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput139 dout1[39] vssd1 vssd1 vccd1 vccd1 input139/X sky130_fd_sc_hd__clkbuf_2
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26742_ _27321_/CLK _26742_/D vssd1 vssd1 vccd1 vccd1 _26742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23954_ _26853_/Q _23539_/X _23954_/S vssd1 vssd1 vccd1 vccd1 _23955_/A sky130_fd_sc_hd__mux2_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22905_ _22905_/A vssd1 vssd1 vccd1 vccd1 _26429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_256_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23885_ _23718_/X _26822_/Q _23893_/S vssd1 vssd1 vccd1 vccd1 _23886_/A sky130_fd_sc_hd__mux2_1
X_26673_ _26673_/CLK _26673_/D vssd1 vssd1 vccd1 vccd1 _26673_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22836_ _26399_/Q _22666_/X _22840_/S vssd1 vssd1 vccd1 vccd1 _22837_/A sky130_fd_sc_hd__mux2_1
XFILLER_260_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25624_ _25624_/CLK _25624_/D vssd1 vssd1 vccd1 vccd1 _25624_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22767_ _26369_/Q _22672_/X _22767_/S vssd1 vssd1 vccd1 vccd1 _22768_/A sky130_fd_sc_hd__mux2_1
X_25555_ _25992_/CLK _25555_/D vssd1 vssd1 vccd1 vccd1 _25555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24506_ _24506_/A vssd1 vssd1 vccd1 vccd1 _24506_/X sky130_fd_sc_hd__clkbuf_2
X_21718_ _21718_/A _21718_/B _21718_/C vssd1 vssd1 vccd1 vccd1 _21719_/A sky130_fd_sc_hd__and3_1
XFILLER_40_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25486_ _26843_/CLK _25486_/D vssd1 vssd1 vccd1 vccd1 _25486_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22698_ _23741_/A vssd1 vssd1 vccd1 vccd1 _22698_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27225_ _27227_/CLK _27225_/D vssd1 vssd1 vccd1 vccd1 _27225_/Q sky130_fd_sc_hd__dfxtp_1
X_24437_ _26306_/Q _24382_/X _24383_/X input219/X _24404_/X vssd1 vssd1 vccd1 vccd1
+ _24437_/X sky130_fd_sc_hd__a221o_1
X_21649_ _21645_/Y _21648_/X _21202_/A vssd1 vssd1 vccd1 vccd1 _21649_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_166_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15170_ _15167_/X _26900_/Q _26772_/Q _15030_/S _15169_/X vssd1 vssd1 vccd1 vccd1
+ _15170_/X sky130_fd_sc_hd__a221o_1
XFILLER_184_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24368_ _24372_/A _24550_/A vssd1 vssd1 vccd1 vccd1 _24368_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27156_ _27156_/CLK _27156_/D vssd1 vssd1 vccd1 vccd1 _27156_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_126_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14121_ _13162_/A _14106_/X _14112_/X _14355_/A _14120_/X vssd1 vssd1 vccd1 vccd1
+ _14121_/X sky130_fd_sc_hd__a311o_1
X_26107_ _26467_/CLK _26107_/D vssd1 vssd1 vccd1 vccd1 _26107_/Q sky130_fd_sc_hd__dfxtp_4
X_23319_ _23319_/A vssd1 vssd1 vccd1 vccd1 _26599_/D sky130_fd_sc_hd__clkbuf_1
X_27087_ _27087_/CLK _27087_/D vssd1 vssd1 vccd1 vccd1 _27087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24299_ _26990_/Q _24301_/C _24298_/Y vssd1 vssd1 vccd1 vccd1 _26990_/D sky130_fd_sc_hd__o21a_1
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14052_ _26913_/Q _26397_/Q _14544_/S vssd1 vssd1 vccd1 vccd1 _14052_/X sky130_fd_sc_hd__mux2_1
X_26038_ _26595_/CLK _26038_/D vssd1 vssd1 vccd1 vccd1 _26038_/Q sky130_fd_sc_hd__dfxtp_2
X_13003_ _13197_/A _12989_/A _13015_/A _13002_/A vssd1 vssd1 vccd1 vccd1 _13003_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_134_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_18860_ _18362_/X _18858_/X _18859_/Y _18321_/A vssd1 vssd1 vccd1 vccd1 _18864_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17811_ _18184_/B _18184_/C _18184_/A vssd1 vssd1 vccd1 vccd1 _18251_/C sky130_fd_sc_hd__a21o_1
X_18791_ _25610_/Q _18719_/X _18789_/X _18790_/X vssd1 vssd1 vccd1 vccd1 _25610_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17742_ _18454_/A vssd1 vssd1 vccd1 vccd1 _17742_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14954_ _12776_/A _26712_/Q _26840_/Q _14963_/S _16484_/A vssd1 vssd1 vccd1 vccd1
+ _14954_/X sky130_fd_sc_hd__a221o_1
XTAP_5884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13905_ _14317_/B vssd1 vssd1 vccd1 vccd1 _15948_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_208_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17673_ _18554_/A vssd1 vssd1 vccd1 vccd1 _17673_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14885_ _14593_/A _14839_/Y _14884_/Y _15079_/A vssd1 vssd1 vccd1 vccd1 _14886_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_35_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19412_ _18895_/X _19396_/X _19411_/X _18927_/X vssd1 vssd1 vccd1 vccd1 _19412_/X
+ sky130_fd_sc_hd__a22o_1
X_16624_ _18975_/A _16624_/B vssd1 vssd1 vccd1 vccd1 _16637_/C sky130_fd_sc_hd__xnor2_4
XFILLER_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_203 _14480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13836_ _13835_/X _26915_/Q _26399_/Q _15514_/S _13814_/X vssd1 vssd1 vccd1 vccd1
+ _13836_/X sky130_fd_sc_hd__a221o_1
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_214 _16901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_225 _23549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_236 _19046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_247 _19256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19343_ _18912_/A _19341_/Y _17774_/X vssd1 vssd1 vccd1 vccd1 _19343_/X sky130_fd_sc_hd__o21a_1
XINSDIODE2_258 _24630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16555_ _16560_/A _16562_/A _16561_/B vssd1 vssd1 vccd1 vccd1 _16558_/A sky130_fd_sc_hd__a21o_1
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13767_ _26916_/Q _26400_/Q _15915_/S vssd1 vssd1 vccd1 vccd1 _13767_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_269 _24335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15506_ _15937_/S vssd1 vssd1 vccd1 vccd1 _16113_/A sky130_fd_sc_hd__buf_4
XFILLER_189_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19274_ _16372_/A _18366_/X _19272_/Y _16794_/B _19273_/Y vssd1 vssd1 vccd1 vccd1
+ _19274_/X sky130_fd_sc_hd__o221a_1
X_12718_ _14956_/A vssd1 vssd1 vccd1 vccd1 _16481_/A sky130_fd_sc_hd__buf_6
XFILLER_188_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16486_ _12760_/B _16482_/X _16485_/X vssd1 vssd1 vccd1 vccd1 _16486_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_231_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13698_ _13698_/A vssd1 vssd1 vccd1 vccd1 _15547_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_188_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18225_ _18336_/A _18225_/B vssd1 vssd1 vccd1 vccd1 _18226_/A sky130_fd_sc_hd__and2_1
XFILLER_248_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15437_ _19105_/S vssd1 vssd1 vccd1 vccd1 _15439_/A sky130_fd_sc_hd__inv_2
XFILLER_50_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18156_ _18440_/A vssd1 vssd1 vccd1 vccd1 _18808_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15368_ _15142_/A _15365_/X _15367_/X _15040_/A vssd1 vssd1 vccd1 vccd1 _15368_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17107_ _17145_/A vssd1 vssd1 vccd1 vccd1 _17107_/X sky130_fd_sc_hd__buf_2
XFILLER_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14319_ _18317_/S _14567_/A vssd1 vssd1 vccd1 vccd1 _16713_/A sky130_fd_sc_hd__nor2_2
XFILLER_144_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18087_ _18035_/X _18037_/X _18039_/X _18086_/X vssd1 vssd1 vccd1 vccd1 _18087_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15299_ _26118_/Q _26019_/Q _15299_/S vssd1 vssd1 vccd1 vccd1 _15299_/X sky130_fd_sc_hd__mux2_1
XFILLER_264_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17038_ _17035_/X _16930_/B _17032_/X input229/X vssd1 vssd1 vccd1 vccd1 _17038_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_172_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18989_ _27150_/Q _19465_/B vssd1 vssd1 vccd1 vccd1 _18989_/X sky130_fd_sc_hd__or2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20951_ _23766_/A vssd1 vssd1 vccd1 vccd1 _20951_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23670_ _26741_/Q _23590_/X _23678_/S vssd1 vssd1 vccd1 vccd1 _23671_/A sky130_fd_sc_hd__mux2_1
X_20882_ _25832_/Q _20881_/X _20885_/S vssd1 vssd1 vccd1 vccd1 _20883_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22621_ _22567_/A _22620_/Y _22614_/X vssd1 vssd1 vccd1 vccd1 _26323_/D sky130_fd_sc_hd__a21oi_1
XFILLER_179_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25340_ _25340_/A vssd1 vssd1 vccd1 vccd1 _27270_/D sky130_fd_sc_hd__clkbuf_1
X_22552_ _22538_/X _22551_/Y _22547_/X vssd1 vssd1 vccd1 vccd1 _26297_/D sky130_fd_sc_hd__a21oi_1
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21503_ _21488_/X _21462_/X _21502_/Y _21451_/X vssd1 vssd1 vccd1 vccd1 _21503_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_179_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25271_ _23715_/X _27240_/Q _25271_/S vssd1 vssd1 vccd1 vccd1 _25272_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22483_ _22483_/A _22491_/B vssd1 vssd1 vccd1 vccd1 _22484_/A sky130_fd_sc_hd__and2_1
XFILLER_158_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24222_ _24222_/A _24222_/B _24227_/C vssd1 vssd1 vccd1 vccd1 _26964_/D sky130_fd_sc_hd__nor3_1
X_27010_ _27044_/CLK _27010_/D vssd1 vssd1 vccd1 vccd1 _27010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21434_ _21429_/X _21432_/X _21433_/X vssd1 vssd1 vccd1 vccd1 _21434_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24153_ _24222_/A hold5/X _24157_/C vssd1 vssd1 vccd1 vccd1 _26941_/D sky130_fd_sc_hd__nor3_1
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21365_ _21587_/A vssd1 vssd1 vccd1 vccd1 _21365_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23104_ _23104_/A vssd1 vssd1 vccd1 vccd1 _26508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20316_ _22522_/A _20334_/C _20315_/Y vssd1 vssd1 vccd1 vccd1 _20317_/C sky130_fd_sc_hd__a21oi_1
X_24084_ _24084_/A vssd1 vssd1 vccd1 vccd1 _26910_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21296_ _21309_/A vssd1 vssd1 vccd1 vccd1 _21556_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23035_ _23788_/B vssd1 vssd1 vccd1 vccd1 _25393_/A sky130_fd_sc_hd__buf_4
X_20247_ _22516_/A _20225_/X _20239_/Y _20246_/X _20223_/X vssd1 vssd1 vccd1 vccd1
+ _25681_/D sky130_fd_sc_hd__o221a_1
XFILLER_27_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20178_ _27120_/Q _20079_/X _20112_/X _20177_/Y vssd1 vssd1 vccd1 vccd1 _20178_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24986_ _24986_/A _24986_/B vssd1 vssd1 vccd1 vccd1 _24986_/Y sky130_fd_sc_hd__nand2_4
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26725_ _26916_/CLK _26725_/D vssd1 vssd1 vccd1 vccd1 _26725_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23937_ _26845_/Q _23514_/X _23943_/S vssd1 vssd1 vccd1 vccd1 _23938_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26656_ _26880_/CLK _26656_/D vssd1 vssd1 vccd1 vccd1 _26656_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ _26358_/Q _26618_/Q _14699_/S vssd1 vssd1 vccd1 vccd1 _14670_/X sky130_fd_sc_hd__mux2_1
XFILLER_233_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23868_ _23868_/A vssd1 vssd1 vccd1 vccd1 _26814_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13621_ _14089_/S vssd1 vssd1 vccd1 vccd1 _15720_/S sky130_fd_sc_hd__clkbuf_4
X_25607_ _25607_/CLK _25607_/D vssd1 vssd1 vccd1 vccd1 _25607_/Q sky130_fd_sc_hd__dfxtp_4
X_22819_ _22875_/A vssd1 vssd1 vccd1 vccd1 _22888_/S sky130_fd_sc_hd__buf_8
X_26587_ _27058_/CLK _26587_/D vssd1 vssd1 vccd1 vccd1 _26587_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23799_ _23699_/X _26784_/Q _23799_/S vssd1 vssd1 vccd1 vccd1 _23800_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16340_ _26545_/Q _26153_/Q _16341_/S vssd1 vssd1 vccd1 vccd1 _16340_/X sky130_fd_sc_hd__mux2_1
X_25538_ _26974_/CLK _25538_/D vssd1 vssd1 vccd1 vccd1 _25538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13552_ _13552_/A _17821_/B vssd1 vssd1 vccd1 vccd1 _13553_/B sky130_fd_sc_hd__nor2_1
XFILLER_12_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13483_ _13941_/A vssd1 vssd1 vccd1 vccd1 _13484_/A sky130_fd_sc_hd__buf_2
X_16271_ _26119_/Q _26020_/Q _16271_/S vssd1 vssd1 vccd1 vccd1 _16271_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25469_ _25598_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 _25469_/Q sky130_fd_sc_hd__dfxtp_1
X_18010_ _18339_/A _18785_/A _18010_/C _18010_/D vssd1 vssd1 vccd1 vccd1 _18010_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27208_ _27230_/CLK _27208_/D vssd1 vssd1 vccd1 vccd1 _27208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15222_ _26932_/Q _16354_/S vssd1 vssd1 vccd1 vccd1 _15222_/X sky130_fd_sc_hd__or2_1
XFILLER_172_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27139_ _27164_/CLK _27139_/D vssd1 vssd1 vccd1 vccd1 _27139_/Q sky130_fd_sc_hd__dfxtp_2
X_15153_ _15634_/S vssd1 vssd1 vccd1 vccd1 _16161_/S sky130_fd_sc_hd__buf_2
XFILLER_10_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14104_ _25874_/Q _14109_/B vssd1 vssd1 vccd1 vccd1 _14104_/X sky130_fd_sc_hd__or2_1
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15084_ _25895_/Q _16419_/B vssd1 vssd1 vccd1 vccd1 _15084_/X sky130_fd_sc_hd__or2_1
X_19961_ _19956_/X _19957_/Y _19959_/Y _19787_/A vssd1 vssd1 vccd1 vccd1 _19961_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_154_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14035_ _14323_/B _14834_/C _12869_/X vssd1 vssd1 vccd1 vccd1 _14035_/X sky130_fd_sc_hd__a21o_1
X_18912_ _18912_/A _18912_/B vssd1 vssd1 vccd1 vccd1 _18912_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19892_ _19763_/X _19878_/X _19891_/Y _20067_/A vssd1 vssd1 vccd1 vccd1 _19892_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_268_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18843_ _25737_/Q _25736_/Q _19946_/A _18843_/D vssd1 vssd1 vccd1 vccd1 _18892_/C
+ sky130_fd_sc_hd__and4_2
XFILLER_95_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18774_ _18741_/X _18772_/X _18773_/X vssd1 vssd1 vccd1 vccd1 _18774_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_110_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15986_ _12769_/A _26888_/Q _26760_/Q _14004_/S vssd1 vssd1 vccd1 vccd1 _15986_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_95_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17725_ _18161_/B _17750_/A _18172_/A _17725_/D vssd1 vssd1 vccd1 vccd1 _17732_/B
+ sky130_fd_sc_hd__and4b_4
XFILLER_208_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14937_ _16409_/B _15954_/C vssd1 vssd1 vccd1 vccd1 _14937_/Y sky130_fd_sc_hd__nor2_1
XFILLER_282_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17656_ _21709_/A _17656_/B vssd1 vssd1 vccd1 vccd1 _25596_/D sky130_fd_sc_hd__nor2_1
X_14868_ _26549_/Q _26157_/Q _14876_/S vssd1 vssd1 vccd1 vccd1 _14868_/X sky130_fd_sc_hd__mux2_1
XFILLER_251_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16607_ _19156_/A vssd1 vssd1 vccd1 vccd1 _19155_/A sky130_fd_sc_hd__inv_2
X_13819_ _26659_/Q _25699_/Q _15768_/S vssd1 vssd1 vccd1 vccd1 _13819_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17587_ _17595_/A _17587_/B vssd1 vssd1 vccd1 vccd1 _25578_/D sky130_fd_sc_hd__nor2_1
XFILLER_223_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14799_ _14747_/A _25788_/Q _14813_/S _26874_/Q _14733_/A vssd1 vssd1 vccd1 vccd1
+ _14799_/X sky130_fd_sc_hd__o221a_1
XFILLER_211_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19326_ _19325_/Y _19292_/B _17787_/Y vssd1 vssd1 vccd1 vccd1 _19327_/B sky130_fd_sc_hd__a21bo_1
XFILLER_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16538_ _26095_/Q _25900_/Q _16541_/S vssd1 vssd1 vccd1 vccd1 _16538_/X sky130_fd_sc_hd__mux2_1
X_19257_ _17317_/X _18439_/X _18441_/X _25558_/Q vssd1 vssd1 vccd1 vccd1 _19257_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16469_ _26683_/Q _25723_/Q _16500_/S vssd1 vssd1 vccd1 vccd1 _16469_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18208_ _17911_/X _17900_/X _18209_/S vssd1 vssd1 vccd1 vccd1 _18208_/X sky130_fd_sc_hd__mux2_1
X_19188_ _19155_/A _19155_/B _17793_/X vssd1 vssd1 vccd1 vccd1 _19189_/B sky130_fd_sc_hd__a21bo_1
XFILLER_157_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18139_ _18381_/A vssd1 vssd1 vccd1 vccd1 _18705_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21150_ _25922_/Q _21148_/X _21149_/X input22/X vssd1 vssd1 vccd1 vccd1 _21151_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_176_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20101_ _19833_/X _20151_/C _20099_/Y _20100_/X vssd1 vssd1 vccd1 vccd1 _20102_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_104_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21081_ _25903_/Q _21074_/X _21077_/X input21/X vssd1 vssd1 vccd1 vccd1 _21082_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20032_ _17995_/A _19914_/A _20189_/B _20089_/A vssd1 vssd1 vccd1 vccd1 _20061_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24840_ _24877_/A vssd1 vssd1 vccd1 vccd1 _24856_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_39_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21983_ _26105_/Q _20900_/X _21983_/S vssd1 vssd1 vccd1 vccd1 _21984_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24771_ _24771_/A vssd1 vssd1 vccd1 vccd1 _24771_/X sky130_fd_sc_hd__buf_2
XFILLER_96_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26510_ _27285_/CLK _26510_/D vssd1 vssd1 vccd1 vccd1 _26510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23722_ _23722_/A vssd1 vssd1 vccd1 vccd1 _23722_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20934_ _20934_/A vssd1 vssd1 vccd1 vccd1 _25848_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26441_ _27280_/CLK _26441_/D vssd1 vssd1 vccd1 vccd1 _26441_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23653_ _23653_/A vssd1 vssd1 vccd1 vccd1 _26733_/D sky130_fd_sc_hd__clkbuf_1
X_20865_ _20865_/A vssd1 vssd1 vccd1 vccd1 _25828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22604_ _26317_/Q _22604_/B vssd1 vssd1 vccd1 vccd1 _22604_/Y sky130_fd_sc_hd__nand2_1
XFILLER_224_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26372_ _26468_/CLK _26372_/D vssd1 vssd1 vccd1 vccd1 _26372_/Q sky130_fd_sc_hd__dfxtp_1
X_23584_ _23584_/A vssd1 vssd1 vccd1 vccd1 _23584_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_241_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20796_ _21718_/A _20796_/B _20796_/C vssd1 vssd1 vccd1 vccd1 _20797_/A sky130_fd_sc_hd__and3_1
XFILLER_195_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25323_ _25391_/S vssd1 vssd1 vccd1 vccd1 _25332_/S sky130_fd_sc_hd__buf_2
X_22535_ _22535_/A _22535_/B vssd1 vssd1 vccd1 vccd1 _26292_/D sky130_fd_sc_hd__nor2_1
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22466_ _26210_/Q _22459_/X _22465_/X _22455_/X vssd1 vssd1 vccd1 vccd1 _26258_/D
+ sky130_fd_sc_hd__o211a_1
X_25254_ _23690_/X _27232_/Q _25260_/S vssd1 vssd1 vccd1 vccd1 _25255_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24205_ _26959_/Q _24205_/B vssd1 vssd1 vccd1 vccd1 _24213_/C sky130_fd_sc_hd__and2_1
X_21417_ _21364_/X _18834_/X _21365_/X _25810_/Q _21403_/X vssd1 vssd1 vccd1 vccd1
+ _21417_/X sky130_fd_sc_hd__a221o_1
X_25185_ _24915_/A _25218_/B _25184_/Y vssd1 vssd1 vccd1 vccd1 _27202_/D sky130_fd_sc_hd__a21oi_1
X_22397_ _22379_/X _22340_/S _22380_/X _22396_/Y vssd1 vssd1 vccd1 vccd1 _26237_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24136_ _26934_/Q _23594_/X _24142_/S vssd1 vssd1 vccd1 vccd1 _24137_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21348_ _21345_/X _21347_/X _21290_/A vssd1 vssd1 vccd1 vccd1 _21348_/X sky130_fd_sc_hd__a21o_1
XFILLER_2_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24067_ _24067_/A vssd1 vssd1 vccd1 vccd1 _26903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21279_ _21279_/A vssd1 vssd1 vccd1 vccd1 _21279_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23018_ _23018_/A vssd1 vssd1 vccd1 vccd1 _26480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15840_ _16183_/S _15838_/X _15839_/X _13274_/A vssd1 vssd1 vccd1 vccd1 _15840_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _15109_/A _25844_/Q _26044_/Q _13492_/X _13363_/A vssd1 vssd1 vccd1 vccd1
+ _15771_/X sky130_fd_sc_hd__a221o_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24969_ _24969_/A _24972_/B vssd1 vssd1 vccd1 vccd1 _24969_/Y sky130_fd_sc_hd__nand2_1
X_12983_ _20868_/A vssd1 vssd1 vccd1 vccd1 _20488_/A sky130_fd_sc_hd__clkinv_2
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17510_ _19603_/A _18088_/A vssd1 vssd1 vccd1 vccd1 _19594_/A sky130_fd_sc_hd__nor2_1
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26708_ _26900_/CLK _26708_/D vssd1 vssd1 vccd1 vccd1 _26708_/Q sky130_fd_sc_hd__dfxtp_1
X_14722_ _14722_/A vssd1 vssd1 vccd1 vccd1 _14723_/A sky130_fd_sc_hd__buf_4
XFILLER_217_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18490_ _18345_/S _18490_/B vssd1 vssd1 vccd1 vccd1 _18490_/X sky130_fd_sc_hd__and2b_1
XFILLER_91_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _25564_/Q _17438_/B _17440_/Y vssd1 vssd1 vccd1 vccd1 _25564_/D sky130_fd_sc_hd__o21a_1
XFILLER_232_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_178_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26683_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14653_ _15635_/B vssd1 vssd1 vccd1 vccd1 _16310_/B sky130_fd_sc_hd__clkbuf_4
X_26639_ _26799_/CLK _26639_/D vssd1 vssd1 vccd1 vccd1 _26639_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_107_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26307_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13604_ _25806_/Q _13043_/A _14254_/S _13603_/X vssd1 vssd1 vccd1 vccd1 _13604_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17372_ _25543_/Q _17372_/B vssd1 vssd1 vccd1 vccd1 _17379_/C sky130_fd_sc_hd__and2_1
XFILLER_159_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14584_ _16368_/S vssd1 vssd1 vccd1 vccd1 _16451_/S sky130_fd_sc_hd__buf_2
XFILLER_158_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19111_ _19235_/B _19576_/C vssd1 vssd1 vccd1 vccd1 _19111_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16323_ _25854_/Q _26054_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _16323_/X sky130_fd_sc_hd__mux2_1
X_13535_ _27273_/Q _26466_/Q _13535_/S vssd1 vssd1 vccd1 vccd1 _13535_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19042_ _19042_/A _19042_/B vssd1 vssd1 vccd1 vccd1 _19042_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16254_ _15085_/A _16252_/X _16253_/X _15318_/X vssd1 vssd1 vccd1 vccd1 _16254_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_71_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13466_ _13466_/A vssd1 vssd1 vccd1 vccd1 _13466_/X sky130_fd_sc_hd__buf_6
XFILLER_9_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15205_ _15205_/A vssd1 vssd1 vccd1 vccd1 _16183_/S sky130_fd_sc_hd__buf_6
XFILLER_154_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16185_ _16185_/A _16185_/B vssd1 vssd1 vccd1 vccd1 _16185_/X sky130_fd_sc_hd__or2_1
X_13397_ _14407_/A _13397_/B _13559_/B _13397_/D vssd1 vssd1 vccd1 vccd1 _13397_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_5_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15136_ _25654_/Q _14609_/A _15135_/X vssd1 vssd1 vccd1 vccd1 _15136_/X sky130_fd_sc_hd__a21o_1
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15067_ _12750_/A _15062_/X _15066_/X vssd1 vssd1 vccd1 vccd1 _15068_/B sky130_fd_sc_hd__o21ai_1
X_19944_ _25572_/Q _19600_/X _19968_/A _19589_/A vssd1 vssd1 vccd1 vccd1 _19944_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14018_ _13009_/A _23530_/A _14017_/X _13027_/A vssd1 vssd1 vccd1 vccd1 _16830_/B
+ sky130_fd_sc_hd__o211a_4
X_19875_ _22487_/A _19721_/X _19863_/X _19871_/X _19874_/X vssd1 vssd1 vccd1 vccd1
+ _25668_/D sky130_fd_sc_hd__o221a_1
XFILLER_96_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18826_ _18826_/A vssd1 vssd1 vccd1 vccd1 _18826_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18757_ _18757_/A vssd1 vssd1 vccd1 vccd1 _19465_/B sky130_fd_sc_hd__clkbuf_1
X_15969_ _26500_/Q _26372_/Q _15988_/S vssd1 vssd1 vccd1 vccd1 _15969_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17708_ _17708_/A _17708_/B vssd1 vssd1 vccd1 vccd1 _17708_/X sky130_fd_sc_hd__or2_1
XFILLER_247_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18688_ _18682_/X _17988_/X _18683_/X _18687_/X vssd1 vssd1 vccd1 vccd1 _18688_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_251_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17639_ _17534_/X _17627_/X _12898_/X _17536_/X _25929_/Q vssd1 vssd1 vccd1 vccd1
+ _17639_/Y sky130_fd_sc_hd__o32ai_1
XFILLER_24_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20650_ _20650_/A _20656_/B vssd1 vssd1 vccd1 vccd1 _20650_/X sky130_fd_sc_hd__or2_1
XFILLER_210_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19309_ _19309_/A _19442_/B vssd1 vssd1 vccd1 vccd1 _19309_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20581_ _20580_/X _25713_/Q _20593_/S vssd1 vssd1 vccd1 vccd1 _20582_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22320_ _26218_/Q _22315_/X _22318_/X _22319_/X vssd1 vssd1 vccd1 vccd1 _26218_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_220_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_opt_10_0_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_48_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22251_ _26196_/Q _22235_/X _22250_/X _22243_/X vssd1 vssd1 vccd1 vccd1 _26196_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21202_ _21202_/A vssd1 vssd1 vccd1 vccd1 _21202_/X sky130_fd_sc_hd__buf_2
XFILLER_191_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22182_ _26178_/Q _22169_/X _22180_/X _22181_/X vssd1 vssd1 vccd1 vccd1 _26178_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_254_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21133_ _21136_/A _21133_/B vssd1 vssd1 vccd1 vccd1 _21134_/A sky130_fd_sc_hd__or2_1
X_26990_ _26992_/CLK _26990_/D vssd1 vssd1 vccd1 vccd1 _26990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25941_ _27058_/CLK _25941_/D vssd1 vssd1 vccd1 vccd1 _25941_/Q sky130_fd_sc_hd__dfxtp_1
X_21064_ _21064_/A vssd1 vssd1 vccd1 vccd1 _25900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20015_ _20015_/A vssd1 vssd1 vccd1 vccd1 _20015_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25872_ _26592_/CLK _25872_/D vssd1 vssd1 vccd1 vccd1 _25872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24823_ _20650_/A _24810_/X _24686_/Y _24811_/X vssd1 vssd1 vccd1 vccd1 _24823_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_104_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_5_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27285_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_261_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24754_ _24974_/A vssd1 vssd1 vccd1 vccd1 _24755_/B sky130_fd_sc_hd__inv_2
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21966_ _26097_/Q _20875_/X _21972_/S vssd1 vssd1 vccd1 vccd1 _21967_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23705_ _23705_/A vssd1 vssd1 vccd1 vccd1 _26753_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20917_ _25843_/Q _20916_/X _20917_/S vssd1 vssd1 vccd1 vccd1 _20918_/A sky130_fd_sc_hd__mux2_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21897_ _21897_/A vssd1 vssd1 vccd1 vccd1 _26066_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24685_ _24706_/A vssd1 vssd1 vccd1 vccd1 _24703_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_230_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_200_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27329_/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26424_ _27264_/CLK _26424_/D vssd1 vssd1 vccd1 vccd1 _26424_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_199_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23636_ _23682_/S vssd1 vssd1 vccd1 vccd1 _23645_/S sky130_fd_sc_hd__buf_6
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20848_ _25820_/Q vssd1 vssd1 vccd1 vccd1 _20849_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_42_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26355_ _26483_/CLK _26355_/D vssd1 vssd1 vccd1 vccd1 _26355_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_196_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23567_ _23567_/A vssd1 vssd1 vccd1 vccd1 _26701_/D sky130_fd_sc_hd__clkbuf_1
X_20779_ _20605_/X _25785_/Q _20783_/S vssd1 vssd1 vccd1 vccd1 _20780_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13320_ _26531_/Q _26139_/Q _15671_/S vssd1 vssd1 vccd1 vccd1 _13321_/B sky130_fd_sc_hd__mux2_1
X_25306_ _25306_/A vssd1 vssd1 vccd1 vccd1 _25315_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_183_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22518_ _22518_/A _22524_/B vssd1 vssd1 vccd1 vccd1 _22519_/A sky130_fd_sc_hd__and2_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23498_ _26679_/Q _23124_/X _23502_/S vssd1 vssd1 vccd1 vccd1 _23499_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26286_ _26286_/CLK _26286_/D vssd1 vssd1 vccd1 vccd1 _26286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13251_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13252_/A sky130_fd_sc_hd__clkbuf_4
X_22449_ _26203_/Q _22446_/X _22448_/X _22442_/X vssd1 vssd1 vccd1 vccd1 _26251_/D
+ sky130_fd_sc_hd__o211a_1
X_25237_ _24988_/X _19614_/D _24771_/X _24755_/B _25219_/X vssd1 vssd1 vccd1 vccd1
+ _25237_/X sky130_fd_sc_hd__a221o_1
XFILLER_109_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13182_ _15659_/A _14833_/A vssd1 vssd1 vccd1 vccd1 _16508_/S sky130_fd_sc_hd__nor2_1
X_25168_ _25755_/Q _25138_/A _25167_/X vssd1 vssd1 vccd1 vccd1 _25168_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_191_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24119_ _24119_/A vssd1 vssd1 vccd1 vccd1 _26926_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ _17990_/A vssd1 vssd1 vccd1 vccd1 _18602_/A sky130_fd_sc_hd__clkbuf_2
X_25099_ _20668_/A _25086_/X _25098_/X vssd1 vssd1 vccd1 vccd1 _25099_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_269_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16941_ _16957_/A _16889_/X _16938_/X _16840_/A _16940_/Y vssd1 vssd1 vccd1 vccd1
+ _16942_/B sky130_fd_sc_hd__o221a_1
XFILLER_265_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19660_ _19607_/A _19607_/B _19659_/Y vssd1 vssd1 vccd1 vccd1 _19675_/A sky130_fd_sc_hd__a21oi_2
X_16872_ _16463_/X _23552_/A _15910_/X _16860_/B vssd1 vssd1 vccd1 vccd1 _16872_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_277_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18611_ _27078_/Q vssd1 vssd1 vccd1 vccd1 _19957_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_237_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15823_ _12745_/A _15822_/X _15720_/S vssd1 vssd1 vccd1 vccd1 _15823_/X sky130_fd_sc_hd__a21o_1
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19591_ _25757_/Q _25756_/Q vssd1 vssd1 vccd1 vccd1 _19633_/C sky130_fd_sc_hd__or2_1
XFILLER_265_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ _19235_/B _19572_/C _18541_/X _18037_/X vssd1 vssd1 vccd1 vccd1 _18542_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_246_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15754_ _13330_/A _15751_/X _15753_/X _13340_/A vssd1 vssd1 vccd1 vccd1 _15754_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12966_ _13803_/B vssd1 vssd1 vccd1 vccd1 _15532_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_90 _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14705_ _15187_/A vssd1 vssd1 vccd1 vccd1 _14706_/A sky130_fd_sc_hd__buf_2
XFILLER_261_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18473_ _18435_/X _18471_/X _18474_/B vssd1 vssd1 vccd1 vccd1 _18473_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15685_ _15406_/A _26112_/Q _26013_/Q _15674_/X _15672_/A vssd1 vssd1 vccd1 vccd1
+ _15685_/X sky130_fd_sc_hd__a221o_1
X_12897_ _14402_/S vssd1 vssd1 vccd1 vccd1 _14488_/S sky130_fd_sc_hd__buf_4
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17424_ _17427_/A _17427_/C _17414_/X vssd1 vssd1 vccd1 vccd1 _17424_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14636_ _14953_/S vssd1 vssd1 vccd1 vccd1 _14692_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _25537_/Q _17353_/B _17354_/Y vssd1 vssd1 vccd1 vccd1 _25537_/D sky130_fd_sc_hd__o21a_1
XFILLER_220_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14567_ _14567_/A vssd1 vssd1 vccd1 vccd1 _17805_/B sky130_fd_sc_hd__inv_2
XFILLER_159_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16306_ _26353_/Q _26613_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _16306_/X sky130_fd_sc_hd__mux2_1
X_13518_ _25807_/Q _27241_/Q _15857_/S vssd1 vssd1 vccd1 vccd1 _13518_/X sky130_fd_sc_hd__mux2_1
X_17286_ _25516_/Q _17284_/B _17285_/Y vssd1 vssd1 vccd1 vccd1 _25516_/D sky130_fd_sc_hd__o21a_1
X_14498_ _13890_/X _25758_/Q _15726_/S _26844_/Q _13124_/A vssd1 vssd1 vccd1 vccd1
+ _14498_/X sky130_fd_sc_hd__o221a_1
XFILLER_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19025_ _27023_/Q _18449_/X _19024_/X _18821_/X vssd1 vssd1 vccd1 vccd1 _19025_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16237_ _25820_/Q _15014_/S _16241_/S _16236_/X vssd1 vssd1 vccd1 vccd1 _16237_/X
+ sky130_fd_sc_hd__o211a_1
X_13449_ _12770_/A _26694_/Q _26822_/Q _15459_/S _13050_/A vssd1 vssd1 vccd1 vccd1
+ _13449_/X sky130_fd_sc_hd__a221o_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_75_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27265_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_161_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16168_ _16150_/X _16167_/X _14591_/A vssd1 vssd1 vccd1 vccd1 _16168_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_114_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15119_ _26122_/Q _26023_/Q _15119_/S vssd1 vssd1 vccd1 vccd1 _15119_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16099_ _15676_/X _27282_/Q _26475_/Q _16273_/S _13532_/X vssd1 vssd1 vccd1 vccd1
+ _16099_/X sky130_fd_sc_hd__a221o_1
XFILLER_173_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19927_ _19766_/A _19925_/Y _19926_/X vssd1 vssd1 vccd1 vccd1 _19927_/X sky130_fd_sc_hd__a21o_1
XFILLER_205_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19858_ _19980_/A _19981_/A vssd1 vssd1 vccd1 vccd1 _19860_/A sky130_fd_sc_hd__and2_1
XFILLER_217_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18809_ _17278_/X _18807_/X _18808_/X _25546_/Q vssd1 vssd1 vccd1 vccd1 _18809_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19789_ _19784_/Y _19785_/Y _19788_/Y vssd1 vssd1 vccd1 vccd1 _19789_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21820_ _21820_/A vssd1 vssd1 vccd1 vccd1 _26039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21751_ _21751_/A vssd1 vssd1 vccd1 vccd1 _26009_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20702_ _26291_/Q _20687_/B _20701_/Y _20697_/X vssd1 vssd1 vccd1 vccd1 _25754_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21682_ _21682_/A vssd1 vssd1 vccd1 vccd1 _25980_/D sky130_fd_sc_hd__clkbuf_1
X_24470_ _24551_/A vssd1 vssd1 vccd1 vccd1 _24470_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_260_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20633_ _20646_/A vssd1 vssd1 vccd1 vccd1 _20633_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_23421_ _23421_/A vssd1 vssd1 vccd1 vccd1 _23430_/S sky130_fd_sc_hd__buf_6
XFILLER_221_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26140_ _26468_/CLK _26140_/D vssd1 vssd1 vccd1 vccd1 _26140_/Q sky130_fd_sc_hd__dfxtp_1
X_23352_ _23352_/A vssd1 vssd1 vccd1 vccd1 _26614_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20564_ _20563_/X _25709_/Q _20572_/S vssd1 vssd1 vccd1 vccd1 _20565_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22303_ _24441_/A vssd1 vssd1 vccd1 vccd1 _22428_/A sky130_fd_sc_hd__clkbuf_4
X_26071_ _26594_/CLK _26071_/D vssd1 vssd1 vccd1 vccd1 _26071_/Q sky130_fd_sc_hd__dfxtp_1
X_23283_ _26584_/Q input247/X _23289_/S vssd1 vssd1 vccd1 vccd1 _23284_/A sky130_fd_sc_hd__mux2_1
X_20495_ _23514_/A vssd1 vssd1 vccd1 vccd1 _23690_/A sky130_fd_sc_hd__buf_2
XFILLER_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22234_ _22315_/A vssd1 vssd1 vccd1 vccd1 _22269_/A sky130_fd_sc_hd__buf_2
X_25022_ _24654_/A _25014_/X _25021_/Y _24773_/X vssd1 vssd1 vccd1 vccd1 _25022_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_279_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22165_ _26173_/Q _22152_/X _22163_/X _22164_/X vssd1 vssd1 vccd1 vccd1 _26173_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_279_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21116_ _21116_/A vssd1 vssd1 vccd1 vccd1 _25912_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26973_ _26974_/CLK _26973_/D vssd1 vssd1 vccd1 vccd1 _26973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22096_ _22096_/A vssd1 vssd1 vccd1 vccd1 _26155_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21047_ _21047_/A vssd1 vssd1 vccd1 vccd1 _25892_/D sky130_fd_sc_hd__clkbuf_1
X_25924_ _27213_/CLK _25924_/D vssd1 vssd1 vccd1 vccd1 _25924_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_8_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25855_ _26483_/CLK _25855_/D vssd1 vssd1 vccd1 vccd1 _25855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12820_ _25472_/Q vssd1 vssd1 vccd1 vccd1 _21300_/A sky130_fd_sc_hd__clkbuf_2
X_24806_ _27107_/Q _24818_/B vssd1 vssd1 vccd1 vccd1 _24806_/Y sky130_fd_sc_hd__nand2_1
XFILLER_228_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25786_ _26677_/CLK _25786_/D vssd1 vssd1 vccd1 vccd1 _25786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_264_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22998_ _26471_/Q _22691_/X _23006_/S vssd1 vssd1 vccd1 vccd1 _22999_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12751_ _12751_/A vssd1 vssd1 vccd1 vccd1 _12760_/B sky130_fd_sc_hd__buf_2
X_24737_ _27091_/Q _24724_/X _24736_/Y _24720_/X vssd1 vssd1 vccd1 vccd1 _24738_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_243_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21949_ _20601_/X _26090_/Q _21955_/S vssd1 vssd1 vccd1 vccd1 _21950_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15174_/A _15467_/X _15469_/X _13144_/A vssd1 vssd1 vccd1 vccd1 _15470_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _13215_/A _25567_/Q vssd1 vssd1 vccd1 vccd1 _17500_/B sky130_fd_sc_hd__and2_1
X_24668_ _24682_/A _24668_/B vssd1 vssd1 vccd1 vccd1 _24668_/Y sky130_fd_sc_hd__nand2_2
XFILLER_202_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14421_ _14421_/A _14421_/B _14421_/C vssd1 vssd1 vccd1 vccd1 _14421_/X sky130_fd_sc_hd__and3_1
X_26407_ _27281_/CLK _26407_/D vssd1 vssd1 vccd1 vccd1 _26407_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23619_ _26718_/Q _23517_/X _23623_/S vssd1 vssd1 vccd1 vccd1 _23620_/A sky130_fd_sc_hd__mux2_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24599_ _27055_/Q _24589_/X _24598_/Y _24593_/X vssd1 vssd1 vccd1 vccd1 _27055_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17140_ _18338_/A vssd1 vssd1 vccd1 vccd1 _17200_/A sky130_fd_sc_hd__clkbuf_2
X_26338_ _27277_/CLK _26338_/D vssd1 vssd1 vccd1 vccd1 _26338_/Q sky130_fd_sc_hd__dfxtp_2
X_14352_ _14350_/X _14351_/X _14352_/S vssd1 vssd1 vccd1 vccd1 _14352_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ _14077_/A vssd1 vssd1 vccd1 vccd1 _13304_/A sky130_fd_sc_hd__buf_4
X_17071_ _25979_/Q _17061_/A _17000_/X _17015_/X vssd1 vssd1 vccd1 vccd1 _17071_/X
+ sky130_fd_sc_hd__a22o_4
X_26269_ _26271_/CLK _26269_/D vssd1 vssd1 vccd1 vccd1 _26269_/Q sky130_fd_sc_hd__dfxtp_1
X_14283_ _14187_/A _16820_/B _14282_/Y vssd1 vssd1 vccd1 vccd1 _14283_/Y sky130_fd_sc_hd__a21oi_1
X_16022_ _16022_/A _16022_/B vssd1 vssd1 vccd1 vccd1 _16022_/X sky130_fd_sc_hd__or2_1
XFILLER_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13234_ _16111_/A vssd1 vssd1 vccd1 vccd1 _15424_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13165_ _14647_/A _13153_/X _13160_/X _14677_/A vssd1 vssd1 vccd1 vccd1 _13165_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13096_ _26531_/Q _26139_/Q _15467_/S vssd1 vssd1 vccd1 vccd1 _13096_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17973_ _17973_/A _18186_/A vssd1 vssd1 vccd1 vccd1 _18271_/B sky130_fd_sc_hd__nor2_2
XFILLER_78_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19712_ _19712_/A _19712_/B vssd1 vssd1 vccd1 vccd1 _19712_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16924_ _16924_/A _16924_/B vssd1 vssd1 vccd1 vccd1 _16925_/A sky130_fd_sc_hd__and2_1
XFILLER_278_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_193_wb_clk_i _26681_/CLK vssd1 vssd1 vccd1 vccd1 _27258_/CLK sky130_fd_sc_hd__clkbuf_16
X_19643_ _27134_/Q _27133_/Q _25218_/A vssd1 vssd1 vccd1 vccd1 _19646_/A sky130_fd_sc_hd__and3b_1
XFILLER_66_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16855_ _16855_/A _16855_/B vssd1 vssd1 vccd1 vccd1 _16855_/Y sky130_fd_sc_hd__nand2_1
XFILLER_226_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_122_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25547_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15806_ _15804_/X _15805_/X _15806_/S vssd1 vssd1 vccd1 vccd1 _15806_/X sky130_fd_sc_hd__mux2_1
XFILLER_265_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19574_ _19574_/A _19574_/B _19574_/C _18941_/Y vssd1 vssd1 vccd1 vccd1 _19574_/X
+ sky130_fd_sc_hd__or4b_1
X_16786_ _16784_/X _16785_/Y _16693_/X vssd1 vssd1 vccd1 vccd1 _16786_/X sky130_fd_sc_hd__a21o_1
XFILLER_207_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13998_ _13992_/X _13997_/X _13998_/S vssd1 vssd1 vccd1 vccd1 _13998_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18525_ _18577_/A vssd1 vssd1 vccd1 vccd1 _19268_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15737_ _13698_/A _15734_/X _15736_/X _13863_/X vssd1 vssd1 vccd1 vccd1 _15737_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12949_ _12944_/X _12945_/X _12948_/Y vssd1 vssd1 vccd1 vccd1 _14486_/B sky130_fd_sc_hd__a21o_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18456_ _18450_/X _18451_/X _18453_/X _18455_/X _18120_/D vssd1 vssd1 vccd1 vccd1
+ _18456_/X sky130_fd_sc_hd__a221o_1
XFILLER_61_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15668_ _15668_/A _15668_/B vssd1 vssd1 vccd1 vccd1 _15668_/Y sky130_fd_sc_hd__nor2_1
X_17407_ _17408_/A _17408_/C _25554_/Q vssd1 vssd1 vccd1 vccd1 _17409_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14619_ _25628_/Q _14597_/X _14615_/X _14618_/X vssd1 vssd1 vccd1 vccd1 _23606_/A
+ sky130_fd_sc_hd__o22a_4
X_18387_ _25506_/Q _18556_/A _18557_/A _17356_/X vssd1 vssd1 vccd1 vccd1 _18387_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15599_ _15676_/A _25846_/Q _26046_/Q _16194_/S _15576_/A vssd1 vssd1 vccd1 vccd1
+ _15599_/X sky130_fd_sc_hd__a221o_1
XFILLER_267_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17338_ _17336_/X _17341_/C _17337_/Y vssd1 vssd1 vccd1 vccd1 _25532_/D sky130_fd_sc_hd__o21a_1
XFILLER_159_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17269_ _17414_/A vssd1 vssd1 vccd1 vccd1 _17269_/X sky130_fd_sc_hd__buf_2
XFILLER_162_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19008_ _25615_/Q _18971_/X _19006_/X _19007_/X vssd1 vssd1 vccd1 vccd1 _25615_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20280_ _20280_/A _20280_/B vssd1 vssd1 vccd1 vccd1 _20280_/Y sky130_fd_sc_hd__nand2_1
XFILLER_283_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23970_ _26860_/Q _23562_/X _23976_/S vssd1 vssd1 vccd1 vccd1 _23971_/A sky130_fd_sc_hd__mux2_1
XFILLER_275_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22921_ _26437_/Q _22685_/X _22923_/S vssd1 vssd1 vccd1 vccd1 _22922_/A sky130_fd_sc_hd__mux2_1
XFILLER_272_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25640_ _25661_/CLK _25640_/D vssd1 vssd1 vccd1 vccd1 _25640_/Q sky130_fd_sc_hd__dfxtp_1
X_22852_ _22852_/A vssd1 vssd1 vccd1 vccd1 _26406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21803_ _26032_/Q _20881_/X _21805_/S vssd1 vssd1 vccd1 vccd1 _21804_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25571_ _26683_/CLK _25571_/D vssd1 vssd1 vccd1 vccd1 _25571_/Q sky130_fd_sc_hd__dfxtp_1
X_22783_ _26376_/Q _22695_/X _22789_/S vssd1 vssd1 vccd1 vccd1 _22784_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27310_ _27310_/CLK _27310_/D vssd1 vssd1 vccd1 vccd1 _27310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_5_0_wb_clk_i INSDIODE2_273/DIODE vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
X_24522_ _24538_/A _24978_/A vssd1 vssd1 vccd1 vccd1 _24522_/Y sky130_fd_sc_hd__nand2_1
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21734_ _21791_/S vssd1 vssd1 vccd1 vccd1 _21743_/S sky130_fd_sc_hd__clkbuf_4
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27241_ _27305_/CLK _27241_/D vssd1 vssd1 vccd1 vccd1 _27241_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24453_ _27020_/Q _24448_/X _24452_/Y _24442_/X vssd1 vssd1 vccd1 vccd1 _27020_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21665_ _23289_/S vssd1 vssd1 vccd1 vccd1 _21674_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23404_ _26637_/Q _23092_/X _23408_/S vssd1 vssd1 vccd1 vccd1 _23405_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20616_ _23606_/A vssd1 vssd1 vccd1 vccd1 _23782_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_27172_ _27176_/CLK _27172_/D vssd1 vssd1 vccd1 vccd1 _27172_/Q sky130_fd_sc_hd__dfxtp_1
X_24384_ _24501_/A vssd1 vssd1 vccd1 vccd1 _24384_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_21596_ _21592_/Y _21595_/X _21556_/X vssd1 vssd1 vccd1 vccd1 _21596_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_20_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26123_ _26900_/CLK _26123_/D vssd1 vssd1 vccd1 vccd1 _26123_/Q sky130_fd_sc_hd__dfxtp_1
X_20547_ _20546_/X _25705_/Q _20551_/S vssd1 vssd1 vccd1 vccd1 _20548_/A sky130_fd_sc_hd__mux2_1
X_23335_ _20571_/X _26607_/Q _23335_/S vssd1 vssd1 vccd1 vccd1 _23336_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26054_ _27288_/CLK _26054_/D vssd1 vssd1 vccd1 vccd1 _26054_/Q sky130_fd_sc_hd__dfxtp_1
X_23266_ _26576_/Q _23114_/X _23266_/S vssd1 vssd1 vccd1 vccd1 _23267_/A sky130_fd_sc_hd__mux2_1
X_20478_ _20478_/A _20478_/B vssd1 vssd1 vccd1 vccd1 _20478_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25005_ _25106_/A vssd1 vssd1 vccd1 vccd1 _25005_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22217_ _22288_/A vssd1 vssd1 vccd1 vccd1 _22217_/X sky130_fd_sc_hd__clkbuf_2
X_23197_ _26545_/Q _23117_/X _23205_/S vssd1 vssd1 vccd1 vccd1 _23198_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22148_ _22195_/A vssd1 vssd1 vccd1 vccd1 _22148_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_267_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput390 _17038_/X vssd1 vssd1 vccd1 vccd1 din0[22] sky130_fd_sc_hd__buf_2
XFILLER_126_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26956_ _26992_/CLK _26956_/D vssd1 vssd1 vccd1 vccd1 _26956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_266_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14970_ _27291_/Q _26484_/Q _14970_/S vssd1 vssd1 vccd1 vccd1 _14970_/X sky130_fd_sc_hd__mux2_1
X_22079_ _22090_/A vssd1 vssd1 vccd1 vccd1 _22088_/S sky130_fd_sc_hd__buf_4
XFILLER_282_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13921_ _17623_/B _13921_/B vssd1 vssd1 vccd1 vccd1 _13921_/Y sky130_fd_sc_hd__nor2_1
X_25907_ _27122_/CLK _25907_/D vssd1 vssd1 vccd1 vccd1 _25907_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_281_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26887_ _27312_/CLK _26887_/D vssd1 vssd1 vccd1 vccd1 _26887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_267_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16640_ _25934_/Q _25935_/Q vssd1 vssd1 vccd1 vccd1 _21075_/B sky130_fd_sc_hd__or2b_2
X_25838_ _26595_/CLK _25838_/D vssd1 vssd1 vccd1 vccd1 _25838_/Q sky130_fd_sc_hd__dfxtp_2
X_13852_ _25731_/Q _14317_/B vssd1 vssd1 vccd1 vccd1 _13852_/X sky130_fd_sc_hd__or2_1
XFILLER_75_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_407 _17045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12803_ _25571_/Q _25570_/Q _17504_/B _13269_/A vssd1 vssd1 vccd1 vccd1 _12803_/X
+ sky130_fd_sc_hd__o31a_2
X_16571_ _16571_/A _19277_/A vssd1 vssd1 vccd1 vccd1 _16776_/A sky130_fd_sc_hd__xnor2_1
XFILLER_262_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25769_ _27305_/CLK _25769_/D vssd1 vssd1 vccd1 vccd1 _25769_/Q sky130_fd_sc_hd__dfxtp_4
X_13783_ _15915_/S vssd1 vssd1 vccd1 vccd1 _15914_/S sky130_fd_sc_hd__buf_6
XINSDIODE2_418 _17014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_429 _12781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18310_ _18317_/S vssd1 vssd1 vccd1 vccd1 _18858_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_231_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15522_ _15510_/X _15513_/X _15521_/Y vssd1 vssd1 vccd1 vccd1 _15522_/Y sky130_fd_sc_hd__o21bai_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ _13249_/A vssd1 vssd1 vccd1 vccd1 _14453_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19290_ _19290_/A vssd1 vssd1 vccd1 vccd1 _19423_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _27008_/Q _19063_/A _18239_/X _18565_/A vssd1 vssd1 vccd1 vccd1 _18241_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15453_ _15453_/A vssd1 vssd1 vccd1 vccd1 _16069_/S sky130_fd_sc_hd__buf_4
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14404_ _14404_/A _14404_/B vssd1 vssd1 vccd1 vccd1 _14404_/Y sky130_fd_sc_hd__nand2_1
X_18172_ _18172_/A vssd1 vssd1 vccd1 vccd1 _18829_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_187_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15384_ _15382_/X _15383_/X _15384_/S vssd1 vssd1 vccd1 vccd1 _15384_/X sky130_fd_sc_hd__mux2_1
X_17123_ _17500_/B _20689_/A vssd1 vssd1 vccd1 vccd1 _17123_/X sky130_fd_sc_hd__or2_1
X_14335_ _13083_/A _26590_/Q _14269_/S _26330_/Q _13022_/A vssd1 vssd1 vccd1 vccd1
+ _14335_/X sky130_fd_sc_hd__o221a_1
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17054_ _26585_/Q _17003_/X _20792_/C _17051_/X vssd1 vssd1 vccd1 vccd1 _17054_/X
+ sky130_fd_sc_hd__a22o_4
X_14266_ _13890_/A _26687_/Q _26815_/Q _14497_/A _13048_/A vssd1 vssd1 vccd1 vccd1
+ _14266_/X sky130_fd_sc_hd__a221o_1
XFILLER_109_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16005_ _26500_/Q _26372_/Q _16005_/S vssd1 vssd1 vccd1 vccd1 _16006_/B sky130_fd_sc_hd__mux2_1
X_13217_ _13955_/A vssd1 vssd1 vccd1 vccd1 _13358_/A sky130_fd_sc_hd__clkbuf_4
X_14197_ _14369_/S vssd1 vssd1 vccd1 vccd1 _15858_/S sky130_fd_sc_hd__buf_4
XFILLER_140_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13148_ _14252_/S vssd1 vssd1 vccd1 vccd1 _14004_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_140_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13079_ _25703_/Q _15635_/B vssd1 vssd1 vccd1 vccd1 _13079_/X sky130_fd_sc_hd__or2_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17956_ _17842_/B _16035_/B _17956_/S vssd1 vssd1 vccd1 vccd1 _17956_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16907_ _16939_/A vssd1 vssd1 vccd1 vccd1 _16907_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17887_ _18058_/S vssd1 vssd1 vccd1 vccd1 _18063_/S sky130_fd_sc_hd__buf_2
XFILLER_239_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19626_ _27068_/Q _19616_/B input177/X _19623_/X _19625_/X vssd1 vssd1 vccd1 vccd1
+ _19626_/X sky130_fd_sc_hd__a311o_1
XFILLER_265_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16838_ _16838_/A _17772_/B vssd1 vssd1 vccd1 vccd1 _16859_/A sky130_fd_sc_hd__nor2_2
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19557_ _25656_/Q _19563_/B vssd1 vssd1 vccd1 vccd1 _19557_/X sky130_fd_sc_hd__or2_1
X_16769_ _16769_/A vssd1 vssd1 vccd1 vccd1 _16769_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18508_ _18508_/A vssd1 vssd1 vccd1 vccd1 _18508_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_222_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19488_ _20657_/A vssd1 vssd1 vccd1 vccd1 _19541_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_179_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18439_ _18439_/A vssd1 vssd1 vccd1 vccd1 _18439_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_178_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_90_wb_clk_i _25501_/CLK vssd1 vssd1 vccd1 vccd1 _25661_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21450_ _21450_/A vssd1 vssd1 vccd1 vccd1 _21450_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20401_ _20352_/A _20352_/B _20398_/Y _20400_/Y vssd1 vssd1 vccd1 vccd1 _20443_/B
+ sky130_fd_sc_hd__o31ai_2
XFILLER_174_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21381_ _21379_/X _21380_/X _21367_/X vssd1 vssd1 vccd1 vccd1 _21381_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20332_ _20332_/A _20351_/B vssd1 vssd1 vccd1 vccd1 _20332_/Y sky130_fd_sc_hd__xnor2_1
X_23120_ _23120_/A vssd1 vssd1 vccd1 vccd1 _26513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23051_ _26492_/Q _23050_/X _23051_/S vssd1 vssd1 vccd1 vccd1 _23052_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20263_ _25682_/Q _20286_/C vssd1 vssd1 vccd1 vccd1 _20265_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22002_ _22002_/A vssd1 vssd1 vccd1 vccd1 _26113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20194_ _20194_/A _20194_/B vssd1 vssd1 vccd1 vccd1 _20194_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput107 dout1[0] vssd1 vssd1 vccd1 vccd1 input107/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26810_ _27293_/CLK _26810_/D vssd1 vssd1 vccd1 vccd1 _26810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput118 dout1[1] vssd1 vssd1 vccd1 vccd1 input118/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput129 dout1[2] vssd1 vssd1 vccd1 vccd1 input129/X sky130_fd_sc_hd__clkbuf_1
XFILLER_276_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26741_ _26929_/CLK _26741_/D vssd1 vssd1 vccd1 vccd1 _26741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23953_ _23953_/A vssd1 vssd1 vccd1 vccd1 _26852_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22904_ _26429_/Q _22659_/X _22912_/S vssd1 vssd1 vccd1 vccd1 _22905_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26672_ _27283_/CLK _26672_/D vssd1 vssd1 vccd1 vccd1 _26672_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23884_ _23930_/S vssd1 vssd1 vccd1 vccd1 _23893_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25623_ _25624_/CLK _25623_/D vssd1 vssd1 vccd1 vccd1 _25623_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22835_ _22835_/A vssd1 vssd1 vccd1 vccd1 _26398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25554_ _25992_/CLK _25554_/D vssd1 vssd1 vccd1 vccd1 _25554_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22766_ _22766_/A vssd1 vssd1 vccd1 vccd1 _26368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24505_ _27029_/Q _24480_/X _24504_/Y _24499_/X vssd1 vssd1 vccd1 vccd1 _27029_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21717_ _20977_/A _21652_/X _16668_/B vssd1 vssd1 vccd1 vccd1 _21718_/C sky130_fd_sc_hd__o21ai_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25485_ _26683_/CLK _25485_/D vssd1 vssd1 vccd1 vccd1 _25485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22697_ _22697_/A vssd1 vssd1 vccd1 vccd1 _26344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27224_ _27228_/CLK _27224_/D vssd1 vssd1 vccd1 vccd1 _27224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24436_ _24494_/A vssd1 vssd1 vccd1 vccd1 _24464_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21648_ _21354_/A _25865_/Q _21647_/Y _21237_/X vssd1 vssd1 vccd1 vccd1 _21648_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_185_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27155_ _27227_/CLK _27155_/D vssd1 vssd1 vccd1 vccd1 _27155_/Q sky130_fd_sc_hd__dfxtp_2
X_24367_ _24645_/B vssd1 vssd1 vccd1 vccd1 _24550_/A sky130_fd_sc_hd__inv_2
XFILLER_181_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21579_ input60/X input95/X _21615_/S vssd1 vssd1 vccd1 vccd1 _21580_/A sky130_fd_sc_hd__mux2_8
X_26106_ _26601_/CLK _26106_/D vssd1 vssd1 vccd1 vccd1 _26106_/Q sky130_fd_sc_hd__dfxtp_2
X_14120_ _13141_/A _14115_/X _14119_/X _14354_/S vssd1 vssd1 vccd1 vccd1 _14120_/X
+ sky130_fd_sc_hd__o211a_1
X_23318_ _20538_/X _26599_/Q _23324_/S vssd1 vssd1 vccd1 vccd1 _23319_/A sky130_fd_sc_hd__mux2_1
X_27086_ _27087_/CLK _27086_/D vssd1 vssd1 vccd1 vccd1 _27086_/Q sky130_fd_sc_hd__dfxtp_1
X_24298_ _26990_/Q _24301_/C _24271_/X vssd1 vssd1 vccd1 vccd1 _24298_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_180_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26037_ _26601_/CLK _26037_/D vssd1 vssd1 vccd1 vccd1 _26037_/Q sky130_fd_sc_hd__dfxtp_4
X_14051_ _27300_/Q _26557_/Q _14544_/S vssd1 vssd1 vccd1 vccd1 _14051_/X sky130_fd_sc_hd__mux2_1
X_23249_ _26568_/Q _23089_/X _23255_/S vssd1 vssd1 vccd1 vccd1 _23250_/A sky130_fd_sc_hd__mux2_1
XFILLER_273_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13002_ _13002_/A vssd1 vssd1 vccd1 vccd1 _23363_/B sky130_fd_sc_hd__buf_2
XFILLER_279_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17810_ _17975_/A _17810_/B vssd1 vssd1 vccd1 vccd1 _18184_/C sky130_fd_sc_hd__nand2_1
X_18790_ _19352_/A vssd1 vssd1 vccd1 vccd1 _18790_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17741_ _18120_/C vssd1 vssd1 vccd1 vccd1 _18454_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14953_ _26648_/Q _26744_/Q _14953_/S vssd1 vssd1 vccd1 vccd1 _14953_/X sky130_fd_sc_hd__mux2_1
X_26939_ _26939_/CLK _26939_/D vssd1 vssd1 vccd1 vccd1 _26939_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13904_ _19828_/A _14124_/B vssd1 vssd1 vccd1 vccd1 _13904_/X sky130_fd_sc_hd__or2_1
X_17672_ _18138_/A _17971_/D vssd1 vssd1 vccd1 vccd1 _18554_/A sky130_fd_sc_hd__or2_1
XFILLER_263_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14884_ _14864_/X _14883_/X _14593_/A vssd1 vssd1 vccd1 vccd1 _14884_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_262_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16623_ _18978_/A vssd1 vssd1 vccd1 vccd1 _16624_/B sky130_fd_sc_hd__clkinv_2
X_19411_ _19196_/X _19409_/Y _19410_/X _19388_/A _19076_/X vssd1 vssd1 vccd1 vccd1
+ _19411_/X sky130_fd_sc_hd__o32a_1
X_13835_ _13835_/A vssd1 vssd1 vccd1 vccd1 _13835_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_204 _14559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_215 _19031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_226 _23549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_237 _19046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16554_ _25161_/A _25166_/A vssd1 vssd1 vccd1 vccd1 _17055_/A sky130_fd_sc_hd__nand2_1
X_19342_ _18554_/X _19340_/X _19341_/Y vssd1 vssd1 vccd1 vccd1 _19342_/Y sky130_fd_sc_hd__a21oi_1
X_13766_ _27303_/Q _26560_/Q _15768_/S vssd1 vssd1 vccd1 vccd1 _13766_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_248 _19256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_259 _20707_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15505_ _15499_/X _15504_/X _14816_/A vssd1 vssd1 vccd1 vccd1 _15505_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_189_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19273_ _19273_/A _19393_/B vssd1 vssd1 vccd1 vccd1 _19273_/Y sky130_fd_sc_hd__nand2_1
X_12717_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14956_/A sky130_fd_sc_hd__buf_2
XFILLER_149_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16485_ _17712_/B _26715_/Q _26843_/Q _16493_/S _17697_/B vssd1 vssd1 vccd1 vccd1
+ _16485_/X sky130_fd_sc_hd__a221o_1
X_13697_ _15645_/S _13693_/X _13696_/X _13031_/A vssd1 vssd1 vccd1 vccd1 _13697_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_176_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18224_ _14398_/X _18013_/X _18223_/Y _18022_/X _25600_/Q vssd1 vssd1 vccd1 vccd1
+ _18225_/B sky130_fd_sc_hd__a32o_1
X_15436_ _17790_/A _15438_/B vssd1 vssd1 vccd1 vccd1 _19105_/S sky130_fd_sc_hd__nand2_2
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18155_ _18438_/A vssd1 vssd1 vccd1 vccd1 _18807_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15367_ _26084_/Q _15351_/B _15031_/A _15366_/X vssd1 vssd1 vccd1 vccd1 _15367_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17106_ _18028_/A _17210_/A vssd1 vssd1 vccd1 vccd1 _17145_/A sky130_fd_sc_hd__nor2_1
X_14318_ _13180_/A _19700_/A _14317_/X vssd1 vssd1 vccd1 vccd1 _14567_/A sky130_fd_sc_hd__o21a_2
X_18086_ _18899_/A _18075_/Y _18085_/X _17503_/X vssd1 vssd1 vccd1 vccd1 _18086_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15298_ _26542_/Q _26150_/Q _15299_/S vssd1 vssd1 vccd1 vccd1 _15298_/X sky130_fd_sc_hd__mux2_1
XFILLER_264_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17037_ _17035_/X _16924_/B _17032_/X input228/X vssd1 vssd1 vccd1 vccd1 _17037_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_116_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14249_ _13084_/A _26395_/Q _14272_/S _14248_/X vssd1 vssd1 vccd1 vccd1 _14249_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _27118_/Q _18748_/X _18986_/X _18987_/X vssd1 vssd1 vccd1 vccd1 _18988_/X
+ sky130_fd_sc_hd__o22a_2
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _17936_/X _17937_/X _18067_/S vssd1 vssd1 vccd1 vccd1 _17939_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20950_ _20950_/A vssd1 vssd1 vccd1 vccd1 _25853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19609_ _27057_/Q _19617_/B _19609_/C vssd1 vssd1 vccd1 vccd1 _19614_/A sky130_fd_sc_hd__and3_1
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20881_ _23696_/A vssd1 vssd1 vccd1 vccd1 _20881_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_242_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22620_ _26323_/Q _22632_/B vssd1 vssd1 vccd1 vccd1 _22620_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22551_ _26297_/Q _22551_/B vssd1 vssd1 vccd1 vccd1 _22551_/Y sky130_fd_sc_hd__nand2_1
XFILLER_250_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21502_ _21502_/A vssd1 vssd1 vccd1 vccd1 _21502_/Y sky130_fd_sc_hd__inv_2
X_25270_ _25270_/A vssd1 vssd1 vccd1 vccd1 _27239_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22482_ _24630_/A vssd1 vssd1 vccd1 vccd1 _22491_/B sky130_fd_sc_hd__clkbuf_1
X_24221_ _26964_/Q _26963_/Q _24221_/C vssd1 vssd1 vccd1 vccd1 _24227_/C sky130_fd_sc_hd__and3_1
X_21433_ _21589_/A vssd1 vssd1 vccd1 vccd1 _21433_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_175_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24152_ _27327_/Q _26941_/Q vssd1 vssd1 vccd1 vccd1 _24157_/C sky130_fd_sc_hd__and2b_1
XFILLER_257_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21364_ _21586_/A vssd1 vssd1 vccd1 vccd1 _21364_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20315_ _25684_/Q _20334_/C _20015_/A vssd1 vssd1 vccd1 vccd1 _20315_/Y sky130_fd_sc_hd__o21ai_1
X_23103_ _26508_/Q _23101_/X _23115_/S vssd1 vssd1 vccd1 vccd1 _23104_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24083_ _26910_/Q _23517_/X _24087_/S vssd1 vssd1 vccd1 vccd1 _24084_/A sky130_fd_sc_hd__mux2_1
X_21295_ _21231_/X _21294_/X _21237_/X vssd1 vssd1 vccd1 vccd1 _21295_/Y sky130_fd_sc_hd__o21bai_2
X_23034_ _23508_/A vssd1 vssd1 vccd1 vccd1 _23034_/X sky130_fd_sc_hd__clkbuf_2
X_20246_ _20179_/X _20245_/X _20186_/X vssd1 vssd1 vccd1 vccd1 _20246_/X sky130_fd_sc_hd__a21o_1
XFILLER_104_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20177_ _20233_/C _20165_/Y _19941_/X _20176_/X vssd1 vssd1 vccd1 vccd1 _20177_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_49_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24985_ _27164_/Q _24913_/X _24984_/Y vssd1 vssd1 vccd1 vccd1 _27164_/D sky130_fd_sc_hd__o21a_1
XFILLER_130_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26724_ _26916_/CLK _26724_/D vssd1 vssd1 vccd1 vccd1 _26724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23936_ _23936_/A vssd1 vssd1 vccd1 vccd1 _26844_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26655_ _26877_/CLK _26655_/D vssd1 vssd1 vccd1 vccd1 _26655_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23867_ _23693_/X _26814_/Q _23871_/S vssd1 vssd1 vccd1 vccd1 _23868_/A sky130_fd_sc_hd__mux2_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13620_ _13410_/X _13616_/X _13619_/X _13071_/A vssd1 vssd1 vccd1 vccd1 _13620_/X
+ sky130_fd_sc_hd__o211a_1
X_25606_ _25607_/CLK _25606_/D vssd1 vssd1 vccd1 vccd1 _25606_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_199_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22818_ _22962_/A _25393_/B vssd1 vssd1 vccd1 vccd1 _22875_/A sky130_fd_sc_hd__nor2_8
X_26586_ _27154_/CLK _26586_/D vssd1 vssd1 vccd1 vccd1 _26586_/Q sky130_fd_sc_hd__dfxtp_4
X_23798_ _23798_/A vssd1 vssd1 vccd1 vccd1 _26783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_260_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25537_ _25545_/CLK _25537_/D vssd1 vssd1 vccd1 vccd1 _25537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13551_ _13552_/A _17821_/B vssd1 vssd1 vccd1 vccd1 _18645_/S sky130_fd_sc_hd__and2_1
X_22749_ _22749_/A vssd1 vssd1 vccd1 vccd1 _26360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16270_ _26543_/Q _26151_/Q _16271_/S vssd1 vssd1 vccd1 vccd1 _16270_/X sky130_fd_sc_hd__mux2_1
X_13482_ _14468_/A vssd1 vssd1 vccd1 vccd1 _13941_/A sky130_fd_sc_hd__clkbuf_2
X_25468_ _27327_/CLK _25468_/D vssd1 vssd1 vccd1 vccd1 _25468_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27207_ _27230_/CLK _27207_/D vssd1 vssd1 vccd1 vccd1 _27207_/Q sky130_fd_sc_hd__dfxtp_1
X_15221_ _27319_/Q _26576_/Q _15221_/S vssd1 vssd1 vccd1 vccd1 _15221_/X sky130_fd_sc_hd__mux2_1
X_24419_ _24434_/A _24932_/A vssd1 vssd1 vccd1 vccd1 _24419_/Y sky130_fd_sc_hd__nand2_1
X_25399_ _25399_/A vssd1 vssd1 vccd1 vccd1 _27296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27138_ _27166_/CLK _27138_/D vssd1 vssd1 vccd1 vccd1 _27138_/Q sky130_fd_sc_hd__dfxtp_1
X_15152_ _16378_/S _15146_/X _15151_/X _15040_/X vssd1 vssd1 vccd1 vccd1 _15152_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14103_ _14520_/S vssd1 vssd1 vccd1 vccd1 _14103_/X sky130_fd_sc_hd__buf_2
X_15083_ _27289_/Q _26482_/Q _15088_/S vssd1 vssd1 vccd1 vccd1 _15083_/X sky130_fd_sc_hd__mux2_1
X_27069_ _27176_/CLK _27069_/D vssd1 vssd1 vccd1 vccd1 _27069_/Q sky130_fd_sc_hd__dfxtp_1
X_19960_ _19956_/X _19957_/Y _19959_/Y vssd1 vssd1 vccd1 vccd1 _19960_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_268_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14034_ _12891_/A _12893_/A _14033_/X _12915_/A _25931_/Q vssd1 vssd1 vccd1 vccd1
+ _14834_/C sky130_fd_sc_hd__o32a_1
X_18911_ _20055_/A _19231_/B vssd1 vssd1 vccd1 vccd1 _18912_/B sky130_fd_sc_hd__nor2_1
XFILLER_180_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19891_ _19879_/X _19889_/X _19890_/X vssd1 vssd1 vccd1 vccd1 _19891_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18842_ _18003_/X _18804_/X _18840_/X _18841_/X vssd1 vssd1 vccd1 vccd1 _18842_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15985_ _26664_/Q _13441_/S _15984_/X _15716_/S vssd1 vssd1 vccd1 vccd1 _15985_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18773_ _19140_/A _19971_/A vssd1 vssd1 vccd1 vccd1 _18773_/X sky130_fd_sc_hd__and2b_1
XTAP_5660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17724_ _25501_/Q _18438_/A _18440_/A _25533_/Q vssd1 vssd1 vccd1 vccd1 _17724_/X
+ sky130_fd_sc_hd__a22o_1
X_14936_ _15706_/B _15706_/C _14936_/C vssd1 vssd1 vccd1 vccd1 _15954_/C sky130_fd_sc_hd__nor3_1
XFILLER_94_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_wb_clk_i clkbuf_opt_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26881_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14867_ _12750_/A _14865_/X _14866_/X vssd1 vssd1 vccd1 vccd1 _14867_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17655_ _20249_/A _17635_/X _17608_/A _17654_/Y vssd1 vssd1 vccd1 vccd1 _17656_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_263_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13818_ _13818_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13818_/Y sky130_fd_sc_hd__nor2_4
X_16606_ _19187_/A _19191_/B vssd1 vssd1 vccd1 vccd1 _16606_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_17_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17586_ _16591_/A _17584_/X _17572_/X _17585_/X vssd1 vssd1 vccd1 vccd1 _17587_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_250_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14798_ _25827_/Q _27261_/Q _14813_/S vssd1 vssd1 vccd1 vccd1 _14798_/X sky130_fd_sc_hd__mux2_1
XFILLER_251_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19325_ _19325_/A vssd1 vssd1 vccd1 vccd1 _19325_/Y sky130_fd_sc_hd__inv_2
X_16537_ _14794_/X _16532_/X _16536_/X _17181_/A vssd1 vssd1 vccd1 vccd1 _16537_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_259_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13749_ _25910_/Q _12902_/A _13570_/A _13748_/Y vssd1 vssd1 vccd1 vccd1 _14486_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_232_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19256_ _19256_/A _19256_/B vssd1 vssd1 vccd1 vccd1 _19256_/Y sky130_fd_sc_hd__nand2_1
X_16468_ _16498_/S vssd1 vssd1 vccd1 vccd1 _16500_/S sky130_fd_sc_hd__buf_2
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18207_ _18206_/X _18081_/X _18210_/S vssd1 vssd1 vccd1 vccd1 _18207_/X sky130_fd_sc_hd__mux2_1
X_15419_ _15406_/X _25849_/Q _26049_/Q _16443_/S _15318_/A vssd1 vssd1 vccd1 vccd1
+ _15419_/X sky130_fd_sc_hd__a221o_1
X_19187_ _19187_/A _19191_/B vssd1 vssd1 vccd1 vccd1 _19187_/X sky130_fd_sc_hd__xor2_4
X_16399_ _25856_/Q _26056_/Q _16399_/S vssd1 vssd1 vccd1 vccd1 _16399_/X sky130_fd_sc_hd__mux2_1
XFILLER_275_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18138_ _18138_/A _18138_/B vssd1 vssd1 vccd1 vccd1 _18381_/A sky130_fd_sc_hd__nor2_1
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18069_ _17934_/X _17949_/X _18070_/S vssd1 vssd1 vccd1 vccd1 _18069_/X sky130_fd_sc_hd__mux2_1
XFILLER_208_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20100_ _20100_/A vssd1 vssd1 vccd1 vccd1 _20100_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21080_ _21080_/A vssd1 vssd1 vccd1 vccd1 _25902_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20031_ _22500_/A _20030_/B _19738_/X vssd1 vssd1 vccd1 vccd1 _20031_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_86_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24770_ _24770_/A _24770_/B vssd1 vssd1 vccd1 vccd1 _27099_/D sky130_fd_sc_hd__nor2_1
X_21982_ _21982_/A vssd1 vssd1 vccd1 vccd1 _26104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23721_ _23721_/A vssd1 vssd1 vccd1 vccd1 _26758_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20933_ _25848_/Q _20932_/X _20933_/S vssd1 vssd1 vccd1 vccd1 _20934_/A sky130_fd_sc_hd__mux2_1
XFILLER_270_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26440_ _26796_/CLK _26440_/D vssd1 vssd1 vccd1 vccd1 _26440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23652_ _26733_/Q _23565_/X _23656_/S vssd1 vssd1 vccd1 vccd1 _23653_/A sky130_fd_sc_hd__mux2_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20864_ _25828_/Q vssd1 vssd1 vccd1 vccd1 _20865_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_26_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22603_ _22593_/X _22602_/Y _22600_/X vssd1 vssd1 vccd1 vccd1 _26316_/D sky130_fd_sc_hd__a21oi_1
X_26371_ _26467_/CLK _26371_/D vssd1 vssd1 vccd1 vccd1 _26371_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_224_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23583_ _23583_/A vssd1 vssd1 vccd1 vccd1 _26706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20795_ _20795_/A vssd1 vssd1 vccd1 vccd1 _25792_/D sky130_fd_sc_hd__clkbuf_1
X_25322_ _25378_/A vssd1 vssd1 vccd1 vccd1 _25391_/S sky130_fd_sc_hd__buf_8
XFILLER_23_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22534_ _22534_/A vssd1 vssd1 vccd1 vccd1 _26291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25253_ _25253_/A vssd1 vssd1 vccd1 vccd1 _27231_/D sky130_fd_sc_hd__clkbuf_1
X_22465_ _26258_/Q _22470_/B vssd1 vssd1 vccd1 vccd1 _22465_/X sky130_fd_sc_hd__or2_1
XFILLER_194_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24204_ _24222_/A _24204_/B _24205_/B vssd1 vssd1 vccd1 vccd1 _26958_/D sky130_fd_sc_hd__nor3_1
XFILLER_136_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21416_ _25481_/Q _21416_/B vssd1 vssd1 vccd1 vccd1 _21416_/X sky130_fd_sc_hd__or2_1
X_25184_ _27202_/Q _25217_/A _25179_/A vssd1 vssd1 vccd1 vccd1 _25184_/Y sky130_fd_sc_hd__o21ai_1
X_22396_ _22340_/S _22381_/X _22392_/X _22395_/Y _22379_/X vssd1 vssd1 vccd1 vccd1
+ _22396_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_175_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24135_ _24135_/A vssd1 vssd1 vccd1 vccd1 _26933_/D sky130_fd_sc_hd__clkbuf_1
X_21347_ _21284_/A _18576_/X _21286_/A _25805_/Q _21346_/X vssd1 vssd1 vccd1 vccd1
+ _21347_/X sky130_fd_sc_hd__a221o_1
XFILLER_123_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24066_ _26903_/Q _23597_/X _24070_/S vssd1 vssd1 vccd1 vccd1 _24067_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21278_ _21278_/A vssd1 vssd1 vccd1 vccd1 _21278_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_23017_ _26480_/Q _22720_/X _23017_/S vssd1 vssd1 vccd1 vccd1 _23018_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20229_ _20679_/A _19727_/X _20228_/Y _19920_/A vssd1 vssd1 vccd1 vccd1 _20259_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_270_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15770_ _13335_/A _15767_/X _15769_/X _13340_/A vssd1 vssd1 vccd1 vccd1 _15770_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _12982_/A _13577_/A vssd1 vssd1 vccd1 vccd1 _20487_/C sky130_fd_sc_hd__nor2_2
X_24968_ _27156_/Q _24957_/X _24967_/Y vssd1 vssd1 vccd1 vccd1 _27156_/D sky130_fd_sc_hd__o21a_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _25754_/Q vssd1 vssd1 vccd1 vccd1 _20701_/A sky130_fd_sc_hd__inv_4
XFILLER_233_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26707_ _26931_/CLK _26707_/D vssd1 vssd1 vccd1 vccd1 _26707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23919_ _23919_/A vssd1 vssd1 vccd1 vccd1 _26837_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24899_ _25206_/D vssd1 vssd1 vccd1 vccd1 _24900_/D sky130_fd_sc_hd__clkinv_2
XFILLER_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _25564_/Q _17438_/B _17414_/X vssd1 vssd1 vccd1 vccd1 _17440_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_217_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26638_ _26823_/CLK _26638_/D vssd1 vssd1 vccd1 vccd1 _26638_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _26874_/Q _25788_/Q _14652_/S vssd1 vssd1 vccd1 vccd1 _14652_/X sky130_fd_sc_hd__mux2_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13603_ _27240_/Q _15972_/B vssd1 vssd1 vccd1 vccd1 _13603_/X sky130_fd_sc_hd__or2_1
XFILLER_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _17380_/A _17371_/B _17372_/B vssd1 vssd1 vccd1 vccd1 _25542_/D sky130_fd_sc_hd__nor3_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26569_ _26797_/CLK _26569_/D vssd1 vssd1 vccd1 vccd1 _26569_/Q sky130_fd_sc_hd__dfxtp_1
X_14583_ _16204_/S vssd1 vssd1 vccd1 vccd1 _16368_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_201_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19110_ _19122_/B _19110_/B vssd1 vssd1 vccd1 vccd1 _19576_/C sky130_fd_sc_hd__nand2_2
XFILLER_41_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16322_ _26805_/Q _26449_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _16322_/X sky130_fd_sc_hd__mux2_1
X_13534_ _26074_/Q _25879_/Q _13534_/S vssd1 vssd1 vccd1 vccd1 _13534_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19041_ _19317_/A _19041_/B vssd1 vssd1 vccd1 vccd1 _19041_/Y sky130_fd_sc_hd__nand2_1
XFILLER_185_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16253_ _14742_/A _25781_/Q _16361_/S _26867_/Q _15308_/S vssd1 vssd1 vccd1 vccd1
+ _16253_/X sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_147_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27176_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13465_ _13465_/A vssd1 vssd1 vccd1 vccd1 _13466_/A sky130_fd_sc_hd__buf_6
XFILLER_199_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15204_ _26120_/Q _26021_/Q _16436_/S vssd1 vssd1 vccd1 vccd1 _15204_/X sky130_fd_sc_hd__mux2_1
X_16184_ _16174_/X _16177_/X _16180_/X _16183_/X _14757_/A _14778_/A vssd1 vssd1 vccd1
+ vccd1 _16185_/B sky130_fd_sc_hd__mux4_1
XFILLER_154_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13396_ _25912_/Q _13737_/A _13395_/Y _25795_/Q vssd1 vssd1 vccd1 vccd1 _13397_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15135_ _15135_/A vssd1 vssd1 vccd1 vccd1 _15135_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15066_ _15065_/X _26710_/Q _26838_/Q _16385_/S _14688_/A vssd1 vssd1 vccd1 vccd1
+ _15066_/X sky130_fd_sc_hd__a221o_1
X_19943_ _20189_/A _19943_/B vssd1 vssd1 vccd1 vccd1 _19968_/A sky130_fd_sc_hd__or2_1
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14017_ _13999_/X _14016_/X _13173_/A vssd1 vssd1 vccd1 vccd1 _14017_/X sky130_fd_sc_hd__a21o_2
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19874_ _21718_/A vssd1 vssd1 vccd1 vccd1 _19874_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18825_ _18825_/A vssd1 vssd1 vccd1 vccd1 _18825_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18756_ _18756_/A vssd1 vssd1 vccd1 vccd1 _18756_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15968_ _26340_/Q _26600_/Q _15988_/S vssd1 vssd1 vccd1 vccd1 _15968_/X sky130_fd_sc_hd__mux2_1
XFILLER_255_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17707_ _17708_/A _19847_/A _24342_/A vssd1 vssd1 vccd1 vccd1 _17735_/A sky130_fd_sc_hd__a21o_1
X_14919_ _14755_/A _14916_/X _14918_/X _14804_/A vssd1 vssd1 vccd1 vccd1 _14919_/X
+ sky130_fd_sc_hd__a211o_1
X_15899_ _14107_/X _15897_/X _15898_/X _13141_/A vssd1 vssd1 vccd1 vccd1 _15899_/X
+ sky130_fd_sc_hd__a211o_1
X_18687_ _13381_/Y _19393_/B _18685_/X _18269_/A _18686_/Y vssd1 vssd1 vccd1 vccd1
+ _18687_/X sky130_fd_sc_hd__a221o_1
XFILLER_247_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17638_ _17650_/A _17638_/B vssd1 vssd1 vccd1 vccd1 _25591_/D sky130_fd_sc_hd__nor2_1
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17569_ _25911_/Q _17568_/X _13573_/B _17525_/X vssd1 vssd1 vccd1 vccd1 _17569_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_19308_ _18806_/X _19298_/X _19307_/X vssd1 vssd1 vccd1 vccd1 _19308_/X sky130_fd_sc_hd__a21o_4
XFILLER_17_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20580_ _23754_/A vssd1 vssd1 vccd1 vccd1 _20580_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19239_ _19235_/B _19576_/D _18636_/A vssd1 vssd1 vccd1 vccd1 _19239_/X sky130_fd_sc_hd__o21a_1
XFILLER_164_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22250_ _26195_/Q _22249_/X _22238_/X _26296_/Q _22241_/X vssd1 vssd1 vccd1 vccd1
+ _22250_/X sky130_fd_sc_hd__a221o_1
XFILLER_219_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21201_ _21309_/A vssd1 vssd1 vccd1 vccd1 _21202_/A sky130_fd_sc_hd__buf_4
X_22181_ _22195_/A vssd1 vssd1 vccd1 vccd1 _22181_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21132_ _25917_/Q _21130_/X _21131_/X input16/X vssd1 vssd1 vccd1 vccd1 _21133_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_235_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25940_ _27058_/CLK _25940_/D vssd1 vssd1 vccd1 vccd1 _25940_/Q sky130_fd_sc_hd__dfxtp_1
X_21063_ _25900_/Q _20970_/X _21063_/S vssd1 vssd1 vccd1 vccd1 _21064_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20014_ _20014_/A _20080_/B vssd1 vssd1 vccd1 vccd1 _20014_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25871_ _27265_/CLK _25871_/D vssd1 vssd1 vccd1 vccd1 _25871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24822_ _27111_/Q _24837_/B vssd1 vssd1 vccd1 vccd1 _24822_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24753_ _24764_/A _24753_/B vssd1 vssd1 vccd1 vccd1 _27094_/D sky130_fd_sc_hd__nor2_1
X_21965_ _21965_/A vssd1 vssd1 vccd1 vccd1 _26096_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23704_ _23702_/X _26753_/Q _23716_/S vssd1 vssd1 vccd1 vccd1 _23705_/A sky130_fd_sc_hd__mux2_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ _23731_/A vssd1 vssd1 vccd1 vccd1 _20916_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_214_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24684_ _24699_/A _24684_/B vssd1 vssd1 vccd1 vccd1 _27078_/D sky130_fd_sc_hd__nor2_1
X_21896_ _20500_/X _26066_/Q _21900_/S vssd1 vssd1 vccd1 vccd1 _21897_/A sky130_fd_sc_hd__mux2_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26423_ _26913_/CLK _26423_/D vssd1 vssd1 vccd1 vccd1 _26423_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23635_ _23635_/A vssd1 vssd1 vccd1 vccd1 _26725_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20847_ _20847_/A vssd1 vssd1 vccd1 vccd1 _25819_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26354_ _27292_/CLK _26354_/D vssd1 vssd1 vccd1 vccd1 _26354_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_168_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23566_ _26701_/Q _23565_/X _23572_/S vssd1 vssd1 vccd1 vccd1 _23567_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20778_ _20778_/A vssd1 vssd1 vccd1 vccd1 _25784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25305_ _25305_/A vssd1 vssd1 vccd1 vccd1 _27255_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22517_ _22517_/A vssd1 vssd1 vccd1 vccd1 _26282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26285_ _26286_/CLK _26285_/D vssd1 vssd1 vccd1 vccd1 _26285_/Q sky130_fd_sc_hd__dfxtp_1
X_23497_ _23497_/A vssd1 vssd1 vccd1 vccd1 _26678_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13250_ _13250_/A vssd1 vssd1 vccd1 vccd1 _13937_/A sky130_fd_sc_hd__buf_2
X_25236_ _27224_/Q _25225_/X _25228_/X _24751_/B _25235_/X vssd1 vssd1 vccd1 vccd1
+ _27224_/D sky130_fd_sc_hd__o221a_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22448_ _26251_/Q _22457_/B vssd1 vssd1 vccd1 vccd1 _22448_/X sky130_fd_sc_hd__or2_1
XFILLER_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25167_ _25691_/Q _25065_/A _25139_/A _25166_/Y _25024_/A vssd1 vssd1 vccd1 vccd1
+ _25167_/X sky130_fd_sc_hd__a221o_1
X_13181_ _14566_/A vssd1 vssd1 vccd1 vccd1 _14833_/A sky130_fd_sc_hd__buf_2
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22379_ _22379_/A vssd1 vssd1 vccd1 vccd1 _22379_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24118_ _26926_/Q _23568_/X _24120_/S vssd1 vssd1 vccd1 vccd1 _24119_/A sky130_fd_sc_hd__mux2_1
XFILLER_269_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25098_ _22507_/A _25092_/X _25087_/X _16637_/C _25079_/X vssd1 vssd1 vccd1 vccd1
+ _25098_/X sky130_fd_sc_hd__a221o_1
XFILLER_145_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16940_ _16940_/A _16954_/A vssd1 vssd1 vccd1 vccd1 _16940_/Y sky130_fd_sc_hd__nand2_1
X_24049_ _24049_/A vssd1 vssd1 vccd1 vccd1 _26895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16871_ _16871_/A vssd1 vssd1 vccd1 vccd1 _16871_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18610_ _27208_/Q _19364_/B vssd1 vssd1 vccd1 vccd1 _18610_/X sky130_fd_sc_hd__and2_1
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15822_ _13085_/A _26890_/Q _26762_/Q _15734_/S vssd1 vssd1 vccd1 vccd1 _15822_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_219_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19590_ _19887_/B vssd1 vssd1 vccd1 vccd1 _19779_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15753_ _15932_/A _15753_/B vssd1 vssd1 vccd1 vccd1 _15753_/X sky130_fd_sc_hd__or2_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18541_ _18541_/A _19289_/B vssd1 vssd1 vccd1 vccd1 _18541_/X sky130_fd_sc_hd__or2_1
X_12965_ _13933_/A vssd1 vssd1 vccd1 vccd1 _13803_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_80 _23702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_91 _24871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14704_ _14956_/A _14704_/B vssd1 vssd1 vccd1 vccd1 _14704_/Y sky130_fd_sc_hd__nand2_1
XFILLER_205_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18472_ _19374_/B _19800_/A vssd1 vssd1 vccd1 vccd1 _18474_/B sky130_fd_sc_hd__and2b_1
X_15684_ _15406_/A _25845_/Q _26045_/Q _15674_/X _13281_/A vssd1 vssd1 vccd1 vccd1
+ _15684_/X sky130_fd_sc_hd__a221o_1
X_12896_ _14033_/S vssd1 vssd1 vccd1 vccd1 _14402_/S sky130_fd_sc_hd__buf_4
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _25559_/Q vssd1 vssd1 vccd1 vccd1 _17427_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14635_ _15014_/S vssd1 vssd1 vccd1 vccd1 _14953_/S sky130_fd_sc_hd__buf_2
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _17382_/A _17360_/C vssd1 vssd1 vccd1 vccd1 _17354_/Y sky130_fd_sc_hd__nor2_1
XFILLER_220_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14566_ _14566_/A _14566_/B vssd1 vssd1 vccd1 vccd1 _17983_/A sky130_fd_sc_hd__or2_2
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13517_ _15292_/A vssd1 vssd1 vccd1 vccd1 _15857_/S sky130_fd_sc_hd__buf_2
XFILLER_147_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16305_ _16305_/A vssd1 vssd1 vccd1 vccd1 _16323_/S sky130_fd_sc_hd__buf_2
X_17285_ _17285_/A _17293_/C vssd1 vssd1 vccd1 vccd1 _17285_/Y sky130_fd_sc_hd__nor2_1
X_14497_ _14497_/A vssd1 vssd1 vccd1 vccd1 _15726_/S sky130_fd_sc_hd__buf_4
XFILLER_174_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19024_ _27151_/Q _19302_/B vssd1 vssd1 vccd1 vccd1 _19024_/X sky130_fd_sc_hd__or2_1
X_16236_ _27254_/Q _16388_/B vssd1 vssd1 vccd1 vccd1 _16236_/X sky130_fd_sc_hd__or2_1
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13448_ _26630_/Q _26726_/Q _15800_/S vssd1 vssd1 vccd1 vccd1 _13448_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16167_ _16167_/A _16167_/B vssd1 vssd1 vccd1 vccd1 _16167_/X sky130_fd_sc_hd__or2_1
X_13379_ _19947_/A _15615_/S _13378_/Y vssd1 vssd1 vccd1 vccd1 _17824_/B sky130_fd_sc_hd__a21oi_4
XFILLER_170_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15118_ _26546_/Q _26154_/Q _15119_/S vssd1 vssd1 vccd1 vccd1 _15118_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_141_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16098_ _15676_/X _26347_/Q _26607_/Q _16273_/S _15672_/A vssd1 vssd1 vccd1 vccd1
+ _16098_/X sky130_fd_sc_hd__a221o_1
XFILLER_69_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15049_ _12774_/A _26902_/Q _26774_/Q _16377_/S _15048_/X vssd1 vssd1 vccd1 vccd1
+ _15049_/X sky130_fd_sc_hd__a221o_1
X_19926_ _19926_/A vssd1 vssd1 vccd1 vccd1 _19926_/X sky130_fd_sc_hd__buf_2
XFILLER_141_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_wb_clk_i clkbuf_opt_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27280_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_269_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19857_ _19736_/B _19853_/X _19854_/Y _19855_/X _19856_/Y vssd1 vssd1 vccd1 vccd1
+ _19981_/A sky130_fd_sc_hd__o2111a_2
XFILLER_69_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18808_ _18808_/A vssd1 vssd1 vccd1 vccd1 _18808_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19788_ _19784_/Y _19785_/Y _20323_/B vssd1 vssd1 vccd1 vccd1 _19788_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_110_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18739_ _18359_/X _18728_/X _18737_/X _18738_/X vssd1 vssd1 vccd1 vccd1 _18739_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_271_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21750_ _20542_/X _26009_/Q _21754_/S vssd1 vssd1 vccd1 vccd1 _21751_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20701_ _20701_/A _20703_/B vssd1 vssd1 vccd1 vccd1 _20701_/Y sky130_fd_sc_hd__nand2_1
XFILLER_224_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21681_ _25980_/Q input192/X _21685_/S vssd1 vssd1 vccd1 vccd1 _21682_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23420_ _23420_/A vssd1 vssd1 vccd1 vccd1 _26644_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_260_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20632_ _26264_/Q _17190_/X _20630_/X _20631_/X vssd1 vssd1 vccd1 vccd1 _25727_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_211_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23351_ _20601_/X _26614_/Q _23357_/S vssd1 vssd1 vccd1 vccd1 _23352_/A sky130_fd_sc_hd__mux2_1
X_20563_ _23741_/A vssd1 vssd1 vccd1 vccd1 _20563_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_221_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22302_ _26212_/Q _22294_/X _22300_/X _26313_/Q _22301_/X vssd1 vssd1 vccd1 vccd1
+ _22302_/X sky130_fd_sc_hd__a221o_1
XFILLER_192_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26070_ _26594_/CLK _26070_/D vssd1 vssd1 vccd1 vccd1 _26070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23282_ _23282_/A vssd1 vssd1 vccd1 vccd1 _26583_/D sky130_fd_sc_hd__clkbuf_1
X_20494_ _20494_/A vssd1 vssd1 vccd1 vccd1 _25692_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25021_ _20630_/A _25003_/X _25020_/X vssd1 vssd1 vccd1 vccd1 _25021_/Y sky130_fd_sc_hd__o21ai_1
X_22233_ _22239_/A _22239_/B vssd1 vssd1 vccd1 vccd1 _22315_/A sky130_fd_sc_hd__nor2_2
XFILLER_180_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22164_ _22195_/A vssd1 vssd1 vccd1 vccd1 _22164_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21115_ _21118_/A _21115_/B vssd1 vssd1 vccd1 vccd1 _21116_/A sky130_fd_sc_hd__or2_1
XFILLER_132_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26972_ _26974_/CLK _26972_/D vssd1 vssd1 vccd1 vccd1 _26972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22095_ _26155_/Q _20958_/X _22099_/S vssd1 vssd1 vccd1 vccd1 _22096_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21046_ _25892_/Q _20945_/X _21048_/S vssd1 vssd1 vccd1 vccd1 _21047_/A sky130_fd_sc_hd__mux2_1
X_25923_ _27213_/CLK _25923_/D vssd1 vssd1 vccd1 vccd1 _25923_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_86_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25854_ _27288_/CLK _25854_/D vssd1 vssd1 vccd1 vccd1 _25854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_274_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24805_ _24803_/Y _24804_/X _24796_/X vssd1 vssd1 vccd1 vccd1 _27106_/D sky130_fd_sc_hd__a21oi_1
XFILLER_262_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25785_ _27257_/CLK _25785_/D vssd1 vssd1 vccd1 vccd1 _25785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22997_ _23019_/A vssd1 vssd1 vccd1 vccd1 _23006_/S sky130_fd_sc_hd__buf_4
XFILLER_262_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _12750_/A vssd1 vssd1 vccd1 vccd1 _12751_/A sky130_fd_sc_hd__clkbuf_4
X_24736_ _24739_/A _24736_/B vssd1 vssd1 vccd1 vccd1 _24736_/Y sky130_fd_sc_hd__nand2_4
XFILLER_216_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21948_ _21948_/A vssd1 vssd1 vccd1 vccd1 _26089_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12681_ _13185_/A vssd1 vssd1 vccd1 vccd1 _13215_/A sky130_fd_sc_hd__clkbuf_4
X_24667_ _24923_/A vssd1 vssd1 vccd1 vccd1 _24668_/B sky130_fd_sc_hd__inv_2
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21879_ _21867_/Y _21876_/X _21877_/X _21878_/X vssd1 vssd1 vccd1 vccd1 _26062_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26406_ _26467_/CLK _26406_/D vssd1 vssd1 vccd1 vccd1 _26406_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_230_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14420_ _13134_/A _14418_/X _14419_/X _14522_/S vssd1 vssd1 vccd1 vccd1 _14421_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_199_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23618_ _23618_/A vssd1 vssd1 vccd1 vccd1 _26717_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24598_ hold2/A _24608_/B vssd1 vssd1 vccd1 vccd1 _24598_/Y sky130_fd_sc_hd__nand2_1
X_26337_ _26433_/CLK _26337_/D vssd1 vssd1 vccd1 vccd1 _26337_/Q sky130_fd_sc_hd__dfxtp_2
X_14351_ _26522_/Q _26130_/Q _14351_/S vssd1 vssd1 vccd1 vccd1 _14351_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23549_ _23549_/A vssd1 vssd1 vccd1 vccd1 _23549_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_195_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13302_ _13365_/A vssd1 vssd1 vccd1 vccd1 _14077_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_155_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17070_ _25978_/Q _17061_/A _16999_/X _17015_/X vssd1 vssd1 vccd1 vccd1 _17070_/X
+ sky130_fd_sc_hd__a22o_4
X_26268_ _26271_/CLK _26268_/D vssd1 vssd1 vccd1 vccd1 _26268_/Q sky130_fd_sc_hd__dfxtp_1
X_14282_ _25575_/Q _14187_/A _14193_/B vssd1 vssd1 vccd1 vccd1 _14282_/Y sky130_fd_sc_hd__o21ai_1
X_16021_ _25809_/Q _27243_/Q _16021_/S vssd1 vssd1 vccd1 vccd1 _16022_/B sky130_fd_sc_hd__mux2_1
XFILLER_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25219_ _25219_/A vssd1 vssd1 vccd1 vccd1 _25219_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13233_ _15924_/A vssd1 vssd1 vccd1 vccd1 _16111_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_237_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26199_ _26250_/CLK _26199_/D vssd1 vssd1 vccd1 vccd1 _26199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13164_ _13164_/A vssd1 vssd1 vccd1 vccd1 _14677_/A sky130_fd_sc_hd__buf_4
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13095_ _26107_/Q _26008_/Q _15467_/S vssd1 vssd1 vccd1 vccd1 _13095_/X sky130_fd_sc_hd__mux2_1
X_17972_ _17970_/X _17971_/X _17978_/A _17219_/A vssd1 vssd1 vccd1 vccd1 _18186_/A
+ sky130_fd_sc_hd__a211o_2
X_19711_ _19675_/A _19675_/B _19710_/Y vssd1 vssd1 vccd1 vccd1 _19712_/B sky130_fd_sc_hd__o21ai_1
X_16923_ _16907_/X _16973_/C _16922_/X vssd1 vssd1 vccd1 vccd1 _16924_/B sky130_fd_sc_hd__o21a_2
XFILLER_238_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19642_ _24848_/A vssd1 vssd1 vccd1 vccd1 _19642_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_77_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16854_ _16983_/B vssd1 vssd1 vccd1 vccd1 _16855_/A sky130_fd_sc_hd__buf_2
XFILLER_238_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _26502_/Q _26374_/Q _15805_/S vssd1 vssd1 vccd1 vccd1 _15805_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19573_ _19573_/A _19573_/B _19573_/C _18328_/X vssd1 vssd1 vccd1 vccd1 _19574_/C
+ sky130_fd_sc_hd__or4b_2
XFILLER_92_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13997_ _13995_/X _13996_/X _14010_/S vssd1 vssd1 vccd1 vccd1 _13997_/X sky130_fd_sc_hd__mux2_1
X_16785_ _21709_/B vssd1 vssd1 vccd1 vccd1 _16785_/Y sky130_fd_sc_hd__inv_2
XFILLER_281_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18524_ _18437_/X _18502_/X _18523_/X vssd1 vssd1 vccd1 vccd1 _18524_/X sky130_fd_sc_hd__a21o_4
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_opt_2_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_15736_ _25812_/Q _13441_/S _15970_/S _15735_/X vssd1 vssd1 vccd1 vccd1 _15736_/X
+ sky130_fd_sc_hd__o211a_1
X_12948_ _13916_/B _13916_/C _12948_/C vssd1 vssd1 vccd1 vccd1 _12948_/Y sky130_fd_sc_hd__nand3_1
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_162_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27122_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18455_ _18455_/A vssd1 vssd1 vccd1 vccd1 _18455_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_261_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12879_ _25471_/Q _25470_/Q _12975_/B vssd1 vssd1 vccd1 vccd1 _12946_/A sky130_fd_sc_hd__nor3_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15667_ _16348_/S _15665_/X _15666_/X _13274_/X vssd1 vssd1 vccd1 vccd1 _15668_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17406_ _17408_/A _17408_/C _17405_/Y vssd1 vssd1 vccd1 vccd1 _25553_/D sky130_fd_sc_hd__o21a_1
XFILLER_222_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14618_ _14618_/A vssd1 vssd1 vccd1 vccd1 _14618_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15598_ _13532_/X _15595_/X _15597_/X _13291_/A vssd1 vssd1 vccd1 vccd1 _15598_/X
+ sky130_fd_sc_hd__o211a_1
X_18386_ _18666_/A _18386_/B vssd1 vssd1 vccd1 vccd1 _18386_/Y sky130_fd_sc_hd__nor2_1
XFILLER_221_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17337_ _17336_/X _17341_/C _17318_/X vssd1 vssd1 vccd1 vccd1 _17337_/Y sky130_fd_sc_hd__a21oi_1
X_14549_ _13540_/A _14545_/X _14548_/X _13210_/A vssd1 vssd1 vccd1 vccd1 _14549_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17268_ _25511_/Q vssd1 vssd1 vccd1 vccd1 _17268_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19007_ _19352_/A vssd1 vssd1 vccd1 vccd1 _19007_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16219_ _26119_/Q _26020_/Q _16240_/S vssd1 vssd1 vccd1 vccd1 _16219_/X sky130_fd_sc_hd__mux2_1
X_17199_ _25493_/Q _17151_/X _17146_/X _19774_/A vssd1 vssd1 vccd1 vccd1 _17200_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19909_ _25734_/Q vssd1 vssd1 vccd1 vccd1 _20650_/A sky130_fd_sc_hd__buf_8
XFILLER_257_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22920_ _22920_/A vssd1 vssd1 vccd1 vccd1 _26436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22851_ _26406_/Q _22688_/X _22851_/S vssd1 vssd1 vccd1 vccd1 _22852_/A sky130_fd_sc_hd__mux2_1
XFILLER_256_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21802_ _21802_/A vssd1 vssd1 vccd1 vccd1 _26031_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25570_ _25596_/CLK _25570_/D vssd1 vssd1 vccd1 vccd1 _25570_/Q sky130_fd_sc_hd__dfxtp_1
X_22782_ _22782_/A vssd1 vssd1 vccd1 vccd1 _26375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24521_ _24370_/S _25626_/Q _24520_/X vssd1 vssd1 vccd1 vccd1 _24978_/A sky130_fd_sc_hd__o21ai_4
X_21733_ _21733_/A vssd1 vssd1 vccd1 vccd1 _26001_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27240_ _27301_/CLK _27240_/D vssd1 vssd1 vccd1 vccd1 _27240_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24452_ _24464_/A _24590_/A vssd1 vssd1 vccd1 vccd1 _24452_/Y sky130_fd_sc_hd__nand2_1
XFILLER_169_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21664_ _21698_/A vssd1 vssd1 vccd1 vccd1 _23289_/S sky130_fd_sc_hd__clkbuf_2
X_23403_ _23403_/A vssd1 vssd1 vccd1 vccd1 _26636_/D sky130_fd_sc_hd__clkbuf_1
X_20615_ _20615_/A vssd1 vssd1 vccd1 vccd1 _25721_/D sky130_fd_sc_hd__clkbuf_1
X_27171_ _27173_/CLK _27171_/D vssd1 vssd1 vccd1 vccd1 _27171_/Q sky130_fd_sc_hd__dfxtp_1
X_24383_ _24474_/A vssd1 vssd1 vccd1 vccd1 _24383_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21595_ _21552_/X _21566_/X _21594_/Y _21581_/X vssd1 vssd1 vccd1 vccd1 _21595_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_137_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26122_ _26483_/CLK _26122_/D vssd1 vssd1 vccd1 vccd1 _26122_/Q sky130_fd_sc_hd__dfxtp_1
X_23334_ _23334_/A vssd1 vssd1 vccd1 vccd1 _26606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20546_ _23728_/A vssd1 vssd1 vccd1 vccd1 _20546_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26053_ _27329_/A _26053_/D vssd1 vssd1 vccd1 vccd1 _26053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23265_ _23265_/A vssd1 vssd1 vccd1 vccd1 _26575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20477_ _20457_/B _20460_/B _20457_/A vssd1 vssd1 vccd1 vccd1 _20478_/B sky130_fd_sc_hd__a21boi_1
XFILLER_146_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25004_ _25114_/A vssd1 vssd1 vccd1 vccd1 _25004_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22216_ _24441_/A vssd1 vssd1 vccd1 vccd1 _22288_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_145_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23196_ _23196_/A vssd1 vssd1 vccd1 vccd1 _23205_/S sky130_fd_sc_hd__buf_6
XFILLER_106_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22147_ _26167_/Q _22113_/X _22115_/X _22146_/X _22137_/X vssd1 vssd1 vccd1 vccd1
+ _22147_/X sky130_fd_sc_hd__a221o_1
XFILLER_106_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput380 _17026_/X vssd1 vssd1 vccd1 vccd1 din0[13] sky130_fd_sc_hd__buf_2
XFILLER_267_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput391 _17040_/X vssd1 vssd1 vccd1 vccd1 din0[23] sky130_fd_sc_hd__buf_2
XFILLER_117_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26955_ _26992_/CLK _26955_/D vssd1 vssd1 vccd1 vccd1 _26955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22078_ _22078_/A vssd1 vssd1 vccd1 vccd1 _26147_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13920_ input121/X input156/X _14320_/S vssd1 vssd1 vccd1 vccd1 _13921_/B sky130_fd_sc_hd__mux2_8
X_21029_ _25884_/Q _20919_/X _21037_/S vssd1 vssd1 vccd1 vccd1 _21030_/A sky130_fd_sc_hd__mux2_1
X_25906_ _26278_/CLK _25906_/D vssd1 vssd1 vccd1 vccd1 _25906_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_75_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26886_ _27278_/CLK _26886_/D vssd1 vssd1 vccd1 vccd1 _26886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13851_ _13638_/A _23533_/A _13850_/Y _13683_/X vssd1 vssd1 vccd1 vccd1 _19824_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_19_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25837_ _27307_/CLK _25837_/D vssd1 vssd1 vccd1 vccd1 _25837_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12802_ _25579_/Q _25577_/Q _14188_/A vssd1 vssd1 vccd1 vccd1 _14189_/A sky130_fd_sc_hd__or3b_1
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13782_ _14727_/A _13780_/X _13781_/X _13479_/A vssd1 vssd1 vccd1 vccd1 _13787_/B
+ sky130_fd_sc_hd__o211a_1
X_16570_ _19240_/S _16573_/A vssd1 vssd1 vccd1 vccd1 _16571_/A sky130_fd_sc_hd__nor2_1
XFILLER_74_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_408 _17046_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_25768_ _27277_/CLK _25768_/D vssd1 vssd1 vccd1 vccd1 _25768_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_419 _17099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15521_ _15521_/A _15521_/B vssd1 vssd1 vccd1 vccd1 _15521_/Y sky130_fd_sc_hd__nor2_1
X_12733_ _25580_/Q vssd1 vssd1 vccd1 vccd1 _13249_/A sky130_fd_sc_hd__inv_2
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24719_ _24725_/A _24719_/B vssd1 vssd1 vccd1 vccd1 _24719_/Y sky130_fd_sc_hd__nand2_2
X_25699_ _26595_/CLK _25699_/D vssd1 vssd1 vccd1 vccd1 _25699_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18240_ _18454_/A vssd1 vssd1 vccd1 vccd1 _18565_/A sky130_fd_sc_hd__clkbuf_2
X_15452_ _15448_/X _15451_/X _15646_/A vssd1 vssd1 vccd1 vccd1 _15452_/X sky130_fd_sc_hd__mux2_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14403_ _14403_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14404_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18171_ _26943_/Q _18826_/A _18827_/A _26975_/Q vssd1 vssd1 vccd1 vccd1 _18171_/X
+ sky130_fd_sc_hd__a22o_1
X_15383_ _26116_/Q _26017_/Q _16053_/S vssd1 vssd1 vccd1 vccd1 _15383_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14334_ _14331_/X _14332_/X _14333_/X _14272_/S vssd1 vssd1 vccd1 vccd1 _14334_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17122_ _17635_/A vssd1 vssd1 vccd1 vccd1 _20689_/A sky130_fd_sc_hd__buf_4
XFILLER_117_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17053_ _16604_/A _16792_/X _16996_/X vssd1 vssd1 vccd1 vccd1 _20792_/C sky130_fd_sc_hd__a21o_2
X_14265_ _26623_/Q _26719_/Q _14265_/S vssd1 vssd1 vccd1 vccd1 _14265_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16004_ _26076_/Q _25881_/Q _16004_/S vssd1 vssd1 vccd1 vccd1 _16004_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13216_ _13808_/A vssd1 vssd1 vccd1 vccd1 _13955_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14196_ _16711_/A vssd1 vssd1 vccd1 vccd1 _17966_/A sky130_fd_sc_hd__buf_2
XFILLER_98_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13147_ _14263_/S vssd1 vssd1 vccd1 vccd1 _14252_/S sky130_fd_sc_hd__buf_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _15468_/B vssd1 vssd1 vccd1 vccd1 _15635_/B sky130_fd_sc_hd__buf_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ _17953_/X _17954_/X _17958_/S vssd1 vssd1 vccd1 vccd1 _17955_/X sky130_fd_sc_hd__mux2_1
XFILLER_257_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16906_ _16906_/A _16938_/B vssd1 vssd1 vccd1 vccd1 _16939_/A sky130_fd_sc_hd__nand2_1
XFILLER_239_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17886_ _17807_/Y _17990_/A _17973_/A vssd1 vssd1 vccd1 vccd1 _17886_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_211_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19625_ _27066_/Q _19617_/B input175/X _19624_/X vssd1 vssd1 vccd1 vccd1 _19625_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_20_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16837_ _17669_/A _17992_/A _17658_/A vssd1 vssd1 vccd1 vccd1 _17772_/B sky130_fd_sc_hd__o21ai_4
XFILLER_54_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19556_ _19551_/X _19267_/X _19553_/X _19555_/X vssd1 vssd1 vccd1 vccd1 _25655_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16768_ _25683_/Q vssd1 vssd1 vccd1 vccd1 _22520_/A sky130_fd_sc_hd__buf_2
XFILLER_65_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18507_ _27076_/Q vssd1 vssd1 vccd1 vccd1 _19896_/B sky130_fd_sc_hd__clkbuf_2
X_15719_ _15717_/X _15718_/X _15990_/S vssd1 vssd1 vccd1 vccd1 _15719_/X sky130_fd_sc_hd__mux2_1
XFILLER_280_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19487_ _25630_/Q _19497_/B vssd1 vssd1 vccd1 vccd1 _19487_/X sky130_fd_sc_hd__or2_1
XFILLER_221_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16699_ _16826_/A vssd1 vssd1 vccd1 vccd1 _16951_/A sky130_fd_sc_hd__buf_4
XFILLER_278_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18438_ _18438_/A vssd1 vssd1 vccd1 vccd1 _18439_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18369_ _18369_/A vssd1 vssd1 vccd1 vccd1 _18734_/A sky130_fd_sc_hd__buf_2
XFILLER_187_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20400_ _20448_/A _20400_/B vssd1 vssd1 vccd1 vccd1 _20400_/Y sky130_fd_sc_hd__nand2_1
XFILLER_179_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21380_ _21364_/X _18663_/X _21365_/X _25807_/Q _21322_/X vssd1 vssd1 vccd1 vccd1
+ _21380_/X sky130_fd_sc_hd__a221o_1
XFILLER_147_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20331_ _20359_/A _20353_/B vssd1 vssd1 vccd1 vccd1 _20351_/B sky130_fd_sc_hd__xnor2_1
X_23050_ _23523_/A vssd1 vssd1 vccd1 vccd1 _23050_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20262_ _20300_/C _20262_/B vssd1 vssd1 vccd1 vccd1 _20262_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_143_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22001_ _26113_/Q _20926_/X _22005_/S vssd1 vssd1 vccd1 vccd1 _22002_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20193_ _25744_/Q vssd1 vssd1 vccd1 vccd1 _20677_/A sky130_fd_sc_hd__buf_8
XFILLER_89_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput108 dout1[10] vssd1 vssd1 vccd1 vccd1 input108/X sky130_fd_sc_hd__clkbuf_1
Xinput119 dout1[20] vssd1 vssd1 vccd1 vccd1 input119/X sky130_fd_sc_hd__clkbuf_1
XFILLER_229_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23952_ _26852_/Q _23536_/X _23954_/S vssd1 vssd1 vccd1 vccd1 _23953_/A sky130_fd_sc_hd__mux2_1
X_26740_ _26900_/CLK _26740_/D vssd1 vssd1 vccd1 vccd1 _26740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22903_ _22960_/S vssd1 vssd1 vccd1 vccd1 _22912_/S sky130_fd_sc_hd__buf_2
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26671_ _26671_/CLK _26671_/D vssd1 vssd1 vccd1 vccd1 _26671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23883_ _23883_/A vssd1 vssd1 vccd1 vccd1 _26821_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22834_ _26398_/Q _22663_/X _22840_/S vssd1 vssd1 vccd1 vccd1 _22835_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25622_ _25624_/CLK _25622_/D vssd1 vssd1 vccd1 vccd1 _25622_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25553_ _25553_/CLK _25553_/D vssd1 vssd1 vccd1 vccd1 _25553_/Q sky130_fd_sc_hd__dfxtp_1
X_22765_ _26368_/Q _22669_/X _22767_/S vssd1 vssd1 vccd1 vccd1 _22766_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24504_ _24518_/A _24969_/A vssd1 vssd1 vccd1 vccd1 _24504_/Y sky130_fd_sc_hd__nand2_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21716_ _21654_/C _21654_/D _21715_/Y _21349_/B vssd1 vssd1 vccd1 vccd1 _21718_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_212_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25484_ _26683_/CLK _25484_/D vssd1 vssd1 vccd1 vccd1 _25484_/Q sky130_fd_sc_hd__dfxtp_2
X_22696_ _26344_/Q _22695_/X _22705_/S vssd1 vssd1 vccd1 vccd1 _22697_/A sky130_fd_sc_hd__mux2_1
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24435_ _27017_/Q _24421_/X _24434_/Y _24415_/X vssd1 vssd1 vccd1 vccd1 _27017_/D
+ sky130_fd_sc_hd__o211a_1
X_27223_ _27228_/CLK _27223_/D vssd1 vssd1 vccd1 vccd1 _27223_/Q sky130_fd_sc_hd__dfxtp_1
X_21647_ _21647_/A vssd1 vssd1 vccd1 vccd1 _21647_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27154_ _27154_/CLK _27154_/D vssd1 vssd1 vccd1 vccd1 _27154_/Q sky130_fd_sc_hd__dfxtp_2
X_24366_ _14407_/X _21876_/X _24370_/S vssd1 vssd1 vccd1 vccd1 _24645_/B sky130_fd_sc_hd__mux2_4
X_21578_ _21544_/X _21577_/X _21537_/X vssd1 vssd1 vccd1 vccd1 _21578_/Y sky130_fd_sc_hd__o21ai_1
X_26105_ _27275_/CLK _26105_/D vssd1 vssd1 vccd1 vccd1 _26105_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_181_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23317_ _23317_/A vssd1 vssd1 vccd1 vccd1 _26598_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20529_ _23715_/A vssd1 vssd1 vccd1 vccd1 _20529_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27085_ _27087_/CLK _27085_/D vssd1 vssd1 vccd1 vccd1 _27085_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_125_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24297_ _26989_/Q _24295_/B _24296_/Y vssd1 vssd1 vccd1 vccd1 _26989_/D sky130_fd_sc_hd__o21a_1
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26036_ _26595_/CLK _26036_/D vssd1 vssd1 vccd1 vccd1 _26036_/Q sky130_fd_sc_hd__dfxtp_1
X_14050_ _14060_/A vssd1 vssd1 vccd1 vccd1 _14544_/S sky130_fd_sc_hd__buf_2
X_23248_ _23248_/A vssd1 vssd1 vccd1 vccd1 _26567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13001_ _13001_/A _25588_/Q vssd1 vssd1 vccd1 vccd1 _13015_/A sky130_fd_sc_hd__and2_1
XFILLER_106_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23179_ _26537_/Q _23092_/X _23183_/S vssd1 vssd1 vccd1 vccd1 _23180_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17740_ _18119_/A _17750_/A _17740_/C vssd1 vssd1 vccd1 vccd1 _18120_/C sky130_fd_sc_hd__and3b_1
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14952_ _14950_/X _14951_/X _14952_/S vssd1 vssd1 vccd1 vccd1 _14952_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26938_ _26938_/CLK _26938_/D vssd1 vssd1 vccd1 vccd1 _26938_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13903_ _25592_/Q vssd1 vssd1 vccd1 vccd1 _19828_/A sky130_fd_sc_hd__buf_8
XFILLER_36_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17671_ _18010_/C vssd1 vssd1 vccd1 vccd1 _17671_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_236_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14883_ _12705_/A _14874_/X _14882_/X _17195_/A vssd1 vssd1 vccd1 vccd1 _14883_/X
+ sky130_fd_sc_hd__a211o_1
X_26869_ _27258_/CLK _26869_/D vssd1 vssd1 vccd1 vccd1 _26869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19410_ _18912_/A _19408_/Y _18998_/X vssd1 vssd1 vccd1 vccd1 _19410_/X sky130_fd_sc_hd__o21a_1
XFILLER_29_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16622_ _17835_/C vssd1 vssd1 vccd1 vccd1 _18978_/A sky130_fd_sc_hd__buf_4
X_13834_ _13834_/A vssd1 vssd1 vccd1 vccd1 _15205_/A sky130_fd_sc_hd__buf_2
XFILLER_35_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_205 _14662_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_216 _20120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_227 _16012_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19341_ _19341_/A _19472_/B vssd1 vssd1 vccd1 vccd1 _19341_/Y sky130_fd_sc_hd__nor2_1
X_13765_ _13762_/X _13763_/X _13764_/X _13359_/X vssd1 vssd1 vccd1 vccd1 _13765_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_238 _16636_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16553_ _19452_/A _16553_/B vssd1 vssd1 vccd1 vccd1 _25166_/A sky130_fd_sc_hd__xor2_4
XFILLER_44_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_249 _16792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15504_ _13347_/A _15502_/X _15503_/X _13305_/A vssd1 vssd1 vccd1 vccd1 _15504_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_188_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19272_ _19392_/A _19277_/A vssd1 vssd1 vccd1 vccd1 _19272_/Y sky130_fd_sc_hd__nor2_1
X_12716_ _15285_/A vssd1 vssd1 vccd1 vccd1 _14881_/A sky130_fd_sc_hd__clkbuf_4
X_13696_ _15063_/A _25837_/Q _26037_/Q _16050_/B _13051_/A vssd1 vssd1 vccd1 vccd1
+ _13696_/X sky130_fd_sc_hd__a221o_1
XFILLER_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16484_ _16484_/A vssd1 vssd1 vccd1 vccd1 _17697_/B sky130_fd_sc_hd__buf_8
XFILLER_203_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18223_ _18968_/A _18223_/B vssd1 vssd1 vccd1 vccd1 _18223_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15435_ _25744_/Q _20194_/A _16204_/S vssd1 vssd1 vccd1 vccd1 _15438_/B sky130_fd_sc_hd__mux2_2
XFILLER_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18154_ _18154_/A vssd1 vssd1 vccd1 vccd1 _18806_/A sky130_fd_sc_hd__buf_2
XFILLER_175_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15366_ _25889_/Q _16310_/B vssd1 vssd1 vccd1 vccd1 _15366_/X sky130_fd_sc_hd__or2_1
XFILLER_156_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17105_ _17210_/A vssd1 vssd1 vccd1 vccd1 _17105_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14317_ _25727_/Q _14317_/B vssd1 vssd1 vccd1 vccd1 _14317_/X sky130_fd_sc_hd__or2_2
X_15297_ _14763_/A _15295_/X _15296_/X vssd1 vssd1 vccd1 vccd1 _15297_/X sky130_fd_sc_hd__o21a_1
X_18085_ _16586_/B _18080_/Y _18084_/X _17990_/A vssd1 vssd1 vccd1 vccd1 _18085_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_14248_ _26911_/Q _14257_/A vssd1 vssd1 vccd1 vccd1 _14248_/X sky130_fd_sc_hd__or2_1
X_17036_ _17035_/X _16919_/B _17032_/X input227/X vssd1 vssd1 vccd1 vccd1 _17036_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_109_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14179_ _26492_/Q _26364_/Q _14518_/S vssd1 vssd1 vccd1 vccd1 _14179_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ _27086_/Q _18751_/X _18752_/X _27184_/Q _18753_/X vssd1 vssd1 vccd1 vccd1
+ _18987_/X sky130_fd_sc_hd__a221o_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _18063_/S vssd1 vssd1 vccd1 vccd1 _18067_/S sky130_fd_sc_hd__buf_2
XFILLER_239_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17869_ _17801_/B _17787_/B _17909_/S vssd1 vssd1 vccd1 vccd1 _17869_/X sky130_fd_sc_hd__mux2_1
XFILLER_254_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19608_ _26061_/Q vssd1 vssd1 vccd1 vccd1 _19617_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20880_ _20880_/A vssd1 vssd1 vccd1 vccd1 _25831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19539_ _19552_/A vssd1 vssd1 vccd1 vccd1 _19549_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_81_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22550_ _22538_/X _22549_/Y _22547_/X vssd1 vssd1 vccd1 vccd1 _26296_/D sky130_fd_sc_hd__a21oi_1
XFILLER_107_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21501_ input53/X input89/X _21553_/S vssd1 vssd1 vccd1 vccd1 _21502_/A sky130_fd_sc_hd__mux2_8
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22481_ _22481_/A vssd1 vssd1 vccd1 vccd1 _26266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24220_ _26963_/Q _24221_/C _26964_/Q vssd1 vssd1 vccd1 vccd1 _24222_/B sky130_fd_sc_hd__a21oi_1
X_21432_ _21430_/X _18876_/X _21431_/X _25811_/Q _21403_/X vssd1 vssd1 vccd1 vccd1
+ _21432_/X sky130_fd_sc_hd__a221o_1
XFILLER_108_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24151_ _26941_/Q _27327_/Q vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__and2b_1
XFILLER_257_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21363_ _23363_/A _21416_/B vssd1 vssd1 vccd1 vccd1 _21363_/X sky130_fd_sc_hd__or2_1
XFILLER_257_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23102_ _23118_/A vssd1 vssd1 vccd1 vccd1 _23115_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_163_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20314_ _19879_/X _20313_/X _19926_/X vssd1 vssd1 vccd1 vccd1 _20317_/B sky130_fd_sc_hd__a21oi_1
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24082_ _24082_/A vssd1 vssd1 vccd1 vccd1 _26909_/D sky130_fd_sc_hd__clkbuf_1
Xinput90 dout0[52] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_1
X_21294_ input76/X input71/X _21327_/S vssd1 vssd1 vccd1 vccd1 _21294_/X sky130_fd_sc_hd__mux2_8
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23033_ _23033_/A vssd1 vssd1 vccd1 vccd1 _26487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20245_ _19649_/A _20242_/Y _20243_/X _20244_/X vssd1 vssd1 vccd1 vccd1 _20245_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_277_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20176_ _19796_/X _20174_/X _20175_/Y _19890_/X vssd1 vssd1 vccd1 vccd1 _20176_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_77_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24984_ _24629_/A _24902_/A _24966_/X vssd1 vssd1 vccd1 vccd1 _24984_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_276_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26723_ _26916_/CLK _26723_/D vssd1 vssd1 vccd1 vccd1 _26723_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23935_ _26844_/Q _23508_/X _23943_/S vssd1 vssd1 vccd1 vccd1 _23936_/A sky130_fd_sc_hd__mux2_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26654_ _26813_/CLK _26654_/D vssd1 vssd1 vccd1 vccd1 _26654_/Q sky130_fd_sc_hd__dfxtp_1
X_23866_ _23866_/A vssd1 vssd1 vccd1 vccd1 _26813_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_260_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25605_ _25607_/CLK _25605_/D vssd1 vssd1 vccd1 vccd1 _25605_/Q sky130_fd_sc_hd__dfxtp_4
X_22817_ _22817_/A _22817_/B _22817_/C vssd1 vssd1 vccd1 vccd1 _25393_/B sky130_fd_sc_hd__or3_4
XFILLER_60_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23797_ _23696_/X _26783_/Q _23799_/S vssd1 vssd1 vccd1 vccd1 _23798_/A sky130_fd_sc_hd__mux2_1
X_26585_ _27156_/CLK _26585_/D vssd1 vssd1 vccd1 vccd1 _26585_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_60_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13550_ _15526_/S _19912_/A _13549_/X vssd1 vssd1 vccd1 vccd1 _17821_/B sky130_fd_sc_hd__a21boi_2
XFILLER_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22748_ _26360_/Q _22640_/X _22756_/S vssd1 vssd1 vccd1 vccd1 _22749_/A sky130_fd_sc_hd__mux2_1
X_25536_ _25545_/CLK _25536_/D vssd1 vssd1 vccd1 vccd1 _25536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13481_ _25581_/Q vssd1 vssd1 vccd1 vccd1 _14468_/A sky130_fd_sc_hd__clkbuf_2
X_25467_ _25467_/A vssd1 vssd1 vccd1 vccd1 _27327_/D sky130_fd_sc_hd__clkbuf_1
X_22679_ _23722_/A vssd1 vssd1 vccd1 vccd1 _22679_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_186_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15220_ _14754_/A _15218_/X _15219_/X _14803_/A vssd1 vssd1 vccd1 vccd1 _15220_/X
+ sky130_fd_sc_hd__a211o_1
X_24418_ _24392_/X _25607_/Q _24417_/X vssd1 vssd1 vccd1 vccd1 _24932_/A sky130_fd_sc_hd__o21ai_4
X_27206_ _27230_/CLK _27206_/D vssd1 vssd1 vccd1 vccd1 _27206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25398_ _23690_/X _27296_/Q _25404_/S vssd1 vssd1 vccd1 vccd1 _25399_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15151_ _25821_/Q _16235_/S _16401_/S _15150_/X vssd1 vssd1 vccd1 vccd1 _15151_/X
+ sky130_fd_sc_hd__o211a_1
X_27137_ _27137_/CLK _27137_/D vssd1 vssd1 vccd1 vccd1 _27137_/Q sky130_fd_sc_hd__dfxtp_2
X_24349_ _24542_/A _24542_/B vssd1 vssd1 vccd1 vccd1 _25206_/C sky130_fd_sc_hd__or2b_1
XFILLER_126_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14102_ _27268_/Q _26461_/Q _14257_/A vssd1 vssd1 vccd1 vccd1 _14102_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27068_ _27133_/CLK _27068_/D vssd1 vssd1 vccd1 vccd1 _27068_/Q sky130_fd_sc_hd__dfxtp_2
X_15082_ _25750_/Q vssd1 vssd1 vccd1 vccd1 _20692_/A sky130_fd_sc_hd__inv_4
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14033_ input128/X input164/X _14033_/S vssd1 vssd1 vccd1 vccd1 _14033_/X sky130_fd_sc_hd__mux2_8
X_26019_ _26611_/CLK _26019_/D vssd1 vssd1 vccd1 vccd1 _26019_/Q sky130_fd_sc_hd__dfxtp_1
X_18910_ _18910_/A vssd1 vssd1 vccd1 vccd1 _18912_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19890_ _19926_/A vssd1 vssd1 vccd1 vccd1 _19890_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_268_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18841_ _18927_/A vssd1 vssd1 vccd1 vccd1 _18841_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18772_ _18742_/X _18745_/X _18771_/X vssd1 vssd1 vccd1 vccd1 _18772_/X sky130_fd_sc_hd__a21o_4
XFILLER_283_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15984_ _25704_/Q _15984_/B vssd1 vssd1 vccd1 vccd1 _15984_/X sky130_fd_sc_hd__or2_1
XFILLER_209_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17723_ _17762_/C _17730_/A vssd1 vssd1 vccd1 vccd1 _18440_/A sky130_fd_sc_hd__and2b_1
XFILLER_282_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14935_ _16556_/A vssd1 vssd1 vccd1 vccd1 _16461_/A sky130_fd_sc_hd__inv_2
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17654_ _25933_/Q _17544_/X _17653_/X vssd1 vssd1 vccd1 vccd1 _17654_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14866_ _12775_/A _26905_/Q _26777_/Q _14846_/B _14688_/A vssd1 vssd1 vccd1 vccd1
+ _14866_/X sky130_fd_sc_hd__a221o_1
XFILLER_235_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16605_ _19156_/A _19156_/B _19158_/S vssd1 vssd1 vccd1 vccd1 _19187_/A sky130_fd_sc_hd__a21oi_4
XFILLER_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13817_ _13346_/A _13815_/X _13816_/X _13366_/A vssd1 vssd1 vccd1 vccd1 _13818_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_223_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17585_ _25915_/Q _17568_/X _14032_/B _17577_/X vssd1 vssd1 vccd1 vccd1 _17585_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14797_ _14795_/X _14796_/X _16524_/A vssd1 vssd1 vccd1 vccd1 _14797_/X sky130_fd_sc_hd__mux2_1
XFILLER_251_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_69_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26465_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_250_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19324_ _18682_/A _18321_/B _18312_/Y _18342_/A vssd1 vssd1 vccd1 vccd1 _19324_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_16536_ _14755_/X _16534_/X _16535_/X _14804_/X vssd1 vssd1 vccd1 vccd1 _16536_/X
+ sky130_fd_sc_hd__a211o_1
X_13748_ _13748_/A _13748_/B vssd1 vssd1 vccd1 vccd1 _13748_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19255_ _25622_/Q _19153_/X _19254_/X _19185_/X vssd1 vssd1 vccd1 vccd1 _25622_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16467_ _16467_/A vssd1 vssd1 vccd1 vccd1 _16498_/S sky130_fd_sc_hd__clkbuf_2
X_13679_ _12738_/D _26105_/Q _26006_/Q _16013_/S _14768_/A vssd1 vssd1 vccd1 vccd1
+ _13679_/X sky130_fd_sc_hd__a221o_1
X_18206_ _17892_/X _17873_/X _18209_/S vssd1 vssd1 vccd1 vccd1 _18206_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15418_ _15318_/X _15415_/X _15417_/X _15313_/X vssd1 vssd1 vccd1 vccd1 _15418_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19186_ _25620_/Q _19153_/X _19184_/X _19185_/X vssd1 vssd1 vccd1 vccd1 _25620_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16398_ _16394_/X _16397_/X _16398_/S vssd1 vssd1 vccd1 vccd1 _16398_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18137_ _18945_/A vssd1 vssd1 vccd1 vccd1 _18910_/A sky130_fd_sc_hd__clkbuf_2
X_15349_ _25618_/Q _14597_/A _15348_/X _14618_/A vssd1 vssd1 vccd1 vccd1 _23574_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_89_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18068_ _18066_/X _18067_/X _18071_/S vssd1 vssd1 vccd1 vccd1 _18068_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17019_ _17015_/X _16850_/B _17017_/X input246/X vssd1 vssd1 vccd1 vccd1 _17019_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_259_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20030_ _25674_/Q _20030_/B vssd1 vssd1 vccd1 vccd1 _20098_/C sky130_fd_sc_hd__and2_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21981_ _26104_/Q _20897_/X _21983_/S vssd1 vssd1 vccd1 vccd1 _21982_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23720_ _23718_/X _26758_/Q _23732_/S vssd1 vssd1 vccd1 vccd1 _23721_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20932_ _23747_/A vssd1 vssd1 vccd1 vccd1 _20932_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_254_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23651_ _23651_/A vssd1 vssd1 vccd1 vccd1 _26732_/D sky130_fd_sc_hd__clkbuf_1
X_20863_ _20863_/A vssd1 vssd1 vccd1 vccd1 _25827_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22602_ _26316_/Q _22604_/B vssd1 vssd1 vccd1 vccd1 _22602_/Y sky130_fd_sc_hd__nand2_1
X_26370_ _27277_/CLK _26370_/D vssd1 vssd1 vccd1 vccd1 _26370_/Q sky130_fd_sc_hd__dfxtp_1
X_23582_ _26706_/Q _23581_/X _23588_/S vssd1 vssd1 vccd1 vccd1 _23583_/A sky130_fd_sc_hd__mux2_1
X_20794_ _22472_/B _20973_/B _20794_/C vssd1 vssd1 vccd1 vccd1 _20795_/A sky130_fd_sc_hd__and3_1
X_25321_ _25321_/A _25321_/B vssd1 vssd1 vccd1 vccd1 _25378_/A sky130_fd_sc_hd__nor2_8
XFILLER_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22533_ _22533_/A _22533_/B vssd1 vssd1 vccd1 vccd1 _22534_/A sky130_fd_sc_hd__and2_1
XFILLER_23_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25252_ _23684_/X _27231_/Q _25260_/S vssd1 vssd1 vccd1 vccd1 _25253_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22464_ _26209_/Q _22459_/X _22463_/X _22455_/X vssd1 vssd1 vccd1 vccd1 _26257_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24203_ _26958_/Q _26957_/Q _24203_/C vssd1 vssd1 vccd1 vccd1 _24205_/B sky130_fd_sc_hd__and3_1
XFILLER_182_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21415_ _21545_/A vssd1 vssd1 vccd1 vccd1 _21415_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25183_ _25206_/B _25206_/C _25206_/D vssd1 vssd1 vccd1 vccd1 _25218_/B sky130_fd_sc_hd__nor3_1
X_22395_ _22395_/A _22395_/B vssd1 vssd1 vccd1 vccd1 _22395_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24134_ _26933_/Q _23590_/X _24142_/S vssd1 vssd1 vccd1 vccd1 _24135_/A sky130_fd_sc_hd__mux2_1
X_21346_ _21346_/A vssd1 vssd1 vccd1 vccd1 _21346_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24065_ _24065_/A vssd1 vssd1 vccd1 vccd1 _26902_/D sky130_fd_sc_hd__clkbuf_1
X_21277_ _21277_/A vssd1 vssd1 vccd1 vccd1 _21278_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23016_ _23016_/A vssd1 vssd1 vccd1 vccd1 _26479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20228_ _20141_/B _19148_/X _19911_/X _20227_/Y vssd1 vssd1 vccd1 vccd1 _20228_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_89_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20159_ _20159_/A _20158_/Y vssd1 vssd1 vccd1 vccd1 _20160_/B sky130_fd_sc_hd__or2b_1
XFILLER_249_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _12981_/A _14610_/B vssd1 vssd1 vccd1 vccd1 _13577_/A sky130_fd_sc_hd__nand2_2
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24967_ _24611_/A _24941_/X _24966_/X vssd1 vssd1 vccd1 vccd1 _24967_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26706_ _27285_/CLK _26706_/D vssd1 vssd1 vccd1 vccd1 _26706_/Q sky130_fd_sc_hd__dfxtp_1
X_14720_ _25595_/Q _18059_/A _14719_/Y vssd1 vssd1 vccd1 vccd1 _14831_/A sky130_fd_sc_hd__o21ai_4
XFILLER_217_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23918_ _23766_/X _26837_/Q _23926_/S vssd1 vssd1 vccd1 vccd1 _23919_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24898_ _24896_/Y _24897_/X _21242_/X vssd1 vssd1 vccd1 vccd1 _27132_/D sky130_fd_sc_hd__a21oi_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26637_ _26797_/CLK _26637_/D vssd1 vssd1 vccd1 vccd1 _26637_/Q sky130_fd_sc_hd__dfxtp_1
X_14651_ _16499_/S _14638_/X _14646_/X _14650_/X vssd1 vssd1 vccd1 vccd1 _14651_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23849_ _23849_/A vssd1 vssd1 vccd1 vccd1 _26806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _14330_/A vssd1 vssd1 vccd1 vccd1 _14254_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_214_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _25541_/Q _25542_/Q _17370_/C vssd1 vssd1 vccd1 vccd1 _17372_/B sky130_fd_sc_hd__and3_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14582_ _16122_/S vssd1 vssd1 vccd1 vccd1 _16204_/S sky130_fd_sc_hd__buf_2
X_26568_ _27282_/CLK _26568_/D vssd1 vssd1 vccd1 vccd1 _26568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16321_ _16317_/X _16320_/X _16398_/S vssd1 vssd1 vccd1 vccd1 _16321_/X sky130_fd_sc_hd__mux2_1
X_13533_ _16004_/S vssd1 vssd1 vccd1 vccd1 _13534_/S sky130_fd_sc_hd__buf_2
X_25519_ _27022_/CLK _25519_/D vssd1 vssd1 vccd1 vccd1 _25519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26499_ _26531_/CLK _26499_/D vssd1 vssd1 vccd1 vccd1 _26499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19040_ _18723_/X _19036_/X _19039_/X _18884_/X vssd1 vssd1 vccd1 vccd1 _19041_/B
+ sky130_fd_sc_hd__a22o_1
X_13464_ _13464_/A vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__buf_2
XFILLER_146_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16252_ _25820_/Q _27254_/Q _16255_/S vssd1 vssd1 vccd1 vccd1 _16252_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15203_ _26544_/Q _26152_/Q _16436_/S vssd1 vssd1 vccd1 vccd1 _15203_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13395_ _14031_/A _13395_/B vssd1 vssd1 vccd1 vccd1 _13395_/Y sky130_fd_sc_hd__nor2_1
X_16183_ _16181_/X _16182_/X _16183_/S vssd1 vssd1 vccd1 vccd1 _16183_/X sky130_fd_sc_hd__mux2_1
X_15134_ _15134_/A _16292_/B vssd1 vssd1 vccd1 vccd1 _15134_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_187_wb_clk_i _26681_/CLK vssd1 vssd1 vccd1 vccd1 _27291_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_116_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26992_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19942_ _19978_/A _19978_/B vssd1 vssd1 vccd1 vccd1 _19951_/A sky130_fd_sc_hd__or2_1
X_15065_ _15065_/A vssd1 vssd1 vccd1 vccd1 _15065_/X sky130_fd_sc_hd__buf_2
X_14016_ _13112_/A _14003_/X _14007_/X _14015_/X _13876_/X vssd1 vssd1 vccd1 vccd1
+ _14016_/X sky130_fd_sc_hd__a311o_1
XFILLER_141_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19873_ _22130_/A vssd1 vssd1 vccd1 vccd1 _21718_/A sky130_fd_sc_hd__buf_6
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18824_ _27050_/Q _18811_/X _18819_/X _18822_/X _18823_/X vssd1 vssd1 vccd1 vccd1
+ _18824_/X sky130_fd_sc_hd__o221a_2
XFILLER_68_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18755_ _27113_/Q _18748_/X _18750_/X _18754_/X vssd1 vssd1 vccd1 vccd1 _18755_/X
+ sky130_fd_sc_hd__o22a_2
XTAP_5480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15967_ _13410_/X _15964_/X _15966_/X _13863_/X vssd1 vssd1 vccd1 vccd1 _15967_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput280 versionID[0] vssd1 vssd1 vccd1 vccd1 input280/X sky130_fd_sc_hd__clkbuf_2
XFILLER_209_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17706_ _17706_/A _17706_/B vssd1 vssd1 vccd1 vccd1 _24342_/A sky130_fd_sc_hd__and2_1
XFILLER_36_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14918_ _14890_/A _25787_/Q _15005_/S _26873_/Q _14917_/X vssd1 vssd1 vccd1 vccd1
+ _14918_/X sky130_fd_sc_hd__o221a_1
XFILLER_224_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18686_ _18686_/A _18686_/B vssd1 vssd1 vccd1 vccd1 _18686_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15898_ _14153_/X _25771_/Q _14103_/X _26857_/Q _14264_/S vssd1 vssd1 vccd1 vccd1
+ _15898_/X sky130_fd_sc_hd__o221a_1
XFILLER_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17637_ _12721_/A _17635_/X _17604_/X _17636_/Y vssd1 vssd1 vccd1 vccd1 _17638_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_36_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14849_ _26873_/Q _25787_/Q _14960_/B vssd1 vssd1 vccd1 vccd1 _14849_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17568_ _17597_/A vssd1 vssd1 vccd1 vccd1 _17568_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19307_ _25527_/Q _18810_/X _19304_/X _19306_/X _18832_/X vssd1 vssd1 vccd1 vccd1
+ _19307_/X sky130_fd_sc_hd__o221a_1
XFILLER_204_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16519_ _16513_/X _25860_/Q _26060_/Q _16526_/S _14773_/X vssd1 vssd1 vccd1 vccd1
+ _16519_/X sky130_fd_sc_hd__a221o_1
X_17499_ _17475_/X _17483_/Y _21221_/A _24454_/A vssd1 vssd1 vccd1 vccd1 _17514_/C
+ sky130_fd_sc_hd__o31a_2
XFILLER_149_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19238_ _19276_/B _19238_/B vssd1 vssd1 vccd1 vccd1 _19576_/D sky130_fd_sc_hd__nand2_1
XFILLER_219_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19169_ _26963_/Q _18826_/X _18827_/X _26995_/Q vssd1 vssd1 vccd1 vccd1 _19169_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21200_ _17020_/A _16674_/A _16679_/B _21199_/X vssd1 vssd1 vccd1 vccd1 _21309_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_145_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22180_ _26177_/Q _22171_/X _22179_/X input276/X _22172_/X vssd1 vssd1 vccd1 vccd1
+ _22180_/X sky130_fd_sc_hd__a221o_1
XFILLER_219_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21131_ _21167_/A vssd1 vssd1 vccd1 vccd1 _21131_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21062_ _21062_/A vssd1 vssd1 vccd1 vccd1 _25899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20013_ _20039_/A _20039_/B vssd1 vssd1 vccd1 vccd1 _20080_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25870_ _27265_/CLK _25870_/D vssd1 vssd1 vccd1 vccd1 _25870_/Q sky130_fd_sc_hd__dfxtp_1
X_24821_ _24877_/A vssd1 vssd1 vccd1 vccd1 _24837_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_246_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21964_ _26096_/Q _20866_/X _21972_/S vssd1 vssd1 vccd1 vccd1 _21965_/A sky130_fd_sc_hd__mux2_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24752_ _27094_/Q _24744_/X _25143_/A _24740_/X vssd1 vssd1 vccd1 vccd1 _24753_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_54_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20915_ _20915_/A vssd1 vssd1 vccd1 vccd1 _25842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23703_ _23786_/S vssd1 vssd1 vccd1 vccd1 _23716_/S sky130_fd_sc_hd__buf_2
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24683_ _19957_/B _24680_/X _24682_/Y _24676_/X vssd1 vssd1 vccd1 vccd1 _24684_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_21895_ _21895_/A vssd1 vssd1 vccd1 vccd1 _26065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23634_ _26725_/Q _23539_/X _23634_/S vssd1 vssd1 vccd1 vccd1 _23635_/A sky130_fd_sc_hd__mux2_1
X_26422_ _27326_/CLK _26422_/D vssd1 vssd1 vccd1 vccd1 _26422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20846_ _25819_/Q vssd1 vssd1 vccd1 vccd1 _20847_/A sky130_fd_sc_hd__clkbuf_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23565_ _23565_/A vssd1 vssd1 vccd1 vccd1 _23565_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26353_ _26677_/CLK _26353_/D vssd1 vssd1 vccd1 vccd1 _26353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20777_ _20601_/X _25784_/Q _20783_/S vssd1 vssd1 vccd1 vccd1 _20778_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22516_ _22516_/A _22524_/B vssd1 vssd1 vccd1 vccd1 _22517_/A sky130_fd_sc_hd__and2_1
X_25304_ _23763_/X _27255_/Q _25304_/S vssd1 vssd1 vccd1 vccd1 _25305_/A sky130_fd_sc_hd__mux2_1
X_26284_ _26286_/CLK _26284_/D vssd1 vssd1 vccd1 vccd1 _26284_/Q sky130_fd_sc_hd__dfxtp_1
X_23496_ _26678_/Q _23121_/X _23502_/S vssd1 vssd1 vccd1 vccd1 _23497_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22447_ _22460_/A vssd1 vssd1 vccd1 vccd1 _22457_/B sky130_fd_sc_hd__clkbuf_1
X_25235_ _19614_/C _25209_/X _25179_/A vssd1 vssd1 vccd1 vccd1 _25235_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25166_ _25166_/A vssd1 vssd1 vccd1 vccd1 _25166_/Y sky130_fd_sc_hd__inv_2
X_13180_ _13180_/A vssd1 vssd1 vccd1 vccd1 _14566_/A sky130_fd_sc_hd__clkbuf_2
X_22378_ _22378_/A vssd1 vssd1 vccd1 vccd1 _26236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24117_ _24117_/A vssd1 vssd1 vccd1 vccd1 _26925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21329_ _21326_/Y _21328_/Y _21297_/X vssd1 vssd1 vccd1 vccd1 _21329_/Y sky130_fd_sc_hd__a21oi_4
X_25097_ _25124_/A vssd1 vssd1 vccd1 vccd1 _25097_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24048_ _26895_/Q _23571_/X _24048_/S vssd1 vssd1 vccd1 vccd1 _24049_/A sky130_fd_sc_hd__mux2_1
XFILLER_278_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_132_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16870_ _16893_/A _16870_/B vssd1 vssd1 vccd1 vccd1 _16871_/A sky130_fd_sc_hd__and2_1
XFILLER_104_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15821_ _26666_/Q _15474_/S _15820_/X _13050_/A vssd1 vssd1 vccd1 vccd1 _15821_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25999_ _26240_/CLK _25999_/D vssd1 vssd1 vccd1 vccd1 _25999_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18540_ _18593_/B _18540_/B vssd1 vssd1 vccd1 vccd1 _19572_/C sky130_fd_sc_hd__and2b_1
X_15752_ _26635_/Q _26731_/Q _15931_/S vssd1 vssd1 vccd1 vccd1 _15753_/B sky130_fd_sc_hd__mux2_1
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12964_ _12964_/A vssd1 vssd1 vccd1 vccd1 _13933_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_70 _20677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_81 _23706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_92 _24871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14703_ _12760_/B _14701_/X _14702_/X vssd1 vssd1 vccd1 vccd1 _14704_/B sky130_fd_sc_hd__o21ai_1
XFILLER_261_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18471_ _18437_/X _18442_/X _18470_/X vssd1 vssd1 vccd1 vccd1 _18471_/X sky130_fd_sc_hd__a21o_4
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _15318_/A _15680_/X _15682_/X _15313_/A vssd1 vssd1 vccd1 vccd1 _15683_/X
+ sky130_fd_sc_hd__o211a_1
X_12895_ _13741_/S vssd1 vssd1 vccd1 vccd1 _14033_/S sky130_fd_sc_hd__buf_2
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _25558_/Q _17420_/B _17421_/Y vssd1 vssd1 vccd1 vccd1 _25558_/D sky130_fd_sc_hd__o21a_1
XFILLER_205_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14634_ _16242_/S vssd1 vssd1 vccd1 vccd1 _15014_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_61_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _25537_/Q _17353_/B vssd1 vssd1 vccd1 vccd1 _17360_/C sky130_fd_sc_hd__and2_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14565_ _16586_/B _16580_/A _14562_/X _14564_/X vssd1 vssd1 vccd1 vccd1 _16706_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16304_ _16378_/S _16301_/X _16303_/X _15040_/X vssd1 vssd1 vccd1 vccd1 _16304_/X
+ sky130_fd_sc_hd__a211o_1
X_13516_ _14365_/S vssd1 vssd1 vccd1 vccd1 _15292_/A sky130_fd_sc_hd__buf_6
XFILLER_202_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17284_ _25516_/Q _17284_/B vssd1 vssd1 vccd1 vccd1 _17293_/C sky130_fd_sc_hd__and2_1
XFILLER_147_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14496_ _13084_/A _26392_/Q _15980_/S _26908_/Q _13862_/A vssd1 vssd1 vccd1 vccd1
+ _14496_/X sky130_fd_sc_hd__o221a_1
XFILLER_186_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19023_ _27119_/Q _18812_/X _19021_/X _19022_/X vssd1 vssd1 vccd1 vccd1 _19023_/X
+ sky130_fd_sc_hd__o22a_2
X_16235_ _26867_/Q _25781_/Q _16235_/S vssd1 vssd1 vccd1 vccd1 _16235_/X sky130_fd_sc_hd__mux2_1
X_13447_ _13445_/X _13446_/X _13698_/A vssd1 vssd1 vccd1 vccd1 _13447_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13378_ _25735_/Q _15615_/S vssd1 vssd1 vccd1 vccd1 _13378_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16166_ _16160_/X _16162_/X _14708_/A _16165_/X vssd1 vssd1 vccd1 vccd1 _16167_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15117_ _16439_/A _15117_/B _15117_/C vssd1 vssd1 vccd1 vccd1 _15117_/X sky130_fd_sc_hd__or3_1
XFILLER_170_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16097_ _15394_/A _16094_/X _16096_/X _13291_/X vssd1 vssd1 vccd1 vccd1 _16097_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_269_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15048_ _15048_/A vssd1 vssd1 vccd1 vccd1 _15048_/X sky130_fd_sc_hd__buf_2
X_19925_ _19951_/B _19925_/B vssd1 vssd1 vccd1 vccd1 _19925_/Y sky130_fd_sc_hd__nand2_1
XFILLER_284_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19856_ _17444_/A _19829_/A _19803_/B _19676_/A _12721_/A vssd1 vssd1 vccd1 vccd1
+ _19856_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_69_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18807_ _18807_/A vssd1 vssd1 vccd1 vccd1 _18807_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19787_ _19787_/A vssd1 vssd1 vccd1 vccd1 _20323_/B sky130_fd_sc_hd__clkbuf_2
X_16999_ _22489_/A _16996_/X _16990_/A _16732_/X vssd1 vssd1 vccd1 vccd1 _16999_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_271_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_84_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26657_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18738_ _18738_/A vssd1 vssd1 vccd1 vccd1 _18738_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_243_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26671_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18669_ _18340_/A _16735_/X _18648_/Y _18668_/X vssd1 vssd1 vccd1 vccd1 _18669_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20700_ _26290_/Q _20687_/B _20699_/X _20697_/X vssd1 vssd1 vccd1 vccd1 _25753_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21680_ _21680_/A vssd1 vssd1 vccd1 vccd1 _25979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20631_ _20644_/A vssd1 vssd1 vccd1 vccd1 _20631_/X sky130_fd_sc_hd__buf_2
XFILLER_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23350_ _23350_/A vssd1 vssd1 vccd1 vccd1 _26613_/D sky130_fd_sc_hd__clkbuf_1
X_20562_ _23565_/A vssd1 vssd1 vccd1 vccd1 _23741_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_220_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22301_ _22317_/A vssd1 vssd1 vccd1 vccd1 _22301_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23281_ _26583_/Q _23136_/X _23281_/S vssd1 vssd1 vccd1 vccd1 _23282_/A sky130_fd_sc_hd__mux2_1
X_20493_ _20484_/X _25692_/Q _20509_/S vssd1 vssd1 vccd1 vccd1 _20494_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25020_ _22476_/A _25015_/X _25004_/X _18230_/B _25005_/X vssd1 vssd1 vccd1 vccd1
+ _25020_/X sky130_fd_sc_hd__a221o_1
XFILLER_118_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22232_ _17094_/B _22113_/X _22231_/X _22217_/X vssd1 vssd1 vccd1 vccd1 _26192_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_192_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22163_ _26172_/Q _22154_/X _22160_/X input271/X _22155_/X vssd1 vssd1 vccd1 vccd1
+ _22163_/X sky130_fd_sc_hd__a221o_1
XFILLER_1_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21114_ _25912_/Q _21112_/X _21113_/X input11/X vssd1 vssd1 vccd1 vccd1 _21115_/B
+ sky130_fd_sc_hd__o22a_1
X_26971_ _26974_/CLK _26971_/D vssd1 vssd1 vccd1 vccd1 _26971_/Q sky130_fd_sc_hd__dfxtp_1
X_22094_ _22094_/A vssd1 vssd1 vccd1 vccd1 _26154_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21045_ _21045_/A vssd1 vssd1 vccd1 vccd1 _25891_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25922_ _27213_/CLK _25922_/D vssd1 vssd1 vccd1 vccd1 _25922_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_120_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25853_ _27329_/A _25853_/D vssd1 vssd1 vccd1 vccd1 _25853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24804_ _20637_/A _24789_/X _24664_/Y _24791_/X vssd1 vssd1 vccd1 vccd1 _24804_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_262_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25784_ _27257_/CLK _25784_/D vssd1 vssd1 vccd1 vccd1 _25784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_274_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22996_ _22996_/A vssd1 vssd1 vccd1 vccd1 _26470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24735_ hold1/A vssd1 vssd1 vccd1 vccd1 _24736_/B sky130_fd_sc_hd__clkinv_2
XFILLER_28_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21947_ _20596_/X _26089_/Q _21955_/S vssd1 vssd1 vccd1 vccd1 _21948_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12680_ _13001_/A vssd1 vssd1 vccd1 vccd1 _13185_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21878_ _21878_/A vssd1 vssd1 vccd1 vccd1 _21878_/X sky130_fd_sc_hd__buf_6
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24666_ _24678_/A _24666_/B vssd1 vssd1 vccd1 vccd1 _27074_/D sky130_fd_sc_hd__nor2_1
XFILLER_215_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26405_ _26468_/CLK _26405_/D vssd1 vssd1 vccd1 vccd1 _26405_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23617_ _26717_/Q _23514_/X _23623_/S vssd1 vssd1 vccd1 vccd1 _23618_/A sky130_fd_sc_hd__mux2_1
X_20829_ _20829_/A vssd1 vssd1 vccd1 vccd1 _25810_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24597_ _24610_/A vssd1 vssd1 vccd1 vccd1 _24608_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26336_ _27275_/CLK _26336_/D vssd1 vssd1 vccd1 vccd1 _26336_/Q sky130_fd_sc_hd__dfxtp_4
X_14350_ _26098_/Q _25999_/Q _14351_/S vssd1 vssd1 vccd1 vccd1 _14350_/X sky130_fd_sc_hd__mux2_1
XFILLER_211_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23548_ _23548_/A vssd1 vssd1 vccd1 vccd1 _26695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13301_ _15321_/A _27274_/Q _26467_/Q _16267_/S _13281_/A vssd1 vssd1 vccd1 vccd1
+ _13301_/X sky130_fd_sc_hd__a221o_1
XFILLER_11_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14281_ _13009_/A _23520_/A _14280_/X vssd1 vssd1 vccd1 vccd1 _16820_/B sky130_fd_sc_hd__o21ai_4
XFILLER_156_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23479_ _23479_/A vssd1 vssd1 vccd1 vccd1 _26670_/D sky130_fd_sc_hd__clkbuf_1
X_26267_ _26271_/CLK _26267_/D vssd1 vssd1 vccd1 vccd1 _26267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16020_ _27307_/Q _26564_/Q _16020_/S vssd1 vssd1 vccd1 vccd1 _16020_/X sky130_fd_sc_hd__mux2_1
X_13232_ _13821_/A vssd1 vssd1 vccd1 vccd1 _15924_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25218_ _25218_/A _25218_/B vssd1 vssd1 vccd1 vccd1 _25219_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26198_ _26250_/CLK _26198_/D vssd1 vssd1 vccd1 vccd1 _26198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13163_ _13163_/A vssd1 vssd1 vccd1 vccd1 _13164_/A sky130_fd_sc_hd__buf_2
X_25149_ _22528_/A _24639_/A _25139_/X _16575_/B _12781_/X vssd1 vssd1 vccd1 vccd1
+ _25149_/X sky130_fd_sc_hd__a221o_1
XFILLER_123_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13094_ _15474_/S vssd1 vssd1 vccd1 vccd1 _15467_/S sky130_fd_sc_hd__buf_2
X_17971_ _17971_/A _17971_/B _17971_/C _17971_/D vssd1 vssd1 vccd1 vccd1 _17971_/X
+ sky130_fd_sc_hd__or4_2
X_19710_ _20115_/A _19666_/X _20091_/A _20628_/A _19673_/B vssd1 vssd1 vccd1 vccd1
+ _19710_/Y sky130_fd_sc_hd__o221ai_2
X_16922_ _16909_/X _16873_/B _16872_/X _16910_/X _16911_/X vssd1 vssd1 vccd1 vccd1
+ _16922_/X sky130_fd_sc_hd__o221a_1
XFILLER_238_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19641_ _24777_/A vssd1 vssd1 vccd1 vccd1 _24848_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_265_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16853_ _16853_/A vssd1 vssd1 vccd1 vccd1 _16983_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_120_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15804_ _26342_/Q _26602_/Q _15805_/S vssd1 vssd1 vccd1 vccd1 _15804_/X sky130_fd_sc_hd__mux2_1
X_19572_ _19572_/A _19572_/B _19572_/C _19572_/D vssd1 vssd1 vccd1 vccd1 _19573_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_219_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16784_ _16834_/A vssd1 vssd1 vccd1 vccd1 _16784_/X sky130_fd_sc_hd__buf_4
XFILLER_219_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13996_ _26786_/Q _26430_/Q _14009_/S vssd1 vssd1 vccd1 vccd1 _13996_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18523_ _17259_/X _18444_/X _18520_/X _18522_/X _18469_/X vssd1 vssd1 vccd1 vccd1
+ _18523_/X sky130_fd_sc_hd__o221a_1
XFILLER_218_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15735_ _27246_/Q _15984_/B vssd1 vssd1 vccd1 vccd1 _15735_/X sky130_fd_sc_hd__or2_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ _12962_/C _12947_/B vssd1 vssd1 vccd1 vccd1 _12948_/C sky130_fd_sc_hd__nor2_1
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18454_ _18454_/A vssd1 vssd1 vccd1 vccd1 _18455_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_179_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15666_ _13267_/X _26892_/Q _26764_/Q _16186_/S _13221_/A vssd1 vssd1 vccd1 vccd1
+ _15666_/X sky130_fd_sc_hd__a221o_1
X_12878_ _21429_/A _12878_/B vssd1 vssd1 vccd1 vccd1 _12878_/Y sky130_fd_sc_hd__nor2_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _17408_/A _17408_/C _17366_/X vssd1 vssd1 vccd1 vccd1 _17405_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_233_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14617_ _14617_/A vssd1 vssd1 vccd1 vccd1 _14618_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18385_ _19769_/A _19374_/B vssd1 vssd1 vccd1 vccd1 _18386_/B sky130_fd_sc_hd__nor2_1
XFILLER_159_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15597_ _15670_/A _15597_/B vssd1 vssd1 vccd1 vccd1 _15597_/X sky130_fd_sc_hd__or2_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ _25532_/Q vssd1 vssd1 vccd1 vccd1 _17336_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14548_ _14043_/X _14546_/X _14547_/X _13277_/A vssd1 vssd1 vccd1 vccd1 _14548_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_147_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17267_ _25510_/Q _17265_/B _17266_/Y vssd1 vssd1 vccd1 vccd1 _25510_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_131_wb_clk_i clkbuf_opt_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27227_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14479_ _14228_/A _14463_/X _14478_/X _13508_/A vssd1 vssd1 vccd1 vccd1 _14479_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_174_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19006_ _16521_/A _18972_/X _18973_/X _19005_/Y vssd1 vssd1 vccd1 vccd1 _19006_/X
+ sky130_fd_sc_hd__a211o_1
X_16218_ _26543_/Q _26151_/Q _16380_/B vssd1 vssd1 vccd1 vccd1 _16218_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17198_ _25492_/Q _17131_/B _17197_/Y _17188_/X vssd1 vssd1 vccd1 vccd1 _25492_/D
+ sky130_fd_sc_hd__o211a_1
X_16149_ _15020_/A _16144_/X _16148_/X _14678_/A vssd1 vssd1 vccd1 vccd1 _16149_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19908_ _19833_/A _19985_/C _19907_/Y _19941_/A vssd1 vssd1 vccd1 vccd1 _19908_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_229_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_257_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19839_ _19839_/A _27074_/Q vssd1 vssd1 vccd1 vccd1 _19841_/A sky130_fd_sc_hd__xnor2_1
XFILLER_96_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22850_ _22850_/A vssd1 vssd1 vccd1 vccd1 _26405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21801_ _26031_/Q _20878_/X _21805_/S vssd1 vssd1 vccd1 vccd1 _21802_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22781_ _26375_/Q _22691_/X _22789_/S vssd1 vssd1 vccd1 vccd1 _22782_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21732_ _20508_/X _26001_/Q _21732_/S vssd1 vssd1 vccd1 vccd1 _21733_/A sky130_fd_sc_hd__mux2_1
X_24520_ _26321_/Q _21869_/X _21871_/X input235/X _24501_/X vssd1 vssd1 vccd1 vccd1
+ _24520_/X sky130_fd_sc_hd__a221o_1
XFILLER_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21663_ _21663_/A vssd1 vssd1 vccd1 vccd1 _25972_/D sky130_fd_sc_hd__clkbuf_1
X_24451_ _24707_/B vssd1 vssd1 vccd1 vccd1 _24590_/A sky130_fd_sc_hd__clkinv_2
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20614_ _20613_/X _25721_/Q _20614_/S vssd1 vssd1 vccd1 vccd1 _20615_/A sky130_fd_sc_hd__mux2_1
X_23402_ _26636_/Q _23089_/X _23408_/S vssd1 vssd1 vccd1 vccd1 _23403_/A sky130_fd_sc_hd__mux2_1
X_24382_ _24473_/A vssd1 vssd1 vccd1 vccd1 _24382_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_27170_ _27173_/CLK _27170_/D vssd1 vssd1 vccd1 vccd1 _27170_/Q sky130_fd_sc_hd__dfxtp_1
X_21594_ _21594_/A vssd1 vssd1 vccd1 vccd1 _21594_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23333_ _20567_/X _26606_/Q _23335_/S vssd1 vssd1 vccd1 vccd1 _23334_/A sky130_fd_sc_hd__mux2_1
X_26121_ _27288_/CLK _26121_/D vssd1 vssd1 vccd1 vccd1 _26121_/Q sky130_fd_sc_hd__dfxtp_1
X_20545_ _23552_/A vssd1 vssd1 vccd1 vccd1 _23728_/A sky130_fd_sc_hd__buf_4
XFILLER_124_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23264_ _26575_/Q _23111_/X _23266_/S vssd1 vssd1 vccd1 vccd1 _23265_/A sky130_fd_sc_hd__mux2_1
X_26052_ _27287_/CLK _26052_/D vssd1 vssd1 vccd1 vccd1 _26052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20476_ _27098_/Q vssd1 vssd1 vccd1 vccd1 _20478_/A sky130_fd_sc_hd__inv_2
XFILLER_146_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22215_ _26187_/Q _22201_/X _22206_/X _22214_/X _22203_/X vssd1 vssd1 vccd1 vccd1
+ _22215_/X sky130_fd_sc_hd__a221o_1
X_25003_ _25138_/A vssd1 vssd1 vccd1 vccd1 _25003_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23195_ _23195_/A vssd1 vssd1 vccd1 vccd1 _26544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_279_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22146_ _22146_/A _22207_/S vssd1 vssd1 vccd1 vccd1 _22146_/X sky130_fd_sc_hd__or2b_1
XFILLER_161_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput370 _25901_/Q vssd1 vssd1 vccd1 vccd1 core_wb_stb_o sky130_fd_sc_hd__buf_2
Xoutput381 _17027_/X vssd1 vssd1 vccd1 vccd1 din0[14] sky130_fd_sc_hd__buf_2
XFILLER_121_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput392 _17041_/X vssd1 vssd1 vccd1 vccd1 din0[24] sky130_fd_sc_hd__buf_2
X_26954_ _26987_/CLK _26954_/D vssd1 vssd1 vccd1 vccd1 _26954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22077_ _26147_/Q _20932_/X _22077_/S vssd1 vssd1 vccd1 vccd1 _22078_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25905_ _26278_/CLK _25905_/D vssd1 vssd1 vccd1 vccd1 _25905_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_86_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21028_ _21050_/A vssd1 vssd1 vccd1 vccd1 _21037_/S sky130_fd_sc_hd__buf_4
XFILLER_75_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26885_ _26916_/CLK _26885_/D vssd1 vssd1 vccd1 vccd1 _26885_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25836_ _26595_/CLK _25836_/D vssd1 vssd1 vccd1 vccd1 _25836_/Q sky130_fd_sc_hd__dfxtp_1
X_13850_ _13818_/Y _13826_/Y _13839_/Y _13849_/Y _13638_/A vssd1 vssd1 vccd1 vccd1
+ _13850_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_75_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12801_ _13215_/A _25578_/Q vssd1 vssd1 vccd1 vccd1 _14188_/A sky130_fd_sc_hd__and2_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25767_ _26594_/CLK _25767_/D vssd1 vssd1 vccd1 vccd1 _25767_/Q sky130_fd_sc_hd__dfxtp_1
X_13781_ _13266_/A _25837_/Q _26037_/Q _13262_/A _13832_/A vssd1 vssd1 vccd1 vccd1
+ _13781_/X sky130_fd_sc_hd__a221o_1
XFILLER_56_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22979_ _22979_/A vssd1 vssd1 vccd1 vccd1 _26462_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_409 _17046_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15520_ _14727_/A _15518_/X _15519_/X _13304_/A vssd1 vssd1 vccd1 vccd1 _15521_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _13943_/A vssd1 vssd1 vccd1 vccd1 _12738_/C sky130_fd_sc_hd__buf_2
X_24718_ hold2/A vssd1 vssd1 vccd1 vccd1 _24719_/B sky130_fd_sc_hd__inv_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25698_ _26594_/CLK _25698_/D vssd1 vssd1 vccd1 vccd1 _25698_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_204_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15451_ _15449_/X _15450_/X _15559_/S vssd1 vssd1 vccd1 vccd1 _15451_/X sky130_fd_sc_hd__mux2_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24649_ _24739_/A _24649_/B vssd1 vssd1 vccd1 vccd1 _24649_/Y sky130_fd_sc_hd__nand2_2
XFILLER_203_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ input118/X input133/X _14402_/S vssd1 vssd1 vccd1 vccd1 _14403_/B sky130_fd_sc_hd__mux2_8
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18170_ _18462_/A vssd1 vssd1 vccd1 vccd1 _18827_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15382_ _26540_/Q _26148_/Q _16053_/S vssd1 vssd1 vccd1 vccd1 _15382_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17121_ _25469_/Q _17114_/X _17117_/X _17120_/X vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__o211a_1
X_26319_ _26319_/CLK _26319_/D vssd1 vssd1 vccd1 vccd1 _26319_/Q sky130_fd_sc_hd__dfxtp_4
X_14333_ _12673_/A _27297_/Q _26554_/Q _14173_/B _13022_/A vssd1 vssd1 vccd1 vccd1
+ _14333_/X sky130_fd_sc_hd__o221a_1
XFILLER_183_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27299_ _27299_/CLK _27299_/D vssd1 vssd1 vccd1 vccd1 _27299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17052_ _26584_/Q _17039_/X _20790_/C _17051_/X vssd1 vssd1 vccd1 vccd1 _17052_/X
+ sky130_fd_sc_hd__a22o_4
X_14264_ _14262_/X _14263_/X _14264_/S vssd1 vssd1 vccd1 vccd1 _14264_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16003_ _15205_/A _16001_/X _16002_/X _13976_/X vssd1 vssd1 vccd1 vccd1 _16003_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_137_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13215_ _13215_/A _25582_/Q vssd1 vssd1 vccd1 vccd1 _13808_/A sky130_fd_sc_hd__nand2_2
X_14195_ _14192_/X _14193_/Y _16585_/A vssd1 vssd1 vccd1 vccd1 _16711_/A sky130_fd_sc_hd__o21a_1
XFILLER_83_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13146_ _14513_/S vssd1 vssd1 vccd1 vccd1 _14263_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_253_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13077_ _15984_/B vssd1 vssd1 vccd1 vccd1 _15468_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_151_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17954_ _15701_/B _15788_/B _17954_/S vssd1 vssd1 vccd1 vccd1 _17954_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16905_ _16905_/A vssd1 vssd1 vccd1 vccd1 _16905_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17885_ _17927_/A _17933_/S vssd1 vssd1 vccd1 vccd1 _17973_/A sky130_fd_sc_hd__or2_2
XFILLER_39_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19624_ _27056_/Q _26061_/Q _19624_/C vssd1 vssd1 vccd1 vccd1 _19624_/X sky130_fd_sc_hd__and3_1
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16836_ _16973_/B vssd1 vssd1 vccd1 vccd1 _16836_/X sky130_fd_sc_hd__buf_2
XFILLER_93_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19555_ _20644_/A vssd1 vssd1 vccd1 vccd1 _19555_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16767_ _22518_/A _16756_/X _16757_/X _16638_/A vssd1 vssd1 vccd1 vccd1 _16767_/X
+ sky130_fd_sc_hd__a22o_2
X_13979_ _13466_/A _23530_/A _13978_/X _13683_/X vssd1 vssd1 vccd1 vccd1 _19800_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_20_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18506_ _27206_/Q _19258_/B vssd1 vssd1 vccd1 vccd1 _18506_/X sky130_fd_sc_hd__and2_1
XFILLER_207_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15718_ _25844_/Q _26044_/Q _15988_/S vssd1 vssd1 vccd1 vccd1 _15718_/X sky130_fd_sc_hd__mux2_1
X_19486_ _19568_/B vssd1 vssd1 vccd1 vccd1 _19497_/B sky130_fd_sc_hd__clkbuf_1
X_16698_ _21190_/A _21709_/B vssd1 vssd1 vccd1 vccd1 _16826_/A sky130_fd_sc_hd__nor2_2
XFILLER_34_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18437_ _18437_/A vssd1 vssd1 vccd1 vccd1 _18437_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_278_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15649_ _26668_/Q _16151_/S _15648_/X _15169_/A vssd1 vssd1 vccd1 vccd1 _15649_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_222_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18368_ _18368_/A vssd1 vssd1 vccd1 vccd1 _18368_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_187_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17319_ _17317_/X _17322_/C _17318_/X vssd1 vssd1 vccd1 vccd1 _17319_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18299_ _26945_/Q _18826_/A _18827_/A _26977_/Q vssd1 vssd1 vccd1 vccd1 _18299_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20330_ _19283_/A _20355_/A _20329_/Y _20357_/A vssd1 vssd1 vccd1 vccd1 _20353_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_190_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20261_ _20261_/A _20261_/B vssd1 vssd1 vccd1 vccd1 _20262_/B sky130_fd_sc_hd__nor2_1
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22000_ _22000_/A vssd1 vssd1 vccd1 vccd1 _26112_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20192_ _20379_/A vssd1 vssd1 vccd1 vccd1 _20426_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput109 dout1[11] vssd1 vssd1 vccd1 vccd1 input109/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23951_ _23951_/A vssd1 vssd1 vccd1 vccd1 _26851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22902_ _22902_/A vssd1 vssd1 vccd1 vccd1 _26428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26670_ _26823_/CLK _26670_/D vssd1 vssd1 vccd1 vccd1 _26670_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23882_ _23715_/X _26821_/Q _23882_/S vssd1 vssd1 vccd1 vccd1 _23883_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25621_ _25624_/CLK _25621_/D vssd1 vssd1 vccd1 vccd1 _25621_/Q sky130_fd_sc_hd__dfxtp_4
X_22833_ _22833_/A vssd1 vssd1 vccd1 vccd1 _26397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25552_ _27000_/CLK _25552_/D vssd1 vssd1 vccd1 vccd1 _25552_/Q sky130_fd_sc_hd__dfxtp_1
X_22764_ _22764_/A vssd1 vssd1 vccd1 vccd1 _26367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_253_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24503_ _24370_/S _25622_/Q _24502_/X vssd1 vssd1 vccd1 vccd1 _24969_/A sky130_fd_sc_hd__o21ai_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21715_ _21715_/A vssd1 vssd1 vccd1 vccd1 _21715_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22695_ _23738_/A vssd1 vssd1 vccd1 vccd1 _22695_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25483_ _25590_/CLK _25483_/D vssd1 vssd1 vccd1 vccd1 _25483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27222_ _27227_/CLK _27222_/D vssd1 vssd1 vccd1 vccd1 _27222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24434_ _24434_/A _24582_/A vssd1 vssd1 vccd1 vccd1 _24434_/Y sky130_fd_sc_hd__nand2_1
X_21646_ input67/X input102/X _21646_/S vssd1 vssd1 vccd1 vccd1 _21647_/A sky130_fd_sc_hd__mux2_8
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27153_ _27156_/CLK _27153_/D vssd1 vssd1 vccd1 vccd1 _27153_/Q sky130_fd_sc_hd__dfxtp_4
X_24365_ _24454_/A vssd1 vssd1 vccd1 vccd1 _24370_/S sky130_fd_sc_hd__clkbuf_4
X_21577_ _19283_/A _21545_/X _21563_/X _21576_/X vssd1 vssd1 vccd1 vccd1 _21577_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_138_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26104_ _26601_/CLK _26104_/D vssd1 vssd1 vccd1 vccd1 _26104_/Q sky130_fd_sc_hd__dfxtp_4
X_23316_ _20533_/X _26598_/Q _23324_/S vssd1 vssd1 vccd1 vccd1 _23317_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20528_ _23539_/A vssd1 vssd1 vccd1 vccd1 _23715_/A sky130_fd_sc_hd__buf_4
X_24296_ _24312_/A _24301_/C vssd1 vssd1 vccd1 vccd1 _24296_/Y sky130_fd_sc_hd__nor2_1
XFILLER_181_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27084_ _27087_/CLK _27084_/D vssd1 vssd1 vccd1 vccd1 _27084_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_126_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26035_ _26594_/CLK _26035_/D vssd1 vssd1 vccd1 vccd1 _26035_/Q sky130_fd_sc_hd__dfxtp_1
X_23247_ _26567_/Q _23085_/X _23255_/S vssd1 vssd1 vccd1 vccd1 _23248_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20459_ _20434_/A _20434_/B _20458_/X vssd1 vssd1 vccd1 vccd1 _20460_/B sky130_fd_sc_hd__o21a_1
XFILLER_273_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13000_ _13185_/A _25589_/Q vssd1 vssd1 vccd1 vccd1 _14354_/S sky130_fd_sc_hd__nand2_4
XFILLER_140_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23178_ _23178_/A vssd1 vssd1 vccd1 vccd1 _26536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_279_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22129_ _26162_/Q _22122_/X _22124_/X input256/X _22118_/X vssd1 vssd1 vccd1 vccd1
+ _22129_/X sky130_fd_sc_hd__a221o_1
XFILLER_279_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26937_ _27324_/CLK _26937_/D vssd1 vssd1 vccd1 vccd1 _26937_/Q sky130_fd_sc_hd__dfxtp_1
X_14951_ _26808_/Q _26452_/Q _14953_/S vssd1 vssd1 vccd1 vccd1 _14951_/X sky130_fd_sc_hd__mux2_1
XTAP_5854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13902_ _13009_/A _23533_/A _13901_/X _13027_/A vssd1 vssd1 vccd1 vccd1 _16833_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17670_ _17769_/A _18307_/A _17670_/C vssd1 vssd1 vccd1 vccd1 _18010_/C sky130_fd_sc_hd__and3_2
XTAP_5898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26868_ _26932_/CLK _26868_/D vssd1 vssd1 vccd1 vccd1 _26868_/Q sky130_fd_sc_hd__dfxtp_1
X_14882_ _14881_/A _14877_/X _14881_/Y _14706_/X vssd1 vssd1 vccd1 vccd1 _14882_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_263_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16621_ _16621_/A _16621_/B vssd1 vssd1 vccd1 vccd1 _17835_/C sky130_fd_sc_hd__nor2_1
XFILLER_63_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13833_ _15509_/A _13829_/X _13831_/X _15311_/A vssd1 vssd1 vccd1 vccd1 _13839_/A
+ sky130_fd_sc_hd__o211a_1
X_25819_ _26900_/CLK _25819_/D vssd1 vssd1 vccd1 vccd1 _25819_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26799_ _26799_/CLK _26799_/D vssd1 vssd1 vccd1 vccd1 _26799_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_206 _20701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19340_ _18555_/X _19330_/X _19339_/X vssd1 vssd1 vccd1 vccd1 _19340_/X sky130_fd_sc_hd__a21o_4
XINSDIODE2_217 _20120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16552_ _16462_/A _16461_/A _16461_/B _19427_/S vssd1 vssd1 vccd1 vccd1 _16553_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_262_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13764_ _13472_/X _26596_/Q _13492_/X _26336_/Q _15606_/A vssd1 vssd1 vccd1 vccd1
+ _13764_/X sky130_fd_sc_hd__o221a_1
XFILLER_44_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_228 _19971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_239 _16636_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15503_ _15491_/X _27281_/Q _26474_/Q _15850_/S _13806_/X vssd1 vssd1 vccd1 vccd1
+ _15503_/X sky130_fd_sc_hd__a221o_1
XFILLER_204_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12715_ _16328_/A vssd1 vssd1 vccd1 vccd1 _15285_/A sky130_fd_sc_hd__buf_2
XFILLER_16_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19271_ _19482_/B _19271_/B _19271_/C vssd1 vssd1 vccd1 vccd1 _19271_/X sky130_fd_sc_hd__or3_4
X_16483_ _16490_/B vssd1 vssd1 vccd1 vccd1 _16493_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_241_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13695_ _13719_/A vssd1 vssd1 vccd1 vccd1 _16050_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_70_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18222_ _18027_/X _18150_/X _18221_/X _18976_/A vssd1 vssd1 vccd1 vccd1 _18223_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_231_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15434_ _19100_/A vssd1 vssd1 vccd1 vccd1 _20194_/A sky130_fd_sc_hd__inv_2
XFILLER_87_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18153_ _19069_/A vssd1 vssd1 vccd1 vccd1 _18154_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_175_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15365_ _27283_/Q _26476_/Q _16161_/S vssd1 vssd1 vccd1 vccd1 _15365_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17104_ _17514_/A vssd1 vssd1 vccd1 vccd1 _17210_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14316_ _13638_/A _23520_/A _14315_/X _13683_/X vssd1 vssd1 vccd1 vccd1 _19700_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_117_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18084_ _18343_/A _18859_/B _18364_/A vssd1 vssd1 vccd1 vccd1 _18084_/X sky130_fd_sc_hd__a21bo_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15296_ _15110_/A _26898_/Q _26770_/Q _15422_/S _14770_/A vssd1 vssd1 vccd1 vccd1
+ _15296_/X sky130_fd_sc_hd__a221o_1
XFILLER_156_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17035_ _17063_/A vssd1 vssd1 vccd1 vccd1 _17035_/X sky130_fd_sc_hd__clkbuf_2
X_14247_ _27298_/Q _26555_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _14247_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14178_ _14176_/X _14177_/X _14178_/S vssd1 vssd1 vccd1 vccd1 _14178_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13129_ _15567_/S vssd1 vssd1 vccd1 vccd1 _14870_/A sky130_fd_sc_hd__clkbuf_4
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _27216_/Q _19462_/B vssd1 vssd1 vccd1 vccd1 _18986_/X sky130_fd_sc_hd__and2_1
XFILLER_258_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ _17801_/B _17787_/B _17949_/S vssd1 vssd1 vccd1 vccd1 _17937_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17868_ _17957_/S vssd1 vssd1 vccd1 vccd1 _17909_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_282_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19607_ _19607_/A _19607_/B vssd1 vssd1 vccd1 vccd1 _19607_/X sky130_fd_sc_hd__or2_1
X_16819_ _16819_/A vssd1 vssd1 vccd1 vccd1 _16819_/X sky130_fd_sc_hd__clkbuf_1
X_17799_ _14192_/X _14193_/Y _17809_/A vssd1 vssd1 vccd1 vccd1 _17986_/A sky130_fd_sc_hd__o21ai_4
XFILLER_282_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19538_ _19551_/A vssd1 vssd1 vccd1 vccd1 _19538_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_207_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19469_ _25564_/Q _18763_/X _19468_/X _18767_/X _18768_/X vssd1 vssd1 vccd1 vccd1
+ _19469_/X sky130_fd_sc_hd__a221o_1
XFILLER_22_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21500_ _25866_/Q vssd1 vssd1 vccd1 vccd1 _21553_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22480_ _22480_/A _22480_/B vssd1 vssd1 vccd1 vccd1 _22481_/A sky130_fd_sc_hd__and2_1
X_21431_ _21587_/A vssd1 vssd1 vccd1 vccd1 _21431_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24150_ _24291_/A vssd1 vssd1 vccd1 vccd1 _24222_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_148_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21362_ _21559_/B vssd1 vssd1 vccd1 vccd1 _21416_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_147_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20313_ _20313_/A _20313_/B vssd1 vssd1 vccd1 vccd1 _20313_/X sky130_fd_sc_hd__or2_1
X_23101_ _23574_/A vssd1 vssd1 vccd1 vccd1 _23101_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_24081_ _26909_/Q _23514_/X _24087_/S vssd1 vssd1 vccd1 vccd1 _24082_/A sky130_fd_sc_hd__mux2_1
X_21293_ _21276_/X _21292_/X _21227_/X vssd1 vssd1 vccd1 vccd1 _21293_/Y sky130_fd_sc_hd__o21ai_1
Xinput80 dout0[43] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput91 dout0[53] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__clkbuf_1
X_23032_ _26487_/Q _22742_/X _23032_/S vssd1 vssd1 vccd1 vccd1 _23033_/A sky130_fd_sc_hd__mux2_1
X_20244_ _27154_/Q _20295_/B vssd1 vssd1 vccd1 vccd1 _20244_/X sky130_fd_sc_hd__and2_1
XFILLER_116_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20175_ _20174_/A _20174_/B _20200_/B vssd1 vssd1 vccd1 vccd1 _20175_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24983_ _27163_/Q _24913_/X _24982_/Y vssd1 vssd1 vccd1 vccd1 _27163_/D sky130_fd_sc_hd__o21a_1
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26722_ _26917_/CLK _26722_/D vssd1 vssd1 vccd1 vccd1 _26722_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23934_ _24002_/S vssd1 vssd1 vccd1 vccd1 _23943_/S sky130_fd_sc_hd__buf_6
XFILLER_18_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26653_ _27295_/CLK _26653_/D vssd1 vssd1 vccd1 vccd1 _26653_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23865_ _23690_/X _26813_/Q _23871_/S vssd1 vssd1 vccd1 vccd1 _23866_/A sky130_fd_sc_hd__mux2_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25604_ _25607_/CLK _25604_/D vssd1 vssd1 vccd1 vccd1 _25604_/Q sky130_fd_sc_hd__dfxtp_4
X_22816_ _22816_/A vssd1 vssd1 vccd1 vccd1 _26391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26584_ _27156_/CLK _26584_/D vssd1 vssd1 vccd1 vccd1 _26584_/Q sky130_fd_sc_hd__dfxtp_4
X_23796_ _23796_/A vssd1 vssd1 vccd1 vccd1 _26782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25535_ _26257_/CLK _25535_/D vssd1 vssd1 vccd1 vccd1 _25535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22747_ _22815_/S vssd1 vssd1 vccd1 vccd1 _22756_/S sky130_fd_sc_hd__buf_2
XFILLER_25_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13480_ _15300_/A _13471_/X _13476_/X _14757_/A vssd1 vssd1 vccd1 vccd1 _13497_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25466_ _25466_/A _25466_/B vssd1 vssd1 vccd1 vccd1 _25467_/A sky130_fd_sc_hd__or2_1
X_22678_ _22678_/A vssd1 vssd1 vccd1 vccd1 _26338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27205_ _27230_/CLK _27205_/D vssd1 vssd1 vccd1 vccd1 _27205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24417_ _26302_/Q _24393_/X _24394_/X input246/X _24395_/X vssd1 vssd1 vccd1 vccd1
+ _24417_/X sky130_fd_sc_hd__a221o_1
XFILLER_12_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21629_ _25965_/Q _21573_/X _21628_/Y _21597_/X vssd1 vssd1 vccd1 vccd1 _25965_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_201_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25397_ _25397_/A vssd1 vssd1 vccd1 vccd1 _27295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27136_ _27166_/CLK _27136_/D vssd1 vssd1 vccd1 vccd1 _27136_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15150_ _27255_/Q _16388_/B vssd1 vssd1 vccd1 vccd1 _15150_/X sky130_fd_sc_hd__or2_1
XFILLER_194_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24348_ _25494_/Q _17470_/A _24350_/S vssd1 vssd1 vccd1 vccd1 _24542_/B sky130_fd_sc_hd__mux2_1
XFILLER_138_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14101_ _12700_/A _14089_/X _14093_/X _14099_/Y _14421_/A vssd1 vssd1 vccd1 vccd1
+ _14101_/X sky130_fd_sc_hd__a221o_1
XFILLER_153_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27067_ _27164_/CLK _27067_/D vssd1 vssd1 vccd1 vccd1 _27067_/Q sky130_fd_sc_hd__dfxtp_1
X_15081_ _19798_/A _16451_/S _15080_/Y vssd1 vssd1 vccd1 vccd1 _17787_/A sky130_fd_sc_hd__o21ai_4
X_24279_ _24312_/A _24284_/C vssd1 vssd1 vccd1 vccd1 _24279_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14032_ _14404_/A _14032_/B vssd1 vssd1 vccd1 vccd1 _15874_/C sky130_fd_sc_hd__nand2_1
X_26018_ _26673_/CLK _26018_/D vssd1 vssd1 vccd1 vccd1 _26018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18840_ _19234_/A _18836_/Y _18837_/X _18848_/B _18839_/X vssd1 vssd1 vccd1 vccd1
+ _18840_/X sky130_fd_sc_hd__o32a_2
XFILLER_122_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18771_ _25513_/Q _18746_/X _18762_/X _18769_/X _18770_/X vssd1 vssd1 vccd1 vccd1
+ _18771_/X sky130_fd_sc_hd__o221a_1
XFILLER_79_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15983_ _15979_/X _15982_/X _15983_/S vssd1 vssd1 vccd1 vccd1 _15983_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17722_ _17747_/B _17722_/B _17736_/A vssd1 vssd1 vccd1 vccd1 _17730_/A sky130_fd_sc_hd__and3_4
XFILLER_76_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14934_ _16458_/A _17852_/B vssd1 vssd1 vccd1 vccd1 _16556_/A sky130_fd_sc_hd__nor2_1
XTAP_5684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17653_ _17653_/A _17653_/B _17653_/C vssd1 vssd1 vccd1 vccd1 _17653_/X sky130_fd_sc_hd__or3_1
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14865_ _26681_/Q _25721_/Q _14878_/S vssd1 vssd1 vccd1 vccd1 _14865_/X sky130_fd_sc_hd__mux2_1
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16604_ _16604_/A _16697_/D vssd1 vssd1 vccd1 vccd1 _20799_/B sky130_fd_sc_hd__nor2_4
X_13816_ _13813_/X _27270_/Q _26463_/Q _13535_/S _15776_/A vssd1 vssd1 vccd1 vccd1
+ _13816_/X sky130_fd_sc_hd__a221o_1
X_17584_ _17635_/A vssd1 vssd1 vccd1 vccd1 _17584_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14796_ _26938_/Q _26422_/Q _14811_/S vssd1 vssd1 vccd1 vccd1 _14796_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19323_ _16454_/B _18548_/X _19321_/Y _16794_/B _19322_/Y vssd1 vssd1 vccd1 vccd1
+ _19323_/X sky130_fd_sc_hd__o221a_1
XFILLER_50_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16535_ _16513_/A _25789_/Q _16541_/S _26875_/Q _16524_/A vssd1 vssd1 vccd1 vccd1
+ _16535_/X sky130_fd_sc_hd__o221a_1
X_13747_ _14031_/A _13747_/B vssd1 vssd1 vccd1 vccd1 _13748_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19254_ _16481_/A _19218_/X _19251_/Y _19252_/X _19253_/X vssd1 vssd1 vccd1 vccd1
+ _19254_/X sky130_fd_sc_hd__a221o_2
X_16466_ _16639_/A _15706_/X _16464_/X _16465_/X vssd1 vssd1 vccd1 vccd1 _23609_/A
+ sky130_fd_sc_hd__a31o_4
X_13678_ _16014_/S vssd1 vssd1 vccd1 vccd1 _16013_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_32_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18205_ _18199_/X _18203_/X _18487_/A vssd1 vssd1 vccd1 vccd1 _18205_/X sky130_fd_sc_hd__mux2_1
X_15417_ _15417_/A _15417_/B vssd1 vssd1 vccd1 vccd1 _15417_/X sky130_fd_sc_hd__or2_1
XPHY_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19185_ _19352_/A vssd1 vssd1 vccd1 vccd1 _19185_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16397_ _16395_/X _16396_/X _16397_/S vssd1 vssd1 vccd1 vccd1 _16397_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26889_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18136_ _18435_/A _18133_/X _18135_/X vssd1 vssd1 vccd1 vccd1 _18136_/Y sky130_fd_sc_hd__a21oi_1
X_15348_ _14601_/A _15346_/Y _15347_/X _15135_/X vssd1 vssd1 vccd1 vccd1 _15348_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_184_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18067_ _17929_/X _17922_/X _18067_/S vssd1 vssd1 vccd1 vccd1 _18067_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15279_ _26802_/Q _26446_/Q _16315_/S vssd1 vssd1 vccd1 vccd1 _15279_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17018_ _17015_/X _16844_/B _17017_/X input245/X vssd1 vssd1 vccd1 vccd1 _17018_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_259_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18969_ _16517_/X _18890_/X _18967_/Y _18968_/X _18933_/X vssd1 vssd1 vccd1 vccd1
+ _18969_/X sky130_fd_sc_hd__a221o_4
XFILLER_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21980_ _21980_/A vssd1 vssd1 vccd1 vccd1 _26103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_255_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20931_ _20931_/A vssd1 vssd1 vccd1 vccd1 _25847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20862_ _25827_/Q vssd1 vssd1 vccd1 vccd1 _20863_/A sky130_fd_sc_hd__clkbuf_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23650_ _26732_/Q _23562_/X _23656_/S vssd1 vssd1 vccd1 vccd1 _23651_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22601_ _22593_/X _22599_/Y _22600_/X vssd1 vssd1 vccd1 vccd1 _26315_/D sky130_fd_sc_hd__a21oi_1
XFILLER_23_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 INSDIODE2_273/DIODE
+ sky130_fd_sc_hd__clkbuf_4
X_23581_ _23581_/A vssd1 vssd1 vccd1 vccd1 _23581_/X sky130_fd_sc_hd__clkbuf_2
X_20793_ _20793_/A vssd1 vssd1 vccd1 vccd1 _25791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25320_ _25320_/A vssd1 vssd1 vccd1 vccd1 _27262_/D sky130_fd_sc_hd__clkbuf_1
X_22532_ _22532_/A vssd1 vssd1 vccd1 vccd1 _26290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25251_ _25319_/S vssd1 vssd1 vccd1 vccd1 _25260_/S sky130_fd_sc_hd__buf_4
XFILLER_33_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22463_ _26257_/Q _22470_/B vssd1 vssd1 vccd1 vccd1 _22463_/X sky130_fd_sc_hd__or2_1
XFILLER_194_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24202_ _26957_/Q _24203_/C _26958_/Q vssd1 vssd1 vccd1 vccd1 _24204_/B sky130_fd_sc_hd__a21oi_1
X_21414_ _21544_/A vssd1 vssd1 vccd1 vccd1 _21414_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22394_ _22394_/A _22406_/A vssd1 vssd1 vccd1 vccd1 _22395_/B sky130_fd_sc_hd__and2_1
XFILLER_176_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25182_ _24649_/B _25172_/X _25175_/X _27201_/Q _25179_/X vssd1 vssd1 vccd1 vccd1
+ _27201_/D sky130_fd_sc_hd__o221a_1
XFILLER_163_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21345_ _25476_/Q _21620_/B vssd1 vssd1 vccd1 vccd1 _21345_/X sky130_fd_sc_hd__or2_1
X_24133_ _24133_/A vssd1 vssd1 vccd1 vccd1 _24142_/S sky130_fd_sc_hd__buf_4
XFILLER_108_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21276_ _21276_/A vssd1 vssd1 vccd1 vccd1 _21276_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_24064_ _26902_/Q _23594_/X _24070_/S vssd1 vssd1 vccd1 vccd1 _24065_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23015_ _26479_/Q _22717_/X _23017_/S vssd1 vssd1 vccd1 vccd1 _23016_/A sky130_fd_sc_hd__mux2_1
X_20227_ _20227_/A _20227_/B vssd1 vssd1 vccd1 vccd1 _20227_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20158_ _27151_/Q _27085_/Q vssd1 vssd1 vccd1 vccd1 _20158_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24966_ _24966_/A vssd1 vssd1 vccd1 vccd1 _24966_/X sky130_fd_sc_hd__buf_2
X_12980_ _13916_/B _13916_/C _12948_/C _12964_/A vssd1 vssd1 vccd1 vccd1 _12982_/A
+ sky130_fd_sc_hd__a31o_1
X_20089_ _20089_/A vssd1 vssd1 vccd1 vccd1 _20125_/B sky130_fd_sc_hd__clkbuf_2
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26705_ _27252_/CLK _26705_/D vssd1 vssd1 vccd1 vccd1 _26705_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23917_ _23917_/A vssd1 vssd1 vccd1 vccd1 _23926_/S sky130_fd_sc_hd__buf_6
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24897_ _20703_/A _19724_/X _24772_/Y _24782_/X vssd1 vssd1 vccd1 vccd1 _24897_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14650_ _14650_/A vssd1 vssd1 vccd1 vccd1 _14650_/X sky130_fd_sc_hd__buf_2
X_26636_ _26799_/CLK _26636_/D vssd1 vssd1 vccd1 vccd1 _26636_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23848_ _23770_/X _26806_/Q _23854_/S vssd1 vssd1 vccd1 vccd1 _23849_/A sky130_fd_sc_hd__mux2_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13601_ _26853_/Q _25767_/Q _15805_/S vssd1 vssd1 vccd1 vccd1 _13601_/X sky130_fd_sc_hd__mux2_1
XFILLER_261_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26567_ _27313_/CLK _26567_/D vssd1 vssd1 vccd1 vccd1 _26567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14581_ _17809_/A vssd1 vssd1 vccd1 vccd1 _16122_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23779_ _23779_/A vssd1 vssd1 vccd1 vccd1 _23779_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16320_ _16318_/X _16319_/X _16320_/S vssd1 vssd1 vccd1 vccd1 _16320_/X sky130_fd_sc_hd__mux2_1
X_13532_ _15836_/A vssd1 vssd1 vccd1 vccd1 _13532_/X sky130_fd_sc_hd__buf_4
X_25518_ _25518_/CLK _25518_/D vssd1 vssd1 vccd1 vccd1 _25518_/Q sky130_fd_sc_hd__dfxtp_1
X_26498_ _27309_/CLK _26498_/D vssd1 vssd1 vccd1 vccd1 _26498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16251_ _13105_/B _16451_/S _15244_/X _16250_/Y vssd1 vssd1 vccd1 vccd1 _17795_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_174_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25449_ _25449_/A vssd1 vssd1 vccd1 vccd1 _27319_/D sky130_fd_sc_hd__clkbuf_1
X_13463_ _15482_/A _16852_/A _13458_/X _15526_/S vssd1 vssd1 vccd1 vccd1 _13552_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_139_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15202_ _15422_/S vssd1 vssd1 vccd1 vccd1 _16436_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_138_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16182_ _25850_/Q _26050_/Q _16182_/S vssd1 vssd1 vccd1 vccd1 _16182_/X sky130_fd_sc_hd__mux2_1
X_13394_ input108/X input143/X _13741_/S vssd1 vssd1 vccd1 vccd1 _13395_/B sky130_fd_sc_hd__mux2_8
XFILLER_139_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15133_ _17846_/A vssd1 vssd1 vccd1 vccd1 _19325_/A sky130_fd_sc_hd__clkbuf_4
X_27119_ _27122_/CLK _27119_/D vssd1 vssd1 vccd1 vccd1 _27119_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19941_ _19941_/A vssd1 vssd1 vccd1 vccd1 _19941_/X sky130_fd_sc_hd__buf_2
X_15064_ _15167_/A vssd1 vssd1 vccd1 vccd1 _15065_/A sky130_fd_sc_hd__buf_2
XFILLER_153_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14015_ _13857_/X _14010_/X _14014_/X _13162_/A vssd1 vssd1 vccd1 vccd1 _14015_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19872_ _25208_/B vssd1 vssd1 vccd1 vccd1 _22130_/A sky130_fd_sc_hd__buf_6
XFILLER_268_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18823_ _18823_/A vssd1 vssd1 vccd1 vccd1 _18823_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_256_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_156_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27196_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_228_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15966_ _25809_/Q _13441_/S _15970_/S _15965_/X vssd1 vssd1 vccd1 vccd1 _15966_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18754_ _27081_/Q _18751_/X _18752_/X _27179_/Q _18753_/X vssd1 vssd1 vccd1 vccd1
+ _18754_/X sky130_fd_sc_hd__a221o_1
XTAP_5470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput270 partID[15] vssd1 vssd1 vccd1 vccd1 input270/X sky130_fd_sc_hd__clkbuf_2
XTAP_5481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput281 versionID[1] vssd1 vssd1 vccd1 vccd1 input281/X sky130_fd_sc_hd__clkbuf_2
XFILLER_283_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17705_ _17697_/A _13105_/B _17703_/X _17739_/C vssd1 vssd1 vccd1 vccd1 _18116_/A
+ sky130_fd_sc_hd__a211o_1
X_14917_ _15095_/S vssd1 vssd1 vccd1 vccd1 _14917_/X sky130_fd_sc_hd__buf_2
XFILLER_76_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15897_ _25810_/Q _27244_/Q _15904_/S vssd1 vssd1 vccd1 vccd1 _15897_/X sky130_fd_sc_hd__mux2_2
X_18685_ _18311_/X _18684_/X _18685_/S vssd1 vssd1 vccd1 vccd1 _18685_/X sky130_fd_sc_hd__mux2_1
XFILLER_252_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17636_ _17534_/X _17627_/X _13385_/X _17536_/X _25928_/Q vssd1 vssd1 vccd1 vccd1
+ _17636_/Y sky130_fd_sc_hd__o32ai_1
X_14848_ _14952_/S _14845_/X _14847_/X _14650_/A vssd1 vssd1 vccd1 vccd1 _14848_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17567_ _17575_/A _17567_/B vssd1 vssd1 vccd1 vccd1 _25573_/D sky130_fd_sc_hd__nor2_1
X_14779_ _14779_/A vssd1 vssd1 vccd1 vccd1 _20119_/A sky130_fd_sc_hd__buf_8
XFILLER_211_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19306_ _25559_/Q _18825_/X _19305_/X _18829_/X _18830_/X vssd1 vssd1 vccd1 vccd1
+ _19306_/X sky130_fd_sc_hd__a221o_1
X_16518_ _26811_/Q _26455_/Q _16523_/S vssd1 vssd1 vccd1 vccd1 _16518_/X sky130_fd_sc_hd__mux2_1
X_17498_ _24340_/S vssd1 vssd1 vccd1 vccd1 _24454_/A sky130_fd_sc_hd__buf_2
XFILLER_17_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19237_ _19237_/A _19237_/B _19237_/C vssd1 vssd1 vccd1 vccd1 _19238_/B sky130_fd_sc_hd__nand3_1
X_16449_ _16281_/S _23597_/A _16448_/X _16282_/A vssd1 vssd1 vccd1 vccd1 _19341_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_104_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19168_ _27059_/Q _18811_/X _19165_/X _19167_/X _18823_/X vssd1 vssd1 vccd1 vccd1
+ _19168_/X sky130_fd_sc_hd__o221a_2
XFILLER_158_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18119_ _18119_/A _18119_/B vssd1 vssd1 vccd1 vccd1 _18120_/D sky130_fd_sc_hd__nor2_1
X_19099_ _18437_/A _19089_/X _19098_/X vssd1 vssd1 vccd1 vccd1 _19099_/X sky130_fd_sc_hd__a21o_4
X_21130_ _21166_/A vssd1 vssd1 vccd1 vccd1 _21130_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21061_ _25899_/Q _20967_/X _21063_/S vssd1 vssd1 vccd1 vccd1 _21062_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20012_ _16591_/A _19914_/X _19774_/B _20089_/A vssd1 vssd1 vccd1 vccd1 _20039_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24820_ _24818_/Y _24819_/X _24816_/X vssd1 vssd1 vccd1 vccd1 _27110_/D sky130_fd_sc_hd__a21oi_1
XFILLER_100_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24751_ _24781_/A _24751_/B vssd1 vssd1 vccd1 vccd1 _25143_/A sky130_fd_sc_hd__nand2_4
X_21963_ _22031_/S vssd1 vssd1 vccd1 vccd1 _21972_/S sky130_fd_sc_hd__buf_2
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23702_ _23702_/A vssd1 vssd1 vccd1 vccd1 _23702_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20914_ _25842_/Q _20913_/X _20917_/S vssd1 vssd1 vccd1 vccd1 _20915_/A sky130_fd_sc_hd__mux2_1
XFILLER_254_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24682_ _24682_/A _24682_/B vssd1 vssd1 vccd1 vccd1 _24682_/Y sky130_fd_sc_hd__nand2_2
X_21894_ _20496_/X _26065_/Q _21900_/S vssd1 vssd1 vccd1 vccd1 _21895_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26421_ _27292_/CLK _26421_/D vssd1 vssd1 vccd1 vccd1 _26421_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23633_ _23633_/A vssd1 vssd1 vccd1 vccd1 _26724_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20845_ _20845_/A vssd1 vssd1 vccd1 vccd1 _25818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26352_ _26611_/CLK _26352_/D vssd1 vssd1 vccd1 vccd1 _26352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23564_ _23564_/A vssd1 vssd1 vccd1 vccd1 _26700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20776_ _20776_/A vssd1 vssd1 vccd1 vccd1 _25783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25303_ _25303_/A vssd1 vssd1 vccd1 vccd1 _27254_/D sky130_fd_sc_hd__clkbuf_1
X_22515_ _22515_/A vssd1 vssd1 vccd1 vccd1 _22524_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_211_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26283_ _26286_/CLK _26283_/D vssd1 vssd1 vccd1 vccd1 _26283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23495_ _23495_/A vssd1 vssd1 vccd1 vccd1 _26677_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25234_ _27223_/Q _25225_/X _25228_/X _24746_/B _25233_/X vssd1 vssd1 vccd1 vccd1
+ _27223_/D sky130_fd_sc_hd__o221a_1
XFILLER_13_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22446_ _22459_/A vssd1 vssd1 vccd1 vccd1 _22446_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25165_ _27197_/Q _25137_/X _25164_/X vssd1 vssd1 vccd1 vccd1 _27197_/D sky130_fd_sc_hd__o21ba_1
XFILLER_108_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22377_ _22377_/A _22377_/B vssd1 vssd1 vccd1 vccd1 _22378_/A sky130_fd_sc_hd__and2_1
XFILLER_129_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24116_ _26925_/Q _23565_/X _24120_/S vssd1 vssd1 vccd1 vccd1 _24117_/A sky130_fd_sc_hd__mux2_1
X_21328_ _21231_/X _21327_/X _21259_/A vssd1 vssd1 vccd1 vccd1 _21328_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_108_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25096_ _27183_/Q _25085_/X _25095_/X vssd1 vssd1 vccd1 vccd1 _27183_/D sky130_fd_sc_hd__o21ba_1
XFILLER_151_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21259_ _21259_/A vssd1 vssd1 vccd1 vccd1 _21259_/X sky130_fd_sc_hd__buf_6
X_24047_ _24047_/A vssd1 vssd1 vccd1 vccd1 _26894_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15820_ _25706_/Q _15820_/B vssd1 vssd1 vccd1 vccd1 _15820_/X sky130_fd_sc_hd__or2_1
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25998_ _26240_/CLK _25998_/D vssd1 vssd1 vccd1 vccd1 _25998_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _26667_/Q _25707_/Q _15930_/S vssd1 vssd1 vccd1 vccd1 _15751_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ _12866_/X _13916_/B _12963_/C _12963_/D vssd1 vssd1 vccd1 vccd1 _12964_/A
+ sky130_fd_sc_hd__and4b_1
X_24949_ _25221_/A vssd1 vssd1 vccd1 vccd1 _24949_/X sky130_fd_sc_hd__dlymetal6s2s_1
XINSDIODE2_60 _20648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_71 _22638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_82 _23712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _12777_/A _26714_/Q _26842_/Q _14652_/S _16484_/A vssd1 vssd1 vccd1 vccd1
+ _14702_/X sky130_fd_sc_hd__a221o_1
X_18470_ _25507_/Q _18444_/X _18457_/X _18467_/X _18469_/X vssd1 vssd1 vccd1 vccd1
+ _18470_/X sky130_fd_sc_hd__o221a_1
XFILLER_205_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_93 _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15682_ _16104_/A _15682_/B vssd1 vssd1 vccd1 vccd1 _15682_/X sky130_fd_sc_hd__or2_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _13561_/A vssd1 vssd1 vccd1 vccd1 _17653_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _17430_/A _17427_/C vssd1 vssd1 vccd1 vccd1 _17421_/Y sky130_fd_sc_hd__nor2_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26619_ _26939_/CLK _26619_/D vssd1 vssd1 vccd1 vccd1 _26619_/Q sky130_fd_sc_hd__dfxtp_1
X_14633_ _16319_/S vssd1 vssd1 vccd1 vccd1 _16242_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _17380_/A _17352_/B _17353_/B vssd1 vssd1 vccd1 vccd1 _25536_/D sky130_fd_sc_hd__nor3_1
XFILLER_159_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14564_ _15615_/S _18059_/B _17810_/B vssd1 vssd1 vccd1 vccd1 _14564_/X sky130_fd_sc_hd__and3_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _25822_/Q _16384_/S _15263_/S _16302_/X vssd1 vssd1 vccd1 vccd1 _16303_/X
+ sky130_fd_sc_hd__o211a_1
X_13515_ _14375_/S vssd1 vssd1 vccd1 vccd1 _14365_/S sky130_fd_sc_hd__buf_2
XFILLER_201_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17283_ _17283_/A _17283_/B _17284_/B vssd1 vssd1 vccd1 vccd1 _25515_/D sky130_fd_sc_hd__nor3_1
X_14495_ _14495_/A vssd1 vssd1 vccd1 vccd1 _15979_/S sky130_fd_sc_hd__buf_4
X_19022_ _27087_/Q _18815_/X _18816_/X _27185_/Q _18817_/X vssd1 vssd1 vccd1 vccd1
+ _19022_/X sky130_fd_sc_hd__a221o_1
XFILLER_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16234_ _14859_/X _16231_/X _16233_/X _15020_/X vssd1 vssd1 vccd1 vccd1 _16234_/X
+ sky130_fd_sc_hd__a211o_1
X_13446_ _25839_/Q _26039_/Q _13616_/S vssd1 vssd1 vccd1 vccd1 _13446_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16165_ _15044_/A _16163_/X _16164_/X _12703_/A _15647_/S vssd1 vssd1 vccd1 vccd1
+ _16165_/X sky130_fd_sc_hd__o2111a_1
XFILLER_127_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13377_ _17809_/A vssd1 vssd1 vccd1 vccd1 _15615_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15116_ _14764_/A _15114_/X _15115_/X _14759_/A vssd1 vssd1 vccd1 vccd1 _15117_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16096_ _16104_/A _16096_/B vssd1 vssd1 vccd1 vccd1 _16096_/X sky130_fd_sc_hd__or2_1
XFILLER_114_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19924_ _19976_/C _19923_/Y _19980_/C vssd1 vssd1 vccd1 vccd1 _19925_/B sky130_fd_sc_hd__a21bo_1
X_15047_ _16325_/S vssd1 vssd1 vccd1 vccd1 _16377_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_141_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19855_ _19855_/A _19829_/A vssd1 vssd1 vccd1 vccd1 _19855_/X sky130_fd_sc_hd__or2b_1
XFILLER_123_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18806_ _18806_/A vssd1 vssd1 vccd1 vccd1 _18806_/X sky130_fd_sc_hd__buf_2
XFILLER_228_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19786_ _20000_/A vssd1 vssd1 vccd1 vccd1 _19787_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_284_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16998_ _22487_/A _16996_/X _16990_/A _18541_/A vssd1 vssd1 vccd1 vccd1 _16998_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_110_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18737_ _18597_/X _18731_/Y _18732_/Y _18602_/X _18736_/X vssd1 vssd1 vccd1 vccd1
+ _18737_/X sky130_fd_sc_hd__o221a_1
XFILLER_83_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15949_ _16585_/A _20008_/A _15948_/Y vssd1 vssd1 vccd1 vccd1 _16037_/A sky130_fd_sc_hd__a21oi_4
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18668_ _18891_/A _18651_/Y _18665_/X _18667_/X _18005_/A vssd1 vssd1 vccd1 vccd1
+ _18668_/X sky130_fd_sc_hd__a221o_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17619_ _17633_/A _17619_/B vssd1 vssd1 vccd1 vccd1 _25586_/D sky130_fd_sc_hd__nor2_1
X_18599_ _18599_/A vssd1 vssd1 vccd1 vccd1 _18599_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_53_wb_clk_i clkbuf_leaf_53_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _27278_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_196_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20630_ _20630_/A _20630_/B vssd1 vssd1 vccd1 vccd1 _20630_/X sky130_fd_sc_hd__or2_1
XFILLER_149_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20561_ _20561_/A vssd1 vssd1 vccd1 vccd1 _25708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22300_ _22630_/B vssd1 vssd1 vccd1 vccd1 _22300_/X sky130_fd_sc_hd__clkbuf_2
X_20492_ _20622_/S vssd1 vssd1 vccd1 vccd1 _20509_/S sky130_fd_sc_hd__buf_2
X_23280_ _23280_/A vssd1 vssd1 vccd1 vccd1 _26582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22231_ _26192_/Q input188/X _22231_/S vssd1 vssd1 vccd1 vccd1 _22231_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22162_ _26172_/Q _22152_/X _22161_/X _22148_/X vssd1 vssd1 vccd1 vccd1 _26172_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_279_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21113_ _21113_/A vssd1 vssd1 vccd1 vccd1 _21113_/X sky130_fd_sc_hd__clkbuf_2
X_26970_ _27001_/CLK _26970_/D vssd1 vssd1 vccd1 vccd1 _26970_/Q sky130_fd_sc_hd__dfxtp_1
X_22093_ _26154_/Q _20955_/X _22099_/S vssd1 vssd1 vccd1 vccd1 _22094_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21044_ _25891_/Q _20942_/X _21048_/S vssd1 vssd1 vccd1 vccd1 _21045_/A sky130_fd_sc_hd__mux2_1
X_25921_ _27087_/CLK _25921_/D vssd1 vssd1 vccd1 vccd1 _25921_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_86_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25852_ _27329_/A _25852_/D vssd1 vssd1 vccd1 vccd1 _25852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24803_ _27106_/Q _24818_/B vssd1 vssd1 vccd1 vccd1 _24803_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25783_ _27324_/CLK _25783_/D vssd1 vssd1 vccd1 vccd1 _25783_/Q sky130_fd_sc_hd__dfxtp_1
X_22995_ _26470_/Q _22688_/X _22995_/S vssd1 vssd1 vccd1 vccd1 _22996_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24734_ _24742_/A _24734_/B vssd1 vssd1 vccd1 vccd1 _27090_/D sky130_fd_sc_hd__nor2_1
XFILLER_55_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21946_ _21946_/A vssd1 vssd1 vccd1 vccd1 _21955_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_243_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24665_ _27074_/Q _24657_/X _24664_/Y _24660_/X vssd1 vssd1 vccd1 vccd1 _24666_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_21877_ _26062_/Q _21885_/B vssd1 vssd1 vccd1 vccd1 _21877_/X sky130_fd_sc_hd__or2_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26404_ _26468_/CLK _26404_/D vssd1 vssd1 vccd1 vccd1 _26404_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_199_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23616_ _23616_/A vssd1 vssd1 vccd1 vccd1 _26716_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20828_ _25810_/Q vssd1 vssd1 vccd1 vccd1 _20829_/A sky130_fd_sc_hd__clkbuf_1
X_24596_ _27054_/Q _24589_/X _24595_/Y _24593_/X vssd1 vssd1 vccd1 vccd1 _27054_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_196_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26335_ _26433_/CLK _26335_/D vssd1 vssd1 vccd1 vccd1 _26335_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_168_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23547_ _26695_/Q _23546_/X _23556_/S vssd1 vssd1 vccd1 vccd1 _23548_/A sky130_fd_sc_hd__mux2_1
X_20759_ _20567_/X _25776_/Q _20761_/S vssd1 vssd1 vccd1 vccd1 _20760_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13300_ _15321_/A _26339_/Q _26599_/Q _16267_/S _13321_/A vssd1 vssd1 vccd1 vccd1
+ _13300_/X sky130_fd_sc_hd__a221o_1
XFILLER_155_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14280_ _13173_/A _14279_/X _13026_/A vssd1 vssd1 vccd1 vccd1 _14280_/X sky130_fd_sc_hd__o21a_1
X_26266_ _26271_/CLK _26266_/D vssd1 vssd1 vccd1 vccd1 _26266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23478_ _26670_/Q _23095_/X _23480_/S vssd1 vssd1 vccd1 vccd1 _23479_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13231_ _16022_/A vssd1 vssd1 vccd1 vccd1 _13821_/A sky130_fd_sc_hd__buf_2
XFILLER_196_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25217_ _25217_/A vssd1 vssd1 vccd1 vccd1 _25217_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22429_ _26196_/Q _22418_/X _22427_/X _22428_/X vssd1 vssd1 vccd1 vccd1 _26244_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26197_ _26250_/CLK _26197_/D vssd1 vssd1 vccd1 vccd1 _26197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13162_ _13162_/A vssd1 vssd1 vccd1 vccd1 _13163_/A sky130_fd_sc_hd__buf_2
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25148_ _27193_/Q _25137_/X _25146_/X _25147_/Y _22380_/X vssd1 vssd1 vccd1 vccd1
+ _27193_/D sky130_fd_sc_hd__o221a_1
XFILLER_108_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13093_ _15645_/S _13092_/X _13071_/A vssd1 vssd1 vccd1 vccd1 _13093_/X sky130_fd_sc_hd__a21o_1
X_25079_ _25106_/A vssd1 vssd1 vccd1 vccd1 _25079_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17970_ _17978_/B _17978_/C vssd1 vssd1 vccd1 vccd1 _17970_/X sky130_fd_sc_hd__or2_1
XFILLER_46_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16921_ _16921_/A _16927_/B vssd1 vssd1 vccd1 vccd1 _16973_/C sky130_fd_sc_hd__nor2_1
XFILLER_172_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19640_ _19640_/A _25114_/A _19634_/B vssd1 vssd1 vccd1 vccd1 _24777_/A sky130_fd_sc_hd__or3b_4
X_16852_ _16852_/A _16859_/A vssd1 vssd1 vccd1 vccd1 _16852_/X sky130_fd_sc_hd__and2_2
XFILLER_1_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15803_ _15460_/S _15800_/X _15802_/X _13159_/A vssd1 vssd1 vccd1 vccd1 _15803_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_92_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19571_ _19571_/A _19571_/B _19571_/C _19571_/D vssd1 vssd1 vccd1 vccd1 _19572_/D
+ sky130_fd_sc_hd__or4_1
X_16783_ _16887_/A vssd1 vssd1 vccd1 vccd1 _16834_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13995_ _25835_/Q _26035_/Q _14009_/S vssd1 vssd1 vccd1 vccd1 _13995_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18522_ _25540_/Q _18459_/X _18521_/X _18436_/A _18466_/X vssd1 vssd1 vccd1 vccd1
+ _18522_/X sky130_fd_sc_hd__a221o_1
X_15734_ _26859_/Q _25773_/Q _15734_/S vssd1 vssd1 vccd1 vccd1 _15734_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12946_ _12946_/A vssd1 vssd1 vccd1 vccd1 _13916_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18453_ _27139_/Q _27043_/Q _19334_/B vssd1 vssd1 vccd1 vccd1 _18453_/X sky130_fd_sc_hd__mux2_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15665_ _13267_/X _26700_/Q _26828_/Q _16186_/S _16088_/A vssd1 vssd1 vccd1 vccd1
+ _15665_/X sky130_fd_sc_hd__a221o_1
X_12877_ _25482_/Q vssd1 vssd1 vccd1 vccd1 _21429_/A sky130_fd_sc_hd__buf_2
XFILLER_34_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _25553_/Q vssd1 vssd1 vccd1 vccd1 _17408_/A sky130_fd_sc_hd__clkbuf_2
X_14616_ _14616_/A vssd1 vssd1 vccd1 vccd1 _14617_/A sky130_fd_sc_hd__buf_2
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18384_ _18577_/A vssd1 vssd1 vccd1 vccd1 _19374_/B sky130_fd_sc_hd__clkbuf_2
X_15596_ _26537_/Q _26145_/Q _15596_/S vssd1 vssd1 vccd1 vccd1 _15597_/B sky130_fd_sc_hd__mux2_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _25531_/Q _17333_/B _17334_/Y vssd1 vssd1 vccd1 vccd1 _25531_/D sky130_fd_sc_hd__o21a_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _13520_/A _25758_/Q _14375_/S _26844_/Q _14458_/S vssd1 vssd1 vccd1 vccd1
+ _14547_/X sky130_fd_sc_hd__o221a_1
XFILLER_202_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17266_ _17285_/A _17273_/C vssd1 vssd1 vccd1 vccd1 _17266_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14478_ _14466_/X _14470_/X _14477_/X _13365_/A vssd1 vssd1 vccd1 vccd1 _14478_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16217_ _15044_/X _16215_/X _16216_/X vssd1 vssd1 vccd1 vccd1 _16217_/X sky130_fd_sc_hd__o21a_1
X_19005_ _19448_/A _18975_/Y _19004_/X vssd1 vssd1 vccd1 vccd1 _19005_/Y sky130_fd_sc_hd__o21ai_4
X_13429_ _15961_/B vssd1 vssd1 vccd1 vccd1 _15800_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_128_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17197_ _17197_/A _17224_/B vssd1 vssd1 vccd1 vccd1 _17197_/Y sky130_fd_sc_hd__nand2_1
X_16148_ _16320_/S _16145_/X _16147_/X _15040_/A vssd1 vssd1 vccd1 vccd1 _16148_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_115_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_171_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26264_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_100_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26238_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16079_ _16077_/X _16078_/X _16079_/S vssd1 vssd1 vccd1 vccd1 _16079_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19907_ _25669_/Q _19906_/C _25670_/Q vssd1 vssd1 vccd1 vccd1 _19907_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19838_ _27108_/Q _19722_/X _19761_/X _19837_/Y vssd1 vssd1 vccd1 vccd1 _19838_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput1 coreIndex[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_4
XFILLER_271_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19769_ _19769_/A _19769_/B vssd1 vssd1 vccd1 vccd1 _19769_/X sky130_fd_sc_hd__or2_1
XFILLER_272_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21800_ _21800_/A vssd1 vssd1 vccd1 vccd1 _26030_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22780_ _22802_/A vssd1 vssd1 vccd1 vccd1 _22789_/S sky130_fd_sc_hd__buf_4
XFILLER_225_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21731_ _21731_/A vssd1 vssd1 vccd1 vccd1 _26000_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24450_ _24361_/S _25613_/Q _24449_/X vssd1 vssd1 vccd1 vccd1 _24707_/B sky130_fd_sc_hd__o21a_4
XFILLER_169_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21662_ _25972_/Q input207/X _21662_/S vssd1 vssd1 vccd1 vccd1 _21663_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23401_ _23401_/A vssd1 vssd1 vccd1 vccd1 _26635_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20613_ _23779_/A vssd1 vssd1 vccd1 vccd1 _20613_/X sky130_fd_sc_hd__clkbuf_2
X_24381_ _24472_/A vssd1 vssd1 vccd1 vccd1 _24381_/X sky130_fd_sc_hd__buf_2
X_21593_ input61/X input96/X _21615_/S vssd1 vssd1 vccd1 vccd1 _21594_/A sky130_fd_sc_hd__mux2_8
XFILLER_138_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26120_ _27329_/A _26120_/D vssd1 vssd1 vccd1 vccd1 _26120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23332_ _23332_/A vssd1 vssd1 vccd1 vccd1 _26605_/D sky130_fd_sc_hd__clkbuf_1
X_20544_ _20544_/A vssd1 vssd1 vccd1 vccd1 _25704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26051_ _26611_/CLK _26051_/D vssd1 vssd1 vccd1 vccd1 _26051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23263_ _23263_/A vssd1 vssd1 vccd1 vccd1 _26574_/D sky130_fd_sc_hd__clkbuf_1
X_20475_ _20465_/Y _20707_/D _20712_/A _20474_/X vssd1 vssd1 vccd1 vccd1 _20475_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_117_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25002_ _25113_/A vssd1 vssd1 vccd1 vccd1 _25138_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_22214_ input5/X input280/X _22226_/S vssd1 vssd1 vccd1 vccd1 _22214_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23194_ _26544_/Q _23114_/X _23194_/S vssd1 vssd1 vccd1 vccd1 _23195_/A sky130_fd_sc_hd__mux2_1
X_22145_ _22210_/A vssd1 vssd1 vccd1 vccd1 _22207_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_279_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput360 _16825_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[4] sky130_fd_sc_hd__buf_2
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput371 _12671_/Y vssd1 vssd1 vccd1 vccd1 core_wb_we_o sky130_fd_sc_hd__buf_2
Xoutput382 _17029_/X vssd1 vssd1 vccd1 vccd1 din0[15] sky130_fd_sc_hd__buf_2
XFILLER_117_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26953_ _26987_/CLK _26953_/D vssd1 vssd1 vccd1 vccd1 _26953_/Q sky130_fd_sc_hd__dfxtp_1
X_22076_ _22076_/A vssd1 vssd1 vccd1 vccd1 _26146_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput393 _17043_/X vssd1 vssd1 vccd1 vccd1 din0[25] sky130_fd_sc_hd__buf_2
XFILLER_273_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21027_ _21027_/A vssd1 vssd1 vccd1 vccd1 _25883_/D sky130_fd_sc_hd__clkbuf_1
X_25904_ _26278_/CLK _25904_/D vssd1 vssd1 vccd1 vccd1 _25904_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26884_ _26916_/CLK _26884_/D vssd1 vssd1 vccd1 vccd1 _26884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25835_ _26462_/CLK _25835_/D vssd1 vssd1 vccd1 vccd1 _25835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_267_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12800_ _17971_/C _18194_/B _12810_/A _17971_/B vssd1 vssd1 vccd1 vccd1 _18001_/A
+ sky130_fd_sc_hd__a211oi_4
X_25766_ _27276_/CLK _25766_/D vssd1 vssd1 vccd1 vccd1 _25766_/Q sky130_fd_sc_hd__dfxtp_2
X_13780_ _26788_/Q _26432_/Q _16110_/S vssd1 vssd1 vccd1 vccd1 _13780_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22978_ _26462_/Q _22663_/X _22984_/S vssd1 vssd1 vccd1 vccd1 _22979_/A sky130_fd_sc_hd__mux2_1
XFILLER_250_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12731_ _12731_/A vssd1 vssd1 vccd1 vccd1 _13943_/A sky130_fd_sc_hd__buf_2
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24717_ _24722_/A _24717_/B vssd1 vssd1 vccd1 vccd1 _27086_/D sky130_fd_sc_hd__nor2_1
XFILLER_215_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21929_ _20563_/X _26081_/Q _21933_/S vssd1 vssd1 vccd1 vccd1 _21930_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25697_ _26593_/CLK _25697_/D vssd1 vssd1 vccd1 vccd1 _25697_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15450_ _13694_/A _26702_/Q _26830_/Q _15464_/B vssd1 vssd1 vccd1 vccd1 _15450_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24648_ _24706_/A vssd1 vssd1 vccd1 vccd1 _24739_/A sky130_fd_sc_hd__buf_4
XFILLER_203_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14401_ _14401_/A _14401_/B vssd1 vssd1 vccd1 vccd1 _14594_/A sky130_fd_sc_hd__nor2_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15381_ _15044_/A _15380_/X _13703_/A vssd1 vssd1 vccd1 vccd1 _15381_/X sky130_fd_sc_hd__a21o_1
XFILLER_212_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24579_ _24936_/A _24582_/B vssd1 vssd1 vccd1 vccd1 _24579_/Y sky130_fd_sc_hd__nand2_1
XFILLER_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17120_ _22377_/A vssd1 vssd1 vccd1 vccd1 _17120_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26318_ _26326_/CLK _26318_/D vssd1 vssd1 vccd1 vccd1 _26318_/Q sky130_fd_sc_hd__dfxtp_2
X_14332_ _25799_/Q _27233_/Q _14332_/S vssd1 vssd1 vccd1 vccd1 _14332_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27298_ _27298_/CLK _27298_/D vssd1 vssd1 vccd1 vccd1 _27298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17051_ _17063_/A vssd1 vssd1 vccd1 vccd1 _17051_/X sky130_fd_sc_hd__buf_2
X_14263_ _25832_/Q _26032_/Q _14263_/S vssd1 vssd1 vccd1 vccd1 _14263_/X sky130_fd_sc_hd__mux2_1
X_26249_ _26250_/CLK _26249_/D vssd1 vssd1 vccd1 vccd1 _26249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16002_ _13835_/X _26888_/Q _26760_/Q _13534_/S _13814_/X vssd1 vssd1 vccd1 vccd1
+ _16002_/X sky130_fd_sc_hd__a221o_1
X_13214_ _13214_/A vssd1 vssd1 vccd1 vccd1 _15127_/A sky130_fd_sc_hd__buf_6
XFILLER_125_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14194_ _16031_/S vssd1 vssd1 vccd1 vccd1 _16585_/A sky130_fd_sc_hd__buf_4
XFILLER_100_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13145_ _14870_/A _13130_/X _13138_/X _14659_/A vssd1 vssd1 vccd1 vccd1 _13145_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13076_ _15972_/B vssd1 vssd1 vccd1 vccd1 _15984_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _16043_/B _16040_/B _17957_/S vssd1 vssd1 vccd1 vccd1 _17953_/X sky130_fd_sc_hd__mux2_1
XFILLER_257_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16904_ _16924_/A _16904_/B vssd1 vssd1 vccd1 vccd1 _16905_/A sky130_fd_sc_hd__and2_1
XFILLER_78_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17884_ _17947_/S vssd1 vssd1 vccd1 vccd1 _17933_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_93_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19623_ _27060_/Q _26061_/Q _19623_/C vssd1 vssd1 vccd1 vccd1 _19623_/X sky130_fd_sc_hd__and3_1
XFILLER_238_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16835_ _16835_/A vssd1 vssd1 vccd1 vccd1 _16835_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_226_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19554_ _20657_/A vssd1 vssd1 vccd1 vccd1 _20644_/A sky130_fd_sc_hd__buf_8
XFILLER_20_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13978_ _13305_/A _13947_/X _13954_/X _13509_/A _13977_/X vssd1 vssd1 vccd1 vccd1
+ _13978_/X sky130_fd_sc_hd__a311o_4
XFILLER_202_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16766_ _25682_/Q vssd1 vssd1 vccd1 vccd1 _22518_/A sky130_fd_sc_hd__buf_2
XFILLER_202_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18505_ _18949_/B vssd1 vssd1 vccd1 vccd1 _19258_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_19_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15717_ _26795_/Q _26439_/Q _15726_/S vssd1 vssd1 vccd1 vccd1 _15717_/X sky130_fd_sc_hd__mux2_1
X_12929_ _12929_/A vssd1 vssd1 vccd1 vccd1 _12929_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19485_ _19552_/A vssd1 vssd1 vccd1 vccd1 _19568_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16697_ _17055_/A _17055_/B _19385_/B _16697_/D vssd1 vssd1 vccd1 vccd1 _21709_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_207_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18436_ _18436_/A vssd1 vssd1 vccd1 vccd1 _18437_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15648_ _25708_/Q _16073_/B vssd1 vssd1 vccd1 vccd1 _15648_/X sky130_fd_sc_hd__or2_1
XFILLER_222_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15579_ _15331_/A _26893_/Q _26765_/Q _16193_/S _13284_/A vssd1 vssd1 vccd1 vccd1
+ _15579_/X sky130_fd_sc_hd__a221o_1
X_18367_ _18603_/A vssd1 vssd1 vccd1 vccd1 _18368_/A sky130_fd_sc_hd__buf_2
XFILLER_147_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17318_ _17414_/A vssd1 vssd1 vccd1 vccd1 _17318_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_193_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18298_ _27041_/Q _18811_/A _18295_/X _18297_/X _18823_/A vssd1 vssd1 vccd1 vccd1
+ _18298_/X sky130_fd_sc_hd__o221a_2
X_17249_ _25505_/Q _17253_/C vssd1 vssd1 vccd1 vccd1 _17252_/A sky130_fd_sc_hd__and2_1
XFILLER_135_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20260_ _20305_/A _20260_/B _20305_/B vssd1 vssd1 vccd1 vccd1 _20261_/B sky130_fd_sc_hd__nor3_1
XFILLER_115_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20191_ _20299_/A vssd1 vssd1 vccd1 vccd1 _20379_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23950_ _26851_/Q _23533_/X _23954_/S vssd1 vssd1 vccd1 vccd1 _23951_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22901_ _26428_/Q _22656_/X _22901_/S vssd1 vssd1 vccd1 vccd1 _22902_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23881_ _23881_/A vssd1 vssd1 vccd1 vccd1 _26820_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25620_ _25624_/CLK _25620_/D vssd1 vssd1 vccd1 vccd1 _25620_/Q sky130_fd_sc_hd__dfxtp_4
X_22832_ _26397_/Q _22659_/X _22840_/S vssd1 vssd1 vccd1 vccd1 _22833_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25551_ _27000_/CLK _25551_/D vssd1 vssd1 vccd1 vccd1 _25551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22763_ _26367_/Q _22666_/X _22767_/S vssd1 vssd1 vccd1 vccd1 _22764_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24502_ _26317_/Q _21869_/X _21871_/X input231/X _24501_/X vssd1 vssd1 vccd1 vccd1
+ _24502_/X sky130_fd_sc_hd__a221o_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21714_ _21714_/A vssd1 vssd1 vccd1 vccd1 _25995_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25482_ _26684_/CLK _25482_/D vssd1 vssd1 vccd1 vccd1 _25482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22694_ _22694_/A vssd1 vssd1 vccd1 vccd1 _26343_/D sky130_fd_sc_hd__clkbuf_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27221_ _27221_/CLK _27221_/D vssd1 vssd1 vccd1 vccd1 _27221_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24433_ _24693_/B vssd1 vssd1 vccd1 vccd1 _24582_/A sky130_fd_sc_hd__clkinv_2
XFILLER_169_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21645_ _21276_/A _21644_/X _21603_/X vssd1 vssd1 vccd1 vccd1 _21645_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27152_ _27156_/CLK _27152_/D vssd1 vssd1 vccd1 vccd1 _27152_/Q sky130_fd_sc_hd__dfxtp_4
X_24364_ _27005_/Q _24357_/X _24363_/Y _22468_/X vssd1 vssd1 vccd1 vccd1 _27005_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21576_ _21574_/X _21575_/X _21512_/X vssd1 vssd1 vccd1 vccd1 _21576_/X sky130_fd_sc_hd__a21o_1
XFILLER_193_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26103_ _26465_/CLK _26103_/D vssd1 vssd1 vccd1 vccd1 _26103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23315_ _23361_/S vssd1 vssd1 vccd1 vccd1 _23324_/S sky130_fd_sc_hd__buf_2
XFILLER_20_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20527_ _20527_/A vssd1 vssd1 vccd1 vccd1 _25700_/D sky130_fd_sc_hd__clkbuf_1
X_27083_ _27087_/CLK _27083_/D vssd1 vssd1 vccd1 vccd1 _27083_/Q sky130_fd_sc_hd__dfxtp_1
X_24295_ _26989_/Q _24295_/B vssd1 vssd1 vccd1 vccd1 _24301_/C sky130_fd_sc_hd__and2_1
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26034_ _26593_/CLK _26034_/D vssd1 vssd1 vccd1 vccd1 _26034_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23246_ _23268_/A vssd1 vssd1 vccd1 vccd1 _23255_/S sky130_fd_sc_hd__buf_4
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20458_ _27162_/Q _20434_/B _20435_/Y vssd1 vssd1 vccd1 vccd1 _20458_/X sky130_fd_sc_hd__a21o_1
XFILLER_4_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23177_ _26536_/Q _23089_/X _23183_/S vssd1 vssd1 vccd1 vccd1 _23178_/A sky130_fd_sc_hd__mux2_1
X_20389_ _20389_/A _20389_/B vssd1 vssd1 vccd1 vccd1 _20391_/A sky130_fd_sc_hd__nand2_1
XFILLER_279_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22128_ _26162_/Q _22110_/X _22127_/X _21878_/X vssd1 vssd1 vccd1 vccd1 _26162_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14950_ _25857_/Q _26057_/Q _14953_/S vssd1 vssd1 vccd1 vccd1 _14950_/X sky130_fd_sc_hd__mux2_1
X_22059_ _22059_/A vssd1 vssd1 vccd1 vccd1 _26138_/D sky130_fd_sc_hd__clkbuf_1
X_26936_ _27259_/CLK _26936_/D vssd1 vssd1 vccd1 vccd1 _26936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13901_ _13877_/X _13900_/X _13173_/A vssd1 vssd1 vccd1 vccd1 _13901_/X sky130_fd_sc_hd__a21o_2
XTAP_5888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14881_ _14881_/A _14881_/B vssd1 vssd1 vccd1 vccd1 _14881_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26867_ _26931_/CLK _26867_/D vssd1 vssd1 vccd1 vccd1 _26867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13832_ _13832_/A vssd1 vssd1 vccd1 vccd1 _15311_/A sky130_fd_sc_hd__buf_2
X_16620_ _17838_/A _16620_/B vssd1 vssd1 vccd1 vccd1 _16621_/A sky130_fd_sc_hd__and2_1
X_25818_ _26744_/CLK _25818_/D vssd1 vssd1 vccd1 vccd1 _25818_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_235_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26798_ _27313_/CLK _26798_/D vssd1 vssd1 vccd1 vccd1 _26798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_207 _20701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16551_ _17857_/A _16551_/B vssd1 vssd1 vccd1 vccd1 _19452_/A sky130_fd_sc_hd__nor2_4
X_13763_ _26496_/Q _26368_/Q _13792_/S vssd1 vssd1 vccd1 vccd1 _13763_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_218 _23562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25749_ _26292_/CLK _25749_/D vssd1 vssd1 vccd1 vccd1 _25749_/Q sky130_fd_sc_hd__dfxtp_4
XINSDIODE2_229 _19971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ _15491_/X _26346_/Q _26606_/Q _15850_/S _15852_/A vssd1 vssd1 vccd1 vccd1
+ _15502_/X sky130_fd_sc_hd__a221o_1
XFILLER_189_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12714_ _16072_/S vssd1 vssd1 vccd1 vccd1 _16328_/A sky130_fd_sc_hd__buf_4
XFILLER_280_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19270_ _18474_/A _19268_/Y _17774_/X vssd1 vssd1 vccd1 vccd1 _19271_/C sky130_fd_sc_hd__o21a_1
X_16482_ _26651_/Q _26747_/Q _16490_/B vssd1 vssd1 vccd1 vccd1 _16482_/X sky130_fd_sc_hd__mux2_1
X_13694_ _13694_/A vssd1 vssd1 vccd1 vccd1 _15063_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18221_ _19078_/A _18151_/Y _18181_/X _18219_/Y _18220_/X vssd1 vssd1 vccd1 vccd1
+ _18221_/X sky130_fd_sc_hd__a32o_1
X_15433_ _16281_/S _23574_/A _15432_/Y _16282_/A vssd1 vssd1 vccd1 vccd1 _19100_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15364_ _15362_/X _15363_/X _16144_/S vssd1 vssd1 vccd1 vccd1 _15364_/X sky130_fd_sc_hd__mux2_1
X_18152_ _18554_/A vssd1 vssd1 vccd1 vccd1 _18741_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_178_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14315_ _13305_/A _14292_/X _14299_/X _13509_/A _14314_/X vssd1 vssd1 vccd1 vccd1
+ _14315_/X sky130_fd_sc_hd__a311o_2
X_17103_ _22515_/A vssd1 vssd1 vccd1 vccd1 _17137_/A sky130_fd_sc_hd__buf_8
XFILLER_183_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18083_ _18349_/S _18413_/A _17984_/Y vssd1 vssd1 vccd1 vccd1 _18859_/B sky130_fd_sc_hd__a21o_1
X_15295_ _26674_/Q _25714_/Q _15414_/A vssd1 vssd1 vccd1 vccd1 _15295_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17034_ _17028_/X _16914_/B _17032_/X input225/X vssd1 vssd1 vccd1 vccd1 _17034_/X
+ sky130_fd_sc_hd__a22o_4
X_14246_ _14244_/X _14245_/X _14246_/S vssd1 vssd1 vccd1 vccd1 _14246_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14177_ _27267_/Q _26460_/Q _14433_/S vssd1 vssd1 vccd1 vccd1 _14177_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_4_0_wb_clk_i INSDIODE2_273/DIODE vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_113_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13128_ _15031_/A _13117_/X _13120_/X _14647_/A vssd1 vssd1 vccd1 vccd1 _13128_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18985_ _25518_/Q _18743_/X _18744_/X _17395_/X vssd1 vssd1 vccd1 vccd1 _18985_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13059_ _15797_/B vssd1 vssd1 vccd1 vccd1 _15474_/S sky130_fd_sc_hd__buf_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17936_ _14570_/B _17780_/B _17949_/S vssd1 vssd1 vccd1 vccd1 _17936_/X sky130_fd_sc_hd__mux2_1
XFILLER_280_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17867_ _17956_/S vssd1 vssd1 vccd1 vccd1 _17957_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_281_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19606_ _19607_/A _19607_/B vssd1 vssd1 vccd1 vccd1 _19606_/Y sky130_fd_sc_hd__nand2_1
X_16818_ _16828_/A _16824_/B _16818_/C vssd1 vssd1 vccd1 vccd1 _16819_/A sky130_fd_sc_hd__and3_4
XFILLER_253_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17798_ _17798_/A _14022_/A vssd1 vssd1 vccd1 vccd1 _17798_/X sky130_fd_sc_hd__or2b_1
XFILLER_235_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19537_ _19525_/X _19072_/X _19536_/X _19528_/X vssd1 vssd1 vccd1 vccd1 _25649_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_207_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16749_ _22502_/A _16742_/X _16743_/X _18932_/B vssd1 vssd1 vccd1 vccd1 _16749_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_235_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19468_ _26972_/Q _18764_/X _18765_/X _27004_/Q vssd1 vssd1 vccd1 vccd1 _19468_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18419_ _18683_/A _18419_/B vssd1 vssd1 vccd1 vccd1 _18419_/X sky130_fd_sc_hd__or2_1
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19399_ _27098_/Q _19058_/X _19059_/X _27196_/Q _19060_/X vssd1 vssd1 vccd1 vccd1
+ _19399_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21430_ _21586_/A vssd1 vssd1 vccd1 vccd1 _21430_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_194_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21361_ _25944_/Q _21310_/X _21360_/Y _21330_/X vssd1 vssd1 vccd1 vccd1 _25944_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_190_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23100_ _23100_/A vssd1 vssd1 vccd1 vccd1 _26507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20312_ _20351_/A _20352_/A vssd1 vssd1 vccd1 vccd1 _20313_/B sky130_fd_sc_hd__and2b_1
X_24080_ _24080_/A vssd1 vssd1 vccd1 vccd1 _26908_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput70 dout0[34] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_1
X_21292_ _20630_/A _21278_/X _21279_/X _21291_/X vssd1 vssd1 vccd1 vccd1 _21292_/X
+ sky130_fd_sc_hd__o211a_1
Xinput81 dout0[44] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput92 dout0[54] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__clkbuf_1
X_23031_ _23031_/A vssd1 vssd1 vccd1 vccd1 _26486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20243_ _20240_/Y _20241_/X _20218_/A _20218_/Y vssd1 vssd1 vccd1 vccd1 _20243_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_107_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20174_ _20174_/A _20174_/B _20200_/B vssd1 vssd1 vccd1 vccd1 _20174_/X sky130_fd_sc_hd__or3_1
XFILLER_89_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24982_ _24627_/A _24902_/A _24966_/X vssd1 vssd1 vccd1 vccd1 _24982_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26721_ _26913_/CLK _26721_/D vssd1 vssd1 vccd1 vccd1 _26721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23933_ _23989_/A vssd1 vssd1 vccd1 vccd1 _24002_/S sky130_fd_sc_hd__clkbuf_8
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26652_ _27295_/CLK _26652_/D vssd1 vssd1 vccd1 vccd1 _26652_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23864_ _23864_/A vssd1 vssd1 vccd1 vccd1 _26812_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_8_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27316_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_25603_ _25607_/CLK _25603_/D vssd1 vssd1 vccd1 vccd1 _25603_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_272_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22815_ _26391_/Q _22742_/X _22815_/S vssd1 vssd1 vccd1 vccd1 _22816_/A sky130_fd_sc_hd__mux2_1
X_26583_ _26939_/CLK _26583_/D vssd1 vssd1 vccd1 vccd1 _26583_/Q sky130_fd_sc_hd__dfxtp_1
X_23795_ _23693_/X _26782_/Q _23799_/S vssd1 vssd1 vccd1 vccd1 _23796_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25534_ _25545_/CLK _25534_/D vssd1 vssd1 vccd1 vccd1 _25534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22746_ _22802_/A vssd1 vssd1 vccd1 vccd1 _22815_/S sky130_fd_sc_hd__buf_6
XFILLER_73_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25465_ _27327_/Q _17224_/A _25465_/S vssd1 vssd1 vccd1 vccd1 _25466_/B sky130_fd_sc_hd__mux2_1
X_22677_ _26338_/Q _22675_/X _22689_/S vssd1 vssd1 vccd1 vccd1 _22678_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27204_ _27230_/CLK _27204_/D vssd1 vssd1 vccd1 vccd1 _27204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24416_ _27013_/Q _24391_/X _24414_/Y _24415_/X vssd1 vssd1 vccd1 vccd1 _27013_/D
+ sky130_fd_sc_hd__o211a_1
X_21628_ _21624_/Y _21627_/X _21202_/A vssd1 vssd1 vccd1 vccd1 _21628_/Y sky130_fd_sc_hd__a21oi_4
X_25396_ _23684_/X _27295_/Q _25404_/S vssd1 vssd1 vccd1 vccd1 _25397_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27135_ _27137_/CLK _27135_/D vssd1 vssd1 vccd1 vccd1 _27135_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24347_ _24347_/A _24347_/B _24347_/C _24346_/X vssd1 vssd1 vccd1 vccd1 _24542_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_201_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21559_ _25492_/Q _21559_/B vssd1 vssd1 vccd1 vccd1 _21559_/X sky130_fd_sc_hd__or2_1
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14100_ _14100_/A vssd1 vssd1 vccd1 vccd1 _14421_/A sky130_fd_sc_hd__buf_2
XFILLER_181_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27066_ _27160_/CLK _27066_/D vssd1 vssd1 vccd1 vccd1 _27066_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_4_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15080_ _16250_/A _15079_/X _14718_/X vssd1 vssd1 vccd1 vccd1 _15080_/Y sky130_fd_sc_hd__o21ai_2
X_24278_ _26983_/Q _24278_/B vssd1 vssd1 vccd1 vccd1 _24284_/C sky130_fd_sc_hd__and2_1
X_14031_ _14031_/A _14031_/B vssd1 vssd1 vccd1 vccd1 _14032_/B sky130_fd_sc_hd__nor2_2
XFILLER_141_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26017_ _27283_/CLK _26017_/D vssd1 vssd1 vccd1 vccd1 _26017_/Q sky130_fd_sc_hd__dfxtp_1
X_23229_ _26559_/Q _23060_/X _23233_/S vssd1 vssd1 vccd1 vccd1 _23230_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18770_ _18832_/A vssd1 vssd1 vccd1 vccd1 _18770_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15982_ _15980_/X _15981_/X _15982_/S vssd1 vssd1 vccd1 vccd1 _15982_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17721_ _18161_/A _17728_/B vssd1 vssd1 vccd1 vccd1 _17762_/C sky130_fd_sc_hd__or2_2
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26919_ _27306_/CLK _26919_/D vssd1 vssd1 vccd1 vccd1 _26919_/Q sky130_fd_sc_hd__dfxtp_1
X_14933_ _16458_/B vssd1 vssd1 vccd1 vccd1 _17852_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_94_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ _24723_/A vssd1 vssd1 vccd1 vccd1 _21709_/A sky130_fd_sc_hd__buf_4
XFILLER_264_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14864_ _17197_/A _14848_/X _14852_/X _14863_/X _14683_/X vssd1 vssd1 vccd1 vccd1
+ _14864_/X sky130_fd_sc_hd__a311o_1
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16603_ _16833_/A _16603_/B vssd1 vssd1 vccd1 vccd1 _16697_/D sky130_fd_sc_hd__nand2_4
X_13815_ _13813_/X _26335_/Q _26595_/Q _13534_/S _13814_/X vssd1 vssd1 vccd1 vccd1
+ _13815_/X sky130_fd_sc_hd__a221o_1
XFILLER_223_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14795_ _27325_/Q _26582_/Q _14811_/S vssd1 vssd1 vccd1 vccd1 _14795_/X sky130_fd_sc_hd__mux2_1
X_17583_ _17595_/A _17583_/B vssd1 vssd1 vccd1 vccd1 _25577_/D sky130_fd_sc_hd__nor2_1
XFILLER_90_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19322_ _19322_/A _19393_/B vssd1 vssd1 vccd1 vccd1 _19322_/Y sky130_fd_sc_hd__nand2_1
X_13746_ input169/X input141/X _14132_/S vssd1 vssd1 vccd1 vccd1 _13747_/B sky130_fd_sc_hd__mux2_8
X_16534_ _25828_/Q _27262_/Q _16541_/S vssd1 vssd1 vccd1 vccd1 _16534_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19253_ _19253_/A vssd1 vssd1 vccd1 vccd1 _19253_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13677_ _13841_/A vssd1 vssd1 vccd1 vccd1 _16014_/S sky130_fd_sc_hd__clkbuf_4
X_16465_ _25661_/Q _24351_/B _13578_/X _25629_/Q vssd1 vssd1 vccd1 vccd1 _16465_/X
+ sky130_fd_sc_hd__a22o_1
X_18204_ _18598_/S vssd1 vssd1 vccd1 vccd1 _18487_/A sky130_fd_sc_hd__clkbuf_2
XPHY_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15416_ _26540_/Q _26148_/Q _16256_/B vssd1 vssd1 vccd1 vccd1 _15417_/B sky130_fd_sc_hd__mux2_1
X_16396_ _26123_/Q _26024_/Q _16396_/S vssd1 vssd1 vccd1 vccd1 _16396_/X sky130_fd_sc_hd__mux2_1
X_19184_ _12722_/B _18890_/X _19182_/Y _19183_/Y _18933_/X vssd1 vssd1 vccd1 vccd1
+ _19184_/X sky130_fd_sc_hd__a221o_2
XPHY_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15347_ _25650_/Q _16212_/B vssd1 vssd1 vccd1 vccd1 _15347_/X sky130_fd_sc_hd__and2_1
XFILLER_8_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18135_ _14480_/X _16517_/X _18577_/A vssd1 vssd1 vccd1 vccd1 _18135_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15278_ _15274_/X _15277_/X _16398_/S vssd1 vssd1 vccd1 vccd1 _15278_/X sky130_fd_sc_hd__mux2_1
X_18066_ _17924_/X _17936_/X _18067_/S vssd1 vssd1 vccd1 vccd1 _18066_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14229_ _14220_/X _14227_/X _14228_/X vssd1 vssd1 vccd1 vccd1 _14229_/X sky130_fd_sc_hd__o21a_1
X_17017_ _17039_/A vssd1 vssd1 vccd1 vccd1 _17017_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_78_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26845_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_160_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18968_ _18968_/A _18968_/B vssd1 vssd1 vccd1 vccd1 _18968_/X sky130_fd_sc_hd__or2_1
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17919_ _18317_/S vssd1 vssd1 vccd1 vccd1 _18729_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18899_ _18899_/A _18936_/B _18936_/C vssd1 vssd1 vccd1 vccd1 _18899_/X sky130_fd_sc_hd__or3_1
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20930_ _25847_/Q _20929_/X _20933_/S vssd1 vssd1 vccd1 vccd1 _20931_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20861_ _20861_/A vssd1 vssd1 vccd1 vccd1 _25826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22600_ _22600_/A vssd1 vssd1 vccd1 vccd1 _22600_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_207_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23580_ _23580_/A vssd1 vssd1 vccd1 vccd1 _26705_/D sky130_fd_sc_hd__clkbuf_1
X_20792_ _22472_/B _20973_/B _20792_/C vssd1 vssd1 vccd1 vccd1 _20793_/A sky130_fd_sc_hd__and3_1
XFILLER_241_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22531_ _22531_/A _22533_/B vssd1 vssd1 vccd1 vccd1 _22532_/A sky130_fd_sc_hd__and2_1
XFILLER_168_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25250_ _25306_/A vssd1 vssd1 vccd1 vccd1 _25319_/S sky130_fd_sc_hd__buf_4
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22462_ _26208_/Q _22459_/X _22461_/X _22455_/X vssd1 vssd1 vccd1 vccd1 _26256_/D
+ sky130_fd_sc_hd__o211a_1
X_24201_ _26957_/Q _24203_/C _24200_/Y vssd1 vssd1 vccd1 vccd1 _26957_/D sky130_fd_sc_hd__o21a_1
XFILLER_210_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21413_ _25948_/Q _21378_/X _21412_/Y _21400_/X vssd1 vssd1 vccd1 vccd1 _25948_/D
+ sky130_fd_sc_hd__a211o_1
X_25181_ _24645_/B _25172_/X _25175_/X _27200_/Q _25179_/X vssd1 vssd1 vccd1 vccd1
+ _27200_/D sky130_fd_sc_hd__o221a_1
X_22393_ _22393_/A vssd1 vssd1 vccd1 vccd1 _22394_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24132_ _24132_/A vssd1 vssd1 vccd1 vccd1 _26932_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21344_ _21507_/A vssd1 vssd1 vccd1 vccd1 _21620_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24063_ _24063_/A vssd1 vssd1 vccd1 vccd1 _26901_/D sky130_fd_sc_hd__clkbuf_1
X_21275_ _21275_/A vssd1 vssd1 vccd1 vccd1 _21276_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23014_ _23014_/A vssd1 vssd1 vccd1 vccd1 _26478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20226_ _25745_/Q vssd1 vssd1 vccd1 vccd1 _20679_/A sky130_fd_sc_hd__buf_8
XFILLER_143_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20157_ _27151_/Q _27085_/Q vssd1 vssd1 vccd1 vccd1 _20159_/A sky130_fd_sc_hd__nor2_1
XFILLER_249_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24965_ _27155_/Q _24953_/X _24964_/Y _24949_/X vssd1 vssd1 vccd1 vccd1 _27155_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20088_ _19981_/A _20081_/X _20086_/Y _20087_/X vssd1 vssd1 vccd1 vccd1 _20205_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_40_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26704_ _27253_/CLK _26704_/D vssd1 vssd1 vccd1 vccd1 _26704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23916_ _23916_/A vssd1 vssd1 vccd1 vccd1 _26836_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24896_ _27132_/Q _24896_/B vssd1 vssd1 vccd1 vccd1 _24896_/Y sky130_fd_sc_hd__nand2_1
XFILLER_246_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26635_ _27313_/CLK _26635_/D vssd1 vssd1 vccd1 vccd1 _26635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23847_ _23847_/A vssd1 vssd1 vccd1 vccd1 _26805_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _14008_/S vssd1 vssd1 vccd1 vccd1 _15805_/S sky130_fd_sc_hd__buf_4
XFILLER_14_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _25688_/Q _16685_/B _14580_/C vssd1 vssd1 vccd1 vccd1 _20798_/B sky130_fd_sc_hd__or3_4
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26566_ _26599_/CLK _26566_/D vssd1 vssd1 vccd1 vccd1 _26566_/Q sky130_fd_sc_hd__dfxtp_1
X_23778_ _23778_/A vssd1 vssd1 vccd1 vccd1 _26776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ _13359_/X _13513_/X _13528_/X _13530_/X vssd1 vssd1 vccd1 vccd1 _13531_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_214_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25517_ _25518_/CLK _25517_/D vssd1 vssd1 vccd1 vccd1 _25517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22729_ _22729_/A vssd1 vssd1 vccd1 vccd1 _26354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26497_ _27304_/CLK _26497_/D vssd1 vssd1 vccd1 vccd1 _26497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16250_ _16250_/A _16932_/A vssd1 vssd1 vccd1 vccd1 _16250_/Y sky130_fd_sc_hd__nor2_1
X_25448_ _23763_/X _27319_/Q _25448_/S vssd1 vssd1 vccd1 vccd1 _25449_/A sky130_fd_sc_hd__mux2_1
X_13462_ _15868_/B vssd1 vssd1 vccd1 vccd1 _15526_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_139_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15201_ _14764_/A _15195_/X _15200_/X vssd1 vssd1 vccd1 vccd1 _15201_/X sky130_fd_sc_hd__o21a_1
X_16181_ _26801_/Q _26445_/Q _16182_/S vssd1 vssd1 vccd1 vccd1 _16181_/X sky130_fd_sc_hd__mux2_1
X_13393_ _15791_/A _14604_/B _15074_/A _13392_/X vssd1 vssd1 vccd1 vccd1 _13393_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_166_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25379_ _27288_/Q _23766_/A _25387_/S vssd1 vssd1 vccd1 vccd1 _25380_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15132_ _19294_/S _15132_/B vssd1 vssd1 vccd1 vccd1 _17846_/A sky130_fd_sc_hd__nor2_1
X_27118_ _27122_/CLK _27118_/D vssd1 vssd1 vccd1 vccd1 _27118_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27049_ _27049_/CLK _27049_/D vssd1 vssd1 vccd1 vccd1 _27049_/Q sky130_fd_sc_hd__dfxtp_1
X_19940_ _22494_/A _19985_/C _19780_/X vssd1 vssd1 vccd1 vccd1 _19940_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15063_ _15063_/A vssd1 vssd1 vccd1 vccd1 _15167_/A sky130_fd_sc_hd__buf_2
XFILLER_153_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14014_ _13431_/A _14011_/X _14013_/X _13863_/A vssd1 vssd1 vccd1 vccd1 _14014_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_4_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19871_ _19642_/X _19869_/X _19870_/X _19651_/X vssd1 vssd1 vccd1 vccd1 _19871_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_136_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18822_ _27018_/Q _18449_/X _18820_/X _18821_/X vssd1 vssd1 vccd1 vccd1 _18822_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_268_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18753_ _18817_/A vssd1 vssd1 vccd1 vccd1 _18753_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15965_ _27243_/Q _15984_/B vssd1 vssd1 vccd1 vccd1 _15965_/X sky130_fd_sc_hd__or2_1
XFILLER_48_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput260 manufacturerID[6] vssd1 vssd1 vccd1 vccd1 input260/X sky130_fd_sc_hd__clkbuf_2
XTAP_5471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput271 partID[1] vssd1 vssd1 vccd1 vccd1 input271/X sky130_fd_sc_hd__clkbuf_1
XFILLER_209_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17704_ _12722_/B _17486_/A _17704_/S vssd1 vssd1 vccd1 vccd1 _17739_/C sky130_fd_sc_hd__mux2_1
Xinput282 versionID[2] vssd1 vssd1 vccd1 vccd1 input282/X sky130_fd_sc_hd__buf_2
XFILLER_264_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14916_ _25826_/Q _27260_/Q _15003_/S vssd1 vssd1 vccd1 vccd1 _14916_/X sky130_fd_sc_hd__mux2_1
X_18684_ _18259_/X _18263_/X _18684_/S vssd1 vssd1 vccd1 vccd1 _18684_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_196_wb_clk_i _26681_/CLK vssd1 vssd1 vccd1 vccd1 _26903_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15896_ _15894_/X _15895_/X _15903_/S vssd1 vssd1 vccd1 vccd1 _15896_/X sky130_fd_sc_hd__mux2_2
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17635_ _17635_/A vssd1 vssd1 vccd1 vccd1 _17635_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_125_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27062_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_24_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14847_ _12776_/A _26421_/Q _14948_/S _14846_/X vssd1 vssd1 vccd1 vccd1 _14847_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17566_ _25573_/Q _17564_/X _17540_/X _17565_/X vssd1 vssd1 vccd1 vccd1 _17567_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_211_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14778_ _14778_/A vssd1 vssd1 vccd1 vccd1 _14779_/A sky130_fd_sc_hd__clkbuf_4
X_19305_ _26967_/Q _18826_/X _18827_/X _26999_/Q vssd1 vssd1 vccd1 vccd1 _19305_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16517_ _16517_/A vssd1 vssd1 vccd1 vccd1 _16517_/X sky130_fd_sc_hd__buf_6
XFILLER_260_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13729_ _13727_/X _13728_/X _15547_/A vssd1 vssd1 vccd1 vccd1 _13729_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17497_ _24350_/S vssd1 vssd1 vccd1 vccd1 _24340_/S sky130_fd_sc_hd__clkbuf_2
X_19236_ _19237_/B _19237_/C _19237_/A vssd1 vssd1 vccd1 vccd1 _19276_/B sky130_fd_sc_hd__a21o_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16448_ _16350_/A _16432_/X _16447_/X vssd1 vssd1 vccd1 vccd1 _16448_/X sky130_fd_sc_hd__a21o_2
XFILLER_9_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19167_ _27027_/Q _18449_/X _19166_/X _18821_/X vssd1 vssd1 vccd1 vccd1 _19167_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_219_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16379_ _27322_/Q _26579_/Q _16384_/S vssd1 vssd1 vccd1 vccd1 _16379_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18118_ _18161_/C vssd1 vssd1 vccd1 vccd1 _18120_/B sky130_fd_sc_hd__clkinv_2
XFILLER_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19098_ _25521_/Q _18444_/A _19095_/X _19097_/X _18469_/A vssd1 vssd1 vccd1 vccd1
+ _19098_/X sky130_fd_sc_hd__o221a_1
XFILLER_172_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18049_ _17903_/X _17898_/X _18062_/S vssd1 vssd1 vccd1 vccd1 _18049_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21060_ _21060_/A vssd1 vssd1 vccd1 vccd1 _25898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20011_ _19661_/X _20009_/X _19771_/X _20656_/A vssd1 vssd1 vccd1 vccd1 _20039_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24750_ _24972_/A vssd1 vssd1 vccd1 vccd1 _24751_/B sky130_fd_sc_hd__clkinv_2
XFILLER_228_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21962_ _22018_/A vssd1 vssd1 vccd1 vccd1 _22031_/S sky130_fd_sc_hd__buf_8
XFILLER_27_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23701_ _23701_/A vssd1 vssd1 vccd1 vccd1 _26752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20913_ _23728_/A vssd1 vssd1 vccd1 vccd1 _20913_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24681_ _24932_/A vssd1 vssd1 vccd1 vccd1 _24682_/B sky130_fd_sc_hd__inv_2
X_21893_ _21893_/A vssd1 vssd1 vccd1 vccd1 _26064_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23632_ _26724_/Q _23536_/X _23634_/S vssd1 vssd1 vccd1 vccd1 _23633_/A sky130_fd_sc_hd__mux2_1
X_26420_ _27291_/CLK _26420_/D vssd1 vssd1 vccd1 vccd1 _26420_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20844_ _25818_/Q vssd1 vssd1 vccd1 vccd1 _20845_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26351_ _26611_/CLK _26351_/D vssd1 vssd1 vccd1 vccd1 _26351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23563_ _26700_/Q _23562_/X _23572_/S vssd1 vssd1 vccd1 vccd1 _23564_/A sky130_fd_sc_hd__mux2_1
X_20775_ _20596_/X _25783_/Q _20783_/S vssd1 vssd1 vccd1 vccd1 _20776_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25302_ _23760_/X _27254_/Q _25304_/S vssd1 vssd1 vccd1 vccd1 _25303_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_390 _17030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22514_ _22514_/A vssd1 vssd1 vccd1 vccd1 _26281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26282_ _26282_/CLK _26282_/D vssd1 vssd1 vccd1 vccd1 _26282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23494_ _26677_/Q _23117_/X _23502_/S vssd1 vssd1 vccd1 vccd1 _23495_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25233_ _27061_/Q _21873_/A input185/X _25214_/X _25178_/A vssd1 vssd1 vccd1 vccd1
+ _25233_/X sky130_fd_sc_hd__a41o_1
X_22445_ _26202_/Q _22432_/X _22444_/X _22442_/X vssd1 vssd1 vccd1 vccd1 _26250_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25164_ _24768_/Y _25124_/X _25163_/Y _17339_/A vssd1 vssd1 vccd1 vccd1 _25164_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_276_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22376_ _17087_/A _26229_/Q _22376_/S vssd1 vssd1 vccd1 vccd1 _22377_/B sky130_fd_sc_hd__mux2_1
XFILLER_159_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24115_ _24115_/A vssd1 vssd1 vccd1 vccd1 _26924_/D sky130_fd_sc_hd__clkbuf_1
X_21327_ input103/X input74/X _21327_/S vssd1 vssd1 vccd1 vccd1 _21327_/X sky130_fd_sc_hd__mux2_8
XFILLER_135_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25095_ _24711_/Y _25070_/X _25094_/Y _25082_/X vssd1 vssd1 vccd1 vccd1 _25095_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_151_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24046_ _26894_/Q _23568_/X _24048_/S vssd1 vssd1 vccd1 vccd1 _24047_/A sky130_fd_sc_hd__mux2_1
X_21258_ _21271_/A _21258_/B vssd1 vssd1 vccd1 vccd1 _21258_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20209_ _22513_/A _20233_/C vssd1 vssd1 vccd1 vccd1 _20209_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21189_ _21189_/A vssd1 vssd1 vccd1 vccd1 _25933_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25997_ _26240_/CLK _25997_/D vssd1 vssd1 vccd1 vccd1 _25997_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ _21320_/A _21300_/A _12962_/C vssd1 vssd1 vccd1 vccd1 _12963_/D sky130_fd_sc_hd__and3_1
X_15750_ _15750_/A vssd1 vssd1 vccd1 vccd1 _23558_/A sky130_fd_sc_hd__buf_6
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_50 _20635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_24948_ _24948_/A _24951_/B vssd1 vssd1 vccd1 vccd1 _24948_/Y sky130_fd_sc_hd__nand2_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_61 _19901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_72 _20681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_83 _23712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ _26650_/Q _26746_/Q _16467_/A vssd1 vssd1 vccd1 vccd1 _14701_/X sky130_fd_sc_hd__mux2_1
XFILLER_261_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_94 _21259_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _12893_/A vssd1 vssd1 vccd1 vccd1 _13561_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15681_ _26536_/Q _26144_/Q _16182_/S vssd1 vssd1 vccd1 vccd1 _15682_/B sky130_fd_sc_hd__mux2_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24879_ _20690_/A _19905_/X _25143_/A _24896_/B vssd1 vssd1 vccd1 vccd1 _24879_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _25558_/Q _17420_/B vssd1 vssd1 vccd1 vccd1 _17427_/C sky130_fd_sc_hd__and2_1
XFILLER_234_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _16305_/A vssd1 vssd1 vccd1 vccd1 _16319_/S sky130_fd_sc_hd__buf_4
X_26618_ _27293_/CLK _26618_/D vssd1 vssd1 vccd1 vccd1 _26618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_260_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _25535_/Q _25536_/Q _17351_/C vssd1 vssd1 vccd1 vccd1 _17353_/B sky130_fd_sc_hd__and3_1
XFILLER_202_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14563_ _14563_/A vssd1 vssd1 vccd1 vccd1 _17810_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26549_ _27291_/CLK _26549_/D vssd1 vssd1 vccd1 vccd1 _26549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16302_ _27256_/Q _16388_/B vssd1 vssd1 vccd1 vccd1 _16302_/X sky130_fd_sc_hd__or2_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ _14054_/A vssd1 vssd1 vccd1 vccd1 _14375_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_9_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17282_ _25514_/Q _25515_/Q _17282_/C vssd1 vssd1 vccd1 vccd1 _17284_/B sky130_fd_sc_hd__and3_1
X_14494_ _14528_/A _14528_/B _13008_/A vssd1 vssd1 vccd1 vccd1 _16809_/B sky130_fd_sc_hd__a21o_4
X_19021_ _27217_/Q _19299_/B vssd1 vssd1 vccd1 vccd1 _19021_/X sky130_fd_sc_hd__and2_1
X_13445_ _26790_/Q _26434_/Q _13589_/S vssd1 vssd1 vccd1 vccd1 _13445_/X sky130_fd_sc_hd__mux2_1
X_16233_ _12775_/A _26415_/Q _15060_/S _16232_/X vssd1 vssd1 vccd1 vccd1 _16233_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_277_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13376_ _16581_/A vssd1 vssd1 vccd1 vccd1 _17809_/A sky130_fd_sc_hd__buf_4
X_16164_ _12773_/A _26897_/Q _26769_/Q _15351_/B _15169_/A vssd1 vssd1 vccd1 vccd1
+ _16164_/X sky130_fd_sc_hd__a221o_1
XFILLER_126_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15115_ _15111_/X _25855_/Q _26055_/Q _15121_/S _14771_/A vssd1 vssd1 vccd1 vccd1
+ _15115_/X sky130_fd_sc_hd__a221o_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16095_ _26507_/Q _26379_/Q _16182_/S vssd1 vssd1 vccd1 vccd1 _16096_/B sky130_fd_sc_hd__mux2_1
XFILLER_141_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19923_ _19923_/A vssd1 vssd1 vccd1 vccd1 _19923_/Y sky130_fd_sc_hd__inv_2
X_15046_ _15255_/A vssd1 vssd1 vccd1 vccd1 _16325_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_272_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19854_ _19777_/A _19804_/X _19808_/A _19830_/C _19805_/X vssd1 vssd1 vccd1 vccd1
+ _19854_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_268_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18805_ _18805_/A vssd1 vssd1 vccd1 vccd1 _19234_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_228_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19785_ _19753_/A _19750_/Y _19752_/B vssd1 vssd1 vccd1 vccd1 _19785_/Y sky130_fd_sc_hd__o21ai_2
X_16997_ _22485_/A _16996_/X _16990_/A _18483_/A vssd1 vssd1 vccd1 vccd1 _16997_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_283_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18736_ _18733_/X _18735_/X _16633_/B vssd1 vssd1 vccd1 vccd1 _18736_/X sky130_fd_sc_hd__a21o_1
XFILLER_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15948_ _25737_/Q _15948_/B vssd1 vssd1 vccd1 vccd1 _15948_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18667_ _18382_/X _18666_/Y _17671_/X vssd1 vssd1 vccd1 vccd1 _18667_/X sky130_fd_sc_hd__o21a_1
X_15879_ _26533_/Q _26141_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _15879_/X sky130_fd_sc_hd__mux2_1
XFILLER_251_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17618_ _17697_/B _17612_/X _17608_/X _17617_/Y vssd1 vssd1 vccd1 vccd1 _17619_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18598_ _18054_/X _18065_/X _18598_/S vssd1 vssd1 vccd1 vccd1 _18599_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17549_ _24277_/A vssd1 vssd1 vccd1 vccd1 _17634_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_260_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20560_ _20559_/X _25708_/Q _20572_/S vssd1 vssd1 vccd1 vccd1 _20561_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19219_ _19219_/A _19252_/B vssd1 vssd1 vccd1 vccd1 _19219_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_93_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26250_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20491_ _20597_/A vssd1 vssd1 vccd1 vccd1 _20622_/S sky130_fd_sc_hd__buf_8
X_22230_ _22337_/A _22230_/B _22230_/C vssd1 vssd1 vccd1 vccd1 _22231_/S sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_22_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26677_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_192_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22161_ _26171_/Q _22154_/X _22160_/X input264/X _22155_/X vssd1 vssd1 vccd1 vccd1
+ _22161_/X sky130_fd_sc_hd__a221o_1
XFILLER_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21112_ _21112_/A vssd1 vssd1 vccd1 vccd1 _21112_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_278_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22092_ _22092_/A vssd1 vssd1 vccd1 vccd1 _26153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21043_ _21043_/A vssd1 vssd1 vccd1 vccd1 _25890_/D sky130_fd_sc_hd__clkbuf_1
X_25920_ _27087_/CLK _25920_/D vssd1 vssd1 vccd1 vccd1 _25920_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_114_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25851_ _26611_/CLK _25851_/D vssd1 vssd1 vccd1 vccd1 _25851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24802_ _24877_/A vssd1 vssd1 vccd1 vccd1 _24818_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22994_ _22994_/A vssd1 vssd1 vccd1 vccd1 _26469_/D sky130_fd_sc_hd__clkbuf_1
X_25782_ _26611_/CLK _25782_/D vssd1 vssd1 vccd1 vccd1 _25782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21945_ _21945_/A vssd1 vssd1 vccd1 vccd1 _26088_/D sky130_fd_sc_hd__clkbuf_1
X_24733_ _27090_/Q _24724_/X _24732_/Y _24720_/X vssd1 vssd1 vccd1 vccd1 _24734_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_199_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24664_ _24682_/A _24664_/B vssd1 vssd1 vccd1 vccd1 _24664_/Y sky130_fd_sc_hd__nand2_2
XFILLER_215_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21876_ _26294_/Q _21869_/X _21871_/X input226/X vssd1 vssd1 vccd1 vccd1 _21876_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26403_ _26467_/CLK _26403_/D vssd1 vssd1 vccd1 vccd1 _26403_/Q sky130_fd_sc_hd__dfxtp_4
X_23615_ _26716_/Q _23508_/X _23623_/S vssd1 vssd1 vccd1 vccd1 _23616_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20827_ _20827_/A vssd1 vssd1 vccd1 vccd1 _25809_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24595_ hold3/A _24595_/B vssd1 vssd1 vccd1 vccd1 _24595_/Y sky130_fd_sc_hd__nand2_1
XFILLER_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26334_ _26462_/CLK _26334_/D vssd1 vssd1 vccd1 vccd1 _26334_/Q sky130_fd_sc_hd__dfxtp_2
X_23546_ _23546_/A vssd1 vssd1 vccd1 vccd1 _23546_/X sky130_fd_sc_hd__clkbuf_2
X_20758_ _20758_/A vssd1 vssd1 vccd1 vccd1 _25775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26265_ _26271_/CLK _26265_/D vssd1 vssd1 vccd1 vccd1 _26265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23477_ _23477_/A vssd1 vssd1 vccd1 vccd1 _26669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20689_ _20689_/A vssd1 vssd1 vccd1 vccd1 _20703_/B sky130_fd_sc_hd__buf_4
XFILLER_149_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13230_ _13773_/A vssd1 vssd1 vccd1 vccd1 _16022_/A sky130_fd_sc_hd__buf_2
X_25216_ _27217_/Q _25204_/X _25207_/X _24719_/B _25215_/X vssd1 vssd1 vccd1 vccd1
+ _27217_/D sky130_fd_sc_hd__o221a_1
X_22428_ _22428_/A vssd1 vssd1 vccd1 vccd1 _22428_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26196_ _26250_/CLK _26196_/D vssd1 vssd1 vccd1 vccd1 _26196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13161_ _14522_/S vssd1 vssd1 vccd1 vccd1 _13162_/A sky130_fd_sc_hd__buf_2
X_25147_ _25147_/A _25151_/B vssd1 vssd1 vccd1 vccd1 _25147_/Y sky130_fd_sc_hd__nand2_1
X_22359_ _22381_/A vssd1 vssd1 vccd1 vccd1 _22360_/C sky130_fd_sc_hd__inv_2
XFILLER_156_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13092_ _13086_/X _26887_/Q _26759_/Q _15653_/S vssd1 vssd1 vccd1 vccd1 _13092_/X
+ sky130_fd_sc_hd__a22o_1
X_25078_ _27180_/Q _25058_/X _25077_/X vssd1 vssd1 vccd1 vccd1 _27180_/D sky130_fd_sc_hd__o21ba_1
X_24029_ _26886_/Q _23542_/X _24037_/S vssd1 vssd1 vccd1 vccd1 _24030_/A sky130_fd_sc_hd__mux2_1
X_16920_ _16920_/A vssd1 vssd1 vccd1 vccd1 _16920_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16851_ _16851_/A vssd1 vssd1 vccd1 vccd1 _16851_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_277_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15802_ _25811_/Q _15474_/S _15806_/S _15801_/X vssd1 vssd1 vccd1 vccd1 _15802_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19570_ _19570_/A _19570_/B _19570_/C _19570_/D vssd1 vssd1 vccd1 vccd1 _19652_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_265_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16782_ _16782_/A vssd1 vssd1 vccd1 vccd1 _16887_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_280_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13994_ _14520_/S vssd1 vssd1 vccd1 vccd1 _14009_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18521_ _26948_/Q _18461_/X _18463_/X _26980_/Q vssd1 vssd1 vccd1 vccd1 _18521_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_280_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15733_ _13135_/A _15730_/X _15732_/X _13126_/A vssd1 vssd1 vccd1 vccd1 _15733_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _12872_/A _12933_/B _12907_/Y _13569_/B _12850_/Y vssd1 vssd1 vccd1 vccd1
+ _12945_/X sky130_fd_sc_hd__a41o_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18452_ _18757_/A vssd1 vssd1 vccd1 vccd1 _19334_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _14791_/A _15661_/X _15663_/X _13242_/X vssd1 vssd1 vccd1 vccd1 _15668_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_234_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12876_ _15954_/A vssd1 vssd1 vccd1 vccd1 _15791_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _25552_/Q _17401_/B _17402_/Y vssd1 vssd1 vccd1 vccd1 _25552_/D sky130_fd_sc_hd__o21a_1
XFILLER_222_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14615_ _14601_/X _14607_/Y _14614_/X vssd1 vssd1 vccd1 vccd1 _14615_/X sky130_fd_sc_hd__o21a_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _18383_/A vssd1 vssd1 vccd1 vccd1 _18666_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15595_ _26797_/Q _26441_/Q _16176_/S vssd1 vssd1 vccd1 vccd1 _15595_/X sky130_fd_sc_hd__mux2_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17334_/A _17341_/C vssd1 vssd1 vccd1 vccd1 _17334_/Y sky130_fd_sc_hd__nor2_1
XFILLER_187_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14546_ _25797_/Q _27231_/Q _14553_/S vssd1 vssd1 vccd1 vccd1 _14546_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17265_ _25510_/Q _17265_/B vssd1 vssd1 vccd1 vccd1 _17273_/C sky130_fd_sc_hd__and2_1
X_14477_ _13309_/B _14473_/X _14476_/X _14076_/A vssd1 vssd1 vccd1 vccd1 _14477_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_197_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19004_ _18976_/X _19001_/X _19002_/Y _19003_/X vssd1 vssd1 vccd1 vccd1 _19004_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16216_ _12774_/A _26899_/Q _26771_/Q _16377_/S _15048_/X vssd1 vssd1 vccd1 vccd1
+ _16216_/X sky130_fd_sc_hd__a221o_1
X_13428_ _14253_/S vssd1 vssd1 vccd1 vccd1 _15961_/B sky130_fd_sc_hd__buf_2
X_17196_ _25491_/Q _17131_/B _17195_/Y _17188_/X vssd1 vssd1 vccd1 vccd1 _25491_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13359_ _13359_/A vssd1 vssd1 vccd1 vccd1 _13359_/X sky130_fd_sc_hd__buf_4
XFILLER_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16147_ _26085_/Q _16319_/S _15031_/A _16146_/X vssd1 vssd1 vccd1 vccd1 _16147_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16078_ _26115_/Q _26016_/Q _16078_/S vssd1 vssd1 vccd1 vccd1 _16078_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19906_ _25670_/Q _25669_/Q _19906_/C vssd1 vssd1 vccd1 vccd1 _19985_/C sky130_fd_sc_hd__and3_1
X_15029_ _26354_/Q _26614_/Q _15030_/S vssd1 vssd1 vccd1 vccd1 _15029_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19837_ _19837_/A _19837_/B vssd1 vssd1 vccd1 vccd1 _19837_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_140_wb_clk_i _25501_/CLK vssd1 vssd1 vccd1 vccd1 _26063_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput2 coreIndex[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_4
X_19768_ _19768_/A _19768_/B vssd1 vssd1 vccd1 vccd1 _19768_/Y sky130_fd_sc_hd__nand2_1
XFILLER_232_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18719_ _18719_/A vssd1 vssd1 vccd1 vccd1 _18719_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_271_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19699_ _20034_/B vssd1 vssd1 vccd1 vccd1 _20252_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_64_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21730_ _20504_/X _26000_/Q _21732_/S vssd1 vssd1 vccd1 vccd1 _21731_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21661_ _21661_/A vssd1 vssd1 vccd1 vccd1 _25971_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23400_ _26635_/Q _23085_/X _23408_/S vssd1 vssd1 vccd1 vccd1 _23401_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20612_ _23603_/A vssd1 vssd1 vccd1 vccd1 _23779_/A sky130_fd_sc_hd__buf_2
X_24380_ _27008_/Q _24357_/X _24378_/Y _24379_/X vssd1 vssd1 vccd1 vccd1 _27008_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_196_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21592_ _21544_/X _21591_/X _21537_/X vssd1 vssd1 vccd1 vccd1 _21592_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23331_ _20563_/X _26605_/Q _23335_/S vssd1 vssd1 vccd1 vccd1 _23332_/A sky130_fd_sc_hd__mux2_1
X_20543_ _20542_/X _25704_/Q _20551_/S vssd1 vssd1 vccd1 vccd1 _20544_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26050_ _27284_/CLK _26050_/D vssd1 vssd1 vccd1 vccd1 _26050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23262_ _26574_/Q _23108_/X _23266_/S vssd1 vssd1 vccd1 vccd1 _23263_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20474_ _19740_/X _20466_/Y _20467_/X _20473_/X _20248_/A vssd1 vssd1 vccd1 vccd1
+ _20474_/X sky130_fd_sc_hd__o311a_1
X_25001_ _25142_/A vssd1 vssd1 vccd1 vccd1 _25137_/A sky130_fd_sc_hd__clkbuf_2
X_22213_ _26187_/Q _22200_/X _22212_/X _22195_/X vssd1 vssd1 vccd1 vccd1 _26187_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23193_ _23193_/A vssd1 vssd1 vccd1 vccd1 _26543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22144_ _26167_/Q _22136_/X _22143_/X _22132_/X vssd1 vssd1 vccd1 vccd1 _26167_/D
+ sky130_fd_sc_hd__o211a_1
Xoutput350 _16944_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[24] sky130_fd_sc_hd__buf_2
XFILLER_273_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput361 _16829_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput372 _16683_/X vssd1 vssd1 vccd1 vccd1 csb0[0] sky130_fd_sc_hd__buf_2
XFILLER_126_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26952_ _26987_/CLK _26952_/D vssd1 vssd1 vccd1 vccd1 _26952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_273_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22075_ _26146_/Q _20929_/X _22077_/S vssd1 vssd1 vccd1 vccd1 _22076_/A sky130_fd_sc_hd__mux2_1
Xoutput383 _17030_/X vssd1 vssd1 vccd1 vccd1 din0[16] sky130_fd_sc_hd__buf_2
XFILLER_248_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput394 _17044_/X vssd1 vssd1 vccd1 vccd1 din0[26] sky130_fd_sc_hd__buf_2
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21026_ _25883_/Q _20916_/X _21026_/S vssd1 vssd1 vccd1 vccd1 _21027_/A sky130_fd_sc_hd__mux2_1
X_25903_ _26278_/CLK _25903_/D vssd1 vssd1 vccd1 vccd1 _25903_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_48_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26883_ _26917_/CLK _26883_/D vssd1 vssd1 vccd1 vccd1 _26883_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_247_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25834_ _27265_/CLK _25834_/D vssd1 vssd1 vccd1 vccd1 _25834_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_274_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22977_ _22977_/A vssd1 vssd1 vccd1 vccd1 _26461_/D sky130_fd_sc_hd__clkbuf_1
X_25765_ _26594_/CLK _25765_/D vssd1 vssd1 vccd1 vccd1 _25765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12730_ _14384_/A vssd1 vssd1 vccd1 vccd1 _12731_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24716_ _27086_/Q _24701_/X _24715_/Y _24697_/X vssd1 vssd1 vccd1 vccd1 _24717_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_21928_ _21928_/A vssd1 vssd1 vccd1 vccd1 _26080_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_6_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_255_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25696_ _26592_/CLK _25696_/D vssd1 vssd1 vccd1 vccd1 _25696_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_203_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21859_ _21859_/A vssd1 vssd1 vccd1 vccd1 _26057_/D sky130_fd_sc_hd__clkbuf_1
X_24647_ _27070_/Q _24636_/X _24646_/Y _24631_/X vssd1 vssd1 vccd1 vccd1 _27070_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_230_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _17941_/A _14562_/B vssd1 vssd1 vccd1 vccd1 _16706_/A sky130_fd_sc_hd__or2_1
XFILLER_169_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15380_ _12773_/A _26896_/Q _26768_/Q _16135_/B vssd1 vssd1 vccd1 vccd1 _15380_/X
+ sky130_fd_sc_hd__a22o_1
X_24578_ _27047_/Q _24576_/X _24577_/Y _24567_/X vssd1 vssd1 vccd1 vccd1 _27047_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_168_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26317_ _26319_/CLK _26317_/D vssd1 vssd1 vccd1 vccd1 _26317_/Q sky130_fd_sc_hd__dfxtp_4
X_14331_ _14331_/A vssd1 vssd1 vccd1 vccd1 _14331_/X sky130_fd_sc_hd__buf_2
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23529_ _23529_/A vssd1 vssd1 vccd1 vccd1 _26689_/D sky130_fd_sc_hd__clkbuf_1
X_27297_ _27297_/CLK _27297_/D vssd1 vssd1 vccd1 vccd1 _27297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14262_ _26783_/Q _26427_/Q _14263_/S vssd1 vssd1 vccd1 vccd1 _14262_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17050_ _16604_/A _16812_/A _16639_/B _16996_/A vssd1 vssd1 vccd1 vccd1 _20790_/C
+ sky130_fd_sc_hd__a31o_2
X_26248_ _26248_/CLK _26248_/D vssd1 vssd1 vccd1 vccd1 _26248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16001_ _13835_/X _26696_/Q _26824_/Q _15514_/S _15999_/A vssd1 vssd1 vccd1 vccd1
+ _16001_/X sky130_fd_sc_hd__a221o_1
X_13213_ _13683_/A vssd1 vssd1 vccd1 vccd1 _13214_/A sky130_fd_sc_hd__buf_4
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14193_ _14694_/A _14193_/B vssd1 vssd1 vccd1 vccd1 _14193_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26179_ _26319_/CLK _26179_/D vssd1 vssd1 vccd1 vccd1 _26179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13144_ _13144_/A vssd1 vssd1 vccd1 vccd1 _14659_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_125_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _14109_/B vssd1 vssd1 vccd1 vccd1 _15972_/B sky130_fd_sc_hd__clkbuf_4
X_17952_ _17948_/X _17951_/X _18071_/S vssd1 vssd1 vccd1 vccd1 _17952_/X sky130_fd_sc_hd__mux2_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16903_ _16812_/A _16957_/B _16902_/X vssd1 vssd1 vccd1 vccd1 _16904_/B sky130_fd_sc_hd__a21boi_4
XFILLER_239_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17883_ _17995_/A _17971_/D vssd1 vssd1 vccd1 vccd1 _17947_/S sky130_fd_sc_hd__nor2_4
XFILLER_266_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19622_ _27055_/Q _21264_/A input179/X _19621_/X vssd1 vssd1 vccd1 vccd1 _19622_/X
+ sky130_fd_sc_hd__a31o_1
X_16834_ _16834_/A _16895_/A _16883_/B vssd1 vssd1 vccd1 vccd1 _16835_/A sky130_fd_sc_hd__and3_2
XFILLER_93_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19553_ _25655_/Q _19563_/B vssd1 vssd1 vccd1 vccd1 _19553_/X sky130_fd_sc_hd__or2_1
XFILLER_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16765_ _22516_/A _16756_/X _16757_/X _16638_/B vssd1 vssd1 vccd1 vccd1 _16765_/X
+ sky130_fd_sc_hd__a22o_2
X_13977_ _13965_/X _13975_/X _13976_/X vssd1 vssd1 vccd1 vccd1 _13977_/X sky130_fd_sc_hd__o21a_1
XFILLER_207_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18504_ _18504_/A vssd1 vssd1 vccd1 vccd1 _18504_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15716_ _15713_/X _15715_/X _15716_/S vssd1 vssd1 vccd1 vccd1 _15716_/X sky130_fd_sc_hd__mux2_1
X_19484_ _19512_/A vssd1 vssd1 vccd1 vccd1 _19484_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_206_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12928_ _14237_/A _14131_/A vssd1 vssd1 vccd1 vccd1 _12929_/A sky130_fd_sc_hd__nand2_1
XFILLER_280_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16696_ _16696_/A _18184_/A vssd1 vssd1 vccd1 vccd1 _18151_/B sky130_fd_sc_hd__xor2_4
XFILLER_262_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18435_ _18435_/A vssd1 vssd1 vccd1 vccd1 _18435_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15647_ _15642_/X _15645_/X _15647_/S vssd1 vssd1 vccd1 vccd1 _15647_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12859_ _25500_/Q _25481_/Q vssd1 vssd1 vccd1 vccd1 _12860_/B sky130_fd_sc_hd__and2b_2
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18366_ _18366_/A vssd1 vssd1 vccd1 vccd1 _18366_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_15_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15578_ _15331_/A _26701_/Q _26829_/Q _15322_/A _16111_/A vssd1 vssd1 vccd1 vccd1
+ _15578_/X sky130_fd_sc_hd__a221o_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17317_ _25526_/Q vssd1 vssd1 vccd1 vccd1 _17317_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14529_ _26780_/Q _26424_/Q _14536_/S vssd1 vssd1 vccd1 vccd1 _14529_/X sky130_fd_sc_hd__mux2_1
X_18297_ _27009_/Q _18756_/A _18296_/X _18821_/A vssd1 vssd1 vccd1 vccd1 _18297_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_159_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17248_ _25504_/Q _17243_/C _17247_/Y vssd1 vssd1 vccd1 vccd1 _25504_/D sky130_fd_sc_hd__o21a_1
XFILLER_190_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17179_ _17179_/A _17195_/B vssd1 vssd1 vccd1 vccd1 _17179_/Y sky130_fd_sc_hd__nand2_1
X_20190_ _20190_/A vssd1 vssd1 vccd1 vccd1 _20299_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22900_ _22900_/A vssd1 vssd1 vccd1 vccd1 _26427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_285_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23880_ _23712_/X _26820_/Q _23882_/S vssd1 vssd1 vccd1 vccd1 _23881_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22831_ _22888_/S vssd1 vssd1 vccd1 vccd1 _22840_/S sky130_fd_sc_hd__buf_2
XFILLER_272_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22762_ _22762_/A vssd1 vssd1 vccd1 vccd1 _26366_/D sky130_fd_sc_hd__clkbuf_1
X_25550_ _27000_/CLK _25550_/D vssd1 vssd1 vccd1 vccd1 _25550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24501_ _24501_/A vssd1 vssd1 vccd1 vccd1 _24501_/X sky130_fd_sc_hd__clkbuf_2
X_21713_ _21718_/A _21713_/B _21713_/C vssd1 vssd1 vccd1 vccd1 _21714_/A sky130_fd_sc_hd__and3_1
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25481_ _26881_/CLK _25481_/D vssd1 vssd1 vccd1 vccd1 _25481_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22693_ _26343_/Q _22691_/X _22705_/S vssd1 vssd1 vccd1 vccd1 _22694_/A sky130_fd_sc_hd__mux2_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27220_ _27221_/CLK _27220_/D vssd1 vssd1 vccd1 vccd1 _27220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24432_ _24381_/X _25610_/Q _24431_/X vssd1 vssd1 vccd1 vccd1 _24693_/B sky130_fd_sc_hd__o21a_4
X_21644_ _25755_/Q _21278_/A _21563_/A _21643_/X vssd1 vssd1 vccd1 vccd1 _21644_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_24_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24363_ _24372_/A _24548_/A vssd1 vssd1 vccd1 vccd1 _24363_/Y sky130_fd_sc_hd__nand2_1
X_27151_ _27227_/CLK _27151_/D vssd1 vssd1 vccd1 vccd1 _27151_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_178_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21575_ _21509_/X _19267_/X _21510_/X _25822_/Q _21547_/X vssd1 vssd1 vccd1 vccd1
+ _21575_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26102_ _26462_/CLK _26102_/D vssd1 vssd1 vccd1 vccd1 _26102_/Q sky130_fd_sc_hd__dfxtp_1
X_23314_ _23314_/A vssd1 vssd1 vccd1 vccd1 _26597_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20526_ _20525_/X _25700_/Q _20530_/S vssd1 vssd1 vccd1 vccd1 _20527_/A sky130_fd_sc_hd__mux2_1
X_27082_ _27196_/CLK _27082_/D vssd1 vssd1 vccd1 vccd1 _27082_/Q sky130_fd_sc_hd__dfxtp_1
X_24294_ _24327_/A _24294_/B _24295_/B vssd1 vssd1 vccd1 vccd1 _26988_/D sky130_fd_sc_hd__nor3_1
XFILLER_166_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26033_ _26592_/CLK _26033_/D vssd1 vssd1 vccd1 vccd1 _26033_/Q sky130_fd_sc_hd__dfxtp_2
X_23245_ _23245_/A vssd1 vssd1 vccd1 vccd1 _26566_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_1_0_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_20457_ _20457_/A _20457_/B vssd1 vssd1 vccd1 vccd1 _20460_/A sky130_fd_sc_hd__nand2_1
XFILLER_107_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23176_ _23176_/A vssd1 vssd1 vccd1 vccd1 _26535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_284_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20388_ _27160_/Q _27094_/Q vssd1 vssd1 vccd1 vccd1 _20389_/B sky130_fd_sc_hd__nand2_1
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22127_ _26161_/Q _22122_/X _22124_/X input255/X _22118_/X vssd1 vssd1 vccd1 vccd1
+ _22127_/X sky130_fd_sc_hd__a221o_1
XFILLER_161_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22058_ _26138_/Q _20903_/X _22066_/S vssd1 vssd1 vccd1 vccd1 _22059_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26935_ _27319_/CLK _26935_/D vssd1 vssd1 vccd1 vccd1 _26935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21009_ _25875_/Q _20891_/X _21015_/S vssd1 vssd1 vccd1 vccd1 _21010_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13900_ _13608_/X _13885_/X _13899_/X _13107_/A vssd1 vssd1 vccd1 vccd1 _13900_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_75_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26866_ _27285_/CLK _26866_/D vssd1 vssd1 vccd1 vccd1 _26866_/Q sky130_fd_sc_hd__dfxtp_1
X_14880_ _12750_/A _14878_/X _14879_/X vssd1 vssd1 vccd1 vccd1 _14881_/B sky130_fd_sc_hd__o21ai_1
XFILLER_130_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13831_ _15999_/A _13831_/B vssd1 vssd1 vccd1 vccd1 _13831_/X sky130_fd_sc_hd__or2_1
X_25817_ _27288_/CLK _25817_/D vssd1 vssd1 vccd1 vccd1 _25817_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26797_ _26797_/CLK _26797_/D vssd1 vssd1 vccd1 vccd1 _26797_/Q sky130_fd_sc_hd__dfxtp_1
X_16550_ _16550_/A _17927_/A vssd1 vssd1 vccd1 vccd1 _16551_/B sky130_fd_sc_hd__nor2_1
XINSDIODE2_208 _19374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13762_ _13762_/A vssd1 vssd1 vccd1 vccd1 _13762_/X sky130_fd_sc_hd__buf_4
X_25748_ _26292_/CLK _25748_/D vssd1 vssd1 vccd1 vccd1 _25748_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_250_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_219 _23562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15501_ _15501_/A vssd1 vssd1 vccd1 vccd1 _15850_/S sky130_fd_sc_hd__buf_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12713_ _13711_/A vssd1 vssd1 vccd1 vccd1 _16072_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16481_ _16481_/A _16481_/B vssd1 vssd1 vccd1 vccd1 _16481_/X sky130_fd_sc_hd__or2_1
XFILLER_231_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13693_ _26788_/Q _26432_/Q _16060_/S vssd1 vssd1 vccd1 vccd1 _13693_/X sky130_fd_sc_hd__mux2_1
X_25679_ _26278_/CLK _25679_/D vssd1 vssd1 vccd1 vccd1 _25679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_280_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18220_ _18552_/A vssd1 vssd1 vccd1 vccd1 _18220_/X sky130_fd_sc_hd__clkbuf_2
X_15432_ _15399_/Y _15413_/Y _15431_/Y _14818_/A _16281_/S vssd1 vssd1 vccd1 vccd1
+ _15432_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_176_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18151_ _18339_/A _18151_/B vssd1 vssd1 vccd1 vccd1 _18151_/Y sky130_fd_sc_hd__nand2_1
X_15363_ _26508_/Q _26380_/Q _15374_/S vssd1 vssd1 vccd1 vccd1 _15363_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17102_ _20978_/A vssd1 vssd1 vccd1 vccd1 _22515_/A sky130_fd_sc_hd__buf_6
X_14314_ _14306_/X _14313_/X _13976_/X vssd1 vssd1 vccd1 vccd1 _14314_/X sky130_fd_sc_hd__o21a_1
XFILLER_184_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18082_ _18347_/S _18081_/X _17981_/Y vssd1 vssd1 vccd1 vccd1 _18413_/A sky130_fd_sc_hd__o21ai_1
X_15294_ _15834_/S vssd1 vssd1 vccd1 vccd1 _15414_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17033_ _17028_/X _16904_/B _17032_/X input224/X vssd1 vssd1 vccd1 vccd1 _17033_/X
+ sky130_fd_sc_hd__a22o_4
X_14245_ _26847_/Q _25761_/Q _14245_/S vssd1 vssd1 vccd1 vccd1 _14245_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14176_ _26068_/Q _25873_/Q _14176_/S vssd1 vssd1 vccd1 vccd1 _14176_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ _15538_/A vssd1 vssd1 vccd1 vccd1 _14647_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _18792_/X _18979_/X _18980_/X _18983_/X vssd1 vssd1 vccd1 vccd1 _18984_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _14001_/B vssd1 vssd1 vccd1 vccd1 _15797_/B sky130_fd_sc_hd__buf_2
X_17935_ _17933_/X _17934_/X _18044_/S vssd1 vssd1 vccd1 vccd1 _17935_/X sky130_fd_sc_hd__mux2_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17866_ _18076_/A _17971_/D vssd1 vssd1 vccd1 vccd1 _17956_/S sky130_fd_sc_hd__or2_4
XFILLER_254_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19605_ _14559_/X _19604_/X _20092_/A _17444_/C vssd1 vssd1 vccd1 vccd1 _19607_/B
+ sky130_fd_sc_hd__o211a_1
X_16817_ _16855_/B vssd1 vssd1 vccd1 vccd1 _16818_/C sky130_fd_sc_hd__clkinv_2
XFILLER_238_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17797_ _13908_/B _17797_/B vssd1 vssd1 vccd1 vccd1 _18539_/B sky130_fd_sc_hd__and2b_1
XFILLER_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19536_ _25649_/Q _19536_/B vssd1 vssd1 vccd1 vccd1 _19536_/X sky130_fd_sc_hd__or2_1
XFILLER_93_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16748_ _16748_/A vssd1 vssd1 vccd1 vccd1 _18932_/B sky130_fd_sc_hd__buf_4
XFILLER_241_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19467_ _27068_/Q _18747_/X _19464_/X _19466_/X _18761_/X vssd1 vssd1 vccd1 vccd1
+ _19467_/X sky130_fd_sc_hd__o221a_2
X_16679_ _25867_/Q _16679_/B _16674_/A vssd1 vssd1 vccd1 vccd1 _16679_/X sky130_fd_sc_hd__or3b_4
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18418_ _18416_/X _18417_/X _18492_/A vssd1 vssd1 vccd1 vccd1 _18419_/B sky130_fd_sc_hd__mux2_1
XFILLER_210_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19398_ _27228_/Q _19462_/B vssd1 vssd1 vccd1 vccd1 _19398_/X sky130_fd_sc_hd__and2_1
XFILLER_148_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18349_ _18347_/X _18348_/X _18349_/S vssd1 vssd1 vccd1 vccd1 _18350_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21360_ _21352_/Y _21358_/X _21359_/X vssd1 vssd1 vccd1 vccd1 _21360_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20311_ _20352_/A _20351_/A vssd1 vssd1 vccd1 vccd1 _20313_/A sky130_fd_sc_hd__and2b_1
X_21291_ _21282_/X _21288_/X _21290_/X vssd1 vssd1 vccd1 vccd1 _21291_/X sky130_fd_sc_hd__a21o_1
Xinput60 dout0[25] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_2
XFILLER_238_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput71 dout0[35] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_1
Xinput82 dout0[45] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__clkbuf_1
Xinput93 dout0[55] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_1
X_23030_ _26486_/Q _22739_/X _23032_/S vssd1 vssd1 vccd1 vccd1 _23031_/A sky130_fd_sc_hd__mux2_1
X_20242_ _20218_/A _20218_/Y _20240_/Y _20241_/X vssd1 vssd1 vccd1 vccd1 _20242_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_89_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20173_ _20173_/A _20173_/B vssd1 vssd1 vccd1 vccd1 _20200_/B sky130_fd_sc_hd__xnor2_1
XFILLER_103_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24981_ _20434_/A _24957_/X _24980_/Y vssd1 vssd1 vccd1 vccd1 _27162_/D sky130_fd_sc_hd__o21a_1
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26720_ _26880_/CLK _26720_/D vssd1 vssd1 vccd1 vccd1 _26720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23932_ _25249_/A _25249_/B _25321_/A vssd1 vssd1 vccd1 vccd1 _23989_/A sky130_fd_sc_hd__nor3_4
XFILLER_130_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26651_ _26715_/CLK _26651_/D vssd1 vssd1 vccd1 vccd1 _26651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23863_ _23684_/X _26812_/Q _23871_/S vssd1 vssd1 vccd1 vccd1 _23864_/A sky130_fd_sc_hd__mux2_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25602_ _25607_/CLK _25602_/D vssd1 vssd1 vccd1 vccd1 _25602_/Q sky130_fd_sc_hd__dfxtp_4
X_22814_ _22814_/A vssd1 vssd1 vccd1 vccd1 _26390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26582_ _27293_/CLK _26582_/D vssd1 vssd1 vccd1 vccd1 _26582_/Q sky130_fd_sc_hd__dfxtp_1
X_23794_ _23794_/A vssd1 vssd1 vccd1 vccd1 _26781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25533_ _26257_/CLK _25533_/D vssd1 vssd1 vccd1 vccd1 _25533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22745_ _23211_/A _23291_/B vssd1 vssd1 vccd1 vccd1 _22802_/A sky130_fd_sc_hd__nor2_8
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22676_ _22743_/S vssd1 vssd1 vccd1 vccd1 _22689_/S sky130_fd_sc_hd__buf_2
XFILLER_201_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25464_ _25464_/A vssd1 vssd1 vccd1 vccd1 _27326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27203_ _27203_/CLK _27203_/D vssd1 vssd1 vccd1 vccd1 _27203_/Q sky130_fd_sc_hd__dfxtp_1
X_24415_ _24415_/A vssd1 vssd1 vccd1 vccd1 _24415_/X sky130_fd_sc_hd__clkbuf_2
X_21627_ _21354_/A _25865_/Q _21626_/Y _21581_/X vssd1 vssd1 vccd1 vccd1 _21627_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_8_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25395_ _25463_/S vssd1 vssd1 vccd1 vccd1 _25404_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_32_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27134_ _27137_/CLK _27134_/D vssd1 vssd1 vccd1 vccd1 _27134_/Q sky130_fd_sc_hd__dfxtp_2
X_21558_ _25959_/Q _21506_/X _21557_/Y _21531_/X vssd1 vssd1 vccd1 vccd1 _25959_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_166_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24346_ _21203_/A _21641_/A _21630_/A _25497_/Q _17701_/X vssd1 vssd1 vccd1 vccd1
+ _24346_/X sky130_fd_sc_hd__a41o_1
X_20509_ _20508_/X _25696_/Q _20509_/S vssd1 vssd1 vccd1 vccd1 _20510_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24277_ _24277_/A vssd1 vssd1 vccd1 vccd1 _24312_/A sky130_fd_sc_hd__buf_2
X_27065_ _27164_/CLK _27065_/D vssd1 vssd1 vccd1 vccd1 _27065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21489_ input52/X input88/X _21489_/S vssd1 vssd1 vccd1 vccd1 _21490_/A sky130_fd_sc_hd__mux2_8
X_14030_ input111/X input146/X _14402_/S vssd1 vssd1 vccd1 vccd1 _14031_/B sky130_fd_sc_hd__mux2_8
XFILLER_180_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23228_ _23228_/A vssd1 vssd1 vccd1 vccd1 _26558_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26016_ _26796_/CLK _26016_/D vssd1 vssd1 vccd1 vccd1 _26016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23159_ _26528_/Q _23063_/X _23161_/S vssd1 vssd1 vccd1 vccd1 _23160_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15981_ _13585_/A _26696_/Q _26824_/Q _15816_/S vssd1 vssd1 vccd1 vccd1 _15981_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17720_ _17725_/D _18161_/B vssd1 vssd1 vccd1 vccd1 _17728_/B sky130_fd_sc_hd__nand2_1
XTAP_5653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26918_ _27278_/CLK _26918_/D vssd1 vssd1 vccd1 vccd1 _26918_/Q sky130_fd_sc_hd__dfxtp_1
X_14932_ _25753_/Q _14931_/Y _15012_/S vssd1 vssd1 vccd1 vccd1 _16458_/B sky130_fd_sc_hd__mux2_2
XTAP_5664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ _24277_/A vssd1 vssd1 vccd1 vccd1 _24723_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26849_ _26913_/CLK _26849_/D vssd1 vssd1 vccd1 vccd1 _26849_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14863_ _14650_/A _14856_/X _14862_/X _14679_/X vssd1 vssd1 vccd1 vccd1 _14863_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16602_ _25671_/Q _16996_/A _18678_/A _16989_/A vssd1 vssd1 vccd1 vccd1 _16660_/A
+ sky130_fd_sc_hd__a22o_4
X_13814_ _13827_/A vssd1 vssd1 vccd1 vccd1 _13814_/X sky130_fd_sc_hd__buf_2
X_17582_ _17995_/B _17564_/X _17572_/X _17581_/Y vssd1 vssd1 vccd1 vccd1 _17583_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14794_ _14794_/A vssd1 vssd1 vccd1 vccd1 _14794_/X sky130_fd_sc_hd__buf_2
XFILLER_204_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19321_ _19392_/A _19327_/A vssd1 vssd1 vccd1 vccd1 _19321_/Y sky130_fd_sc_hd__nor2_1
XFILLER_244_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16533_ _16533_/A vssd1 vssd1 vccd1 vccd1 _16541_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_232_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13745_ _15245_/A _13744_/X _12929_/X vssd1 vssd1 vccd1 vccd1 _13745_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19252_ _19252_/A _19252_/B vssd1 vssd1 vccd1 vccd1 _19252_/X sky130_fd_sc_hd__or2_1
X_16464_ _12860_/B _12869_/X _12878_/Y _12941_/A _12868_/Y vssd1 vssd1 vccd1 vccd1
+ _16464_/X sky130_fd_sc_hd__a41o_1
XFILLER_92_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13676_ _14459_/S vssd1 vssd1 vccd1 vccd1 _13841_/A sky130_fd_sc_hd__clkbuf_4
X_18203_ _18200_/X _18201_/X _18345_/S vssd1 vssd1 vccd1 vccd1 _18203_/X sky130_fd_sc_hd__mux2_1
X_15415_ _26800_/Q _26444_/Q _16361_/S vssd1 vssd1 vccd1 vccd1 _15415_/X sky130_fd_sc_hd__mux2_1
XPHY_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19183_ _19449_/A _19183_/B vssd1 vssd1 vccd1 vccd1 _19183_/Y sky130_fd_sc_hd__nand2_1
XPHY_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16395_ _26547_/Q _26155_/Q _16395_/S vssd1 vssd1 vccd1 vccd1 _16395_/X sky130_fd_sc_hd__mux2_1
XPHY_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18134_ _18303_/S vssd1 vssd1 vccd1 vccd1 _18577_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_200_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15346_ _15245_/X _15345_/X _14604_/A vssd1 vssd1 vccd1 vccd1 _15346_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18065_ _18061_/Y _18064_/X _18202_/A vssd1 vssd1 vccd1 vccd1 _18065_/X sky130_fd_sc_hd__mux2_2
XFILLER_8_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15277_ _15275_/X _15276_/X _16324_/S vssd1 vssd1 vccd1 vccd1 _15277_/X sky130_fd_sc_hd__mux2_1
XFILLER_208_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17016_ _17016_/A vssd1 vssd1 vccd1 vccd1 _17039_/A sky130_fd_sc_hd__clkbuf_2
X_14228_ _14228_/A vssd1 vssd1 vccd1 vccd1 _14228_/X sky130_fd_sc_hd__buf_2
XFILLER_113_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14159_ _26784_/Q _26428_/Q _15902_/S vssd1 vssd1 vccd1 vccd1 _14159_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18967_ _18967_/A _18967_/B vssd1 vssd1 vccd1 vccd1 _18967_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_47_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26531_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17918_ _17897_/X _17915_/X _18492_/A vssd1 vssd1 vccd1 vccd1 _17918_/X sky130_fd_sc_hd__mux2_1
X_18898_ _18898_/A _18898_/B vssd1 vssd1 vccd1 vccd1 _18936_/C sky130_fd_sc_hd__nor2_1
XFILLER_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17849_ _17852_/A _17852_/B vssd1 vssd1 vccd1 vccd1 _17849_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20860_ _25826_/Q vssd1 vssd1 vccd1 vccd1 _20861_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_54_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19519_ _25642_/Q _19523_/B vssd1 vssd1 vccd1 vccd1 _19519_/X sky130_fd_sc_hd__or2_1
XFILLER_263_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20791_ _20791_/A vssd1 vssd1 vccd1 vccd1 _25790_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_550 _25818_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22530_ _22530_/A _22535_/B vssd1 vssd1 vccd1 vccd1 _26289_/D sky130_fd_sc_hd__nor2_1
XFILLER_167_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22461_ _26256_/Q _22470_/B vssd1 vssd1 vccd1 vccd1 _22461_/X sky130_fd_sc_hd__or2_1
XFILLER_210_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24200_ _26957_/Q _24203_/C _17414_/X vssd1 vssd1 vccd1 vccd1 _24200_/Y sky130_fd_sc_hd__a21oi_1
X_21412_ _21408_/Y _21411_/X _21359_/X vssd1 vssd1 vccd1 vccd1 _21412_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_182_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25180_ _24781_/B _25172_/X _25175_/X _27199_/Q _25179_/X vssd1 vssd1 vccd1 vccd1
+ _27199_/D sky130_fd_sc_hd__o221a_1
X_22392_ _22405_/A _22383_/X _22389_/X _22391_/X vssd1 vssd1 vccd1 vccd1 _22392_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24131_ _26932_/Q _23587_/X _24131_/S vssd1 vssd1 vccd1 vccd1 _24132_/A sky130_fd_sc_hd__mux2_1
X_21343_ _21545_/A vssd1 vssd1 vccd1 vccd1 _21343_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24062_ _26901_/Q _23590_/X _24070_/S vssd1 vssd1 vccd1 vccd1 _24063_/A sky130_fd_sc_hd__mux2_1
X_21274_ _25938_/Q _21202_/X _21273_/Y _21262_/X vssd1 vssd1 vccd1 vccd1 _25938_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_190_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23013_ _26478_/Q _22714_/X _23017_/S vssd1 vssd1 vccd1 vccd1 _23014_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20225_ _20225_/A vssd1 vssd1 vccd1 vccd1 _20225_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_270_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20156_ _20135_/A _20134_/B _20134_/A vssd1 vssd1 vccd1 vccd1 _20160_/A sky130_fd_sc_hd__a21boi_1
XFILLER_281_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24964_ hold1/X _24972_/B vssd1 vssd1 vccd1 vccd1 _24964_/Y sky130_fd_sc_hd__nand2_1
X_20087_ _19982_/A _19982_/B _20081_/B vssd1 vssd1 vccd1 vccd1 _20087_/X sky130_fd_sc_hd__a21o_1
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26703_ _27314_/CLK _26703_/D vssd1 vssd1 vccd1 vccd1 _26703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23915_ _23763_/X _26836_/Q _23915_/S vssd1 vssd1 vccd1 vccd1 _23916_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24895_ _24893_/Y _24894_/X _21242_/X vssd1 vssd1 vccd1 vccd1 _27131_/D sky130_fd_sc_hd__a21oi_1
XFILLER_245_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26634_ _27309_/CLK _26634_/D vssd1 vssd1 vccd1 vccd1 _26634_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23846_ _23766_/X _26805_/Q _23854_/S vssd1 vssd1 vccd1 vccd1 _23847_/A sky130_fd_sc_hd__mux2_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26565_ _27308_/CLK _26565_/D vssd1 vssd1 vccd1 vccd1 _26565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20989_ _20989_/A vssd1 vssd1 vccd1 vccd1 _25866_/D sky130_fd_sc_hd__clkbuf_2
X_23777_ _23776_/X _26776_/Q _23780_/S vssd1 vssd1 vccd1 vccd1 _23778_/A sky130_fd_sc_hd__mux2_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13530_ _14806_/A vssd1 vssd1 vccd1 vccd1 _13530_/X sky130_fd_sc_hd__buf_4
X_25516_ _27062_/CLK _25516_/D vssd1 vssd1 vccd1 vccd1 _25516_/Q sky130_fd_sc_hd__dfxtp_1
X_22728_ _26354_/Q _22727_/X _22737_/S vssd1 vssd1 vccd1 vccd1 _22729_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26496_ _27303_/CLK _26496_/D vssd1 vssd1 vccd1 vccd1 _26496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25447_ _25447_/A vssd1 vssd1 vccd1 vccd1 _27318_/D sky130_fd_sc_hd__clkbuf_1
X_13461_ _16031_/S vssd1 vssd1 vccd1 vccd1 _15868_/B sky130_fd_sc_hd__buf_2
X_22659_ _23702_/A vssd1 vssd1 vccd1 vccd1 _22659_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_201_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ _14743_/A _26900_/Q _26772_/Q _15228_/S _14771_/A vssd1 vssd1 vccd1 vccd1
+ _15200_/X sky130_fd_sc_hd__a221o_1
XFILLER_173_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16180_ _16336_/A _16178_/X _16179_/X vssd1 vssd1 vccd1 vccd1 _16180_/X sky130_fd_sc_hd__o21a_1
X_13392_ _12913_/A _13391_/X _12929_/X vssd1 vssd1 vccd1 vccd1 _13392_/X sky130_fd_sc_hd__a21o_1
X_25378_ _25378_/A vssd1 vssd1 vccd1 vccd1 _25387_/S sky130_fd_sc_hd__buf_4
XFILLER_127_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15131_ _17787_/A _17786_/A vssd1 vssd1 vccd1 vccd1 _15132_/B sky130_fd_sc_hd__and2_1
X_27117_ _27117_/CLK _27117_/D vssd1 vssd1 vccd1 vccd1 _27117_/Q sky130_fd_sc_hd__dfxtp_4
X_24329_ _24335_/A _24329_/B vssd1 vssd1 vccd1 vccd1 _24329_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27048_ _27049_/CLK _27048_/D vssd1 vssd1 vccd1 vccd1 _27048_/Q sky130_fd_sc_hd__dfxtp_1
X_15062_ _26646_/Q _26742_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _15062_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14013_ _26070_/Q _14001_/B _14495_/A _14012_/X vssd1 vssd1 vccd1 vccd1 _14013_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19870_ _19870_/A _19870_/B vssd1 vssd1 vccd1 vccd1 _19870_/X sky130_fd_sc_hd__or2_1
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18821_ _18821_/A vssd1 vssd1 vccd1 vccd1 _18821_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_191_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18752_ _18816_/A vssd1 vssd1 vccd1 vccd1 _18752_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15964_ _26856_/Q _25770_/Q _15964_/S vssd1 vssd1 vccd1 vccd1 _15964_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput250 localMemory_wb_sel_i[3] vssd1 vssd1 vccd1 vccd1 input250/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput261 manufacturerID[7] vssd1 vssd1 vccd1 vccd1 _22146_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17703_ _24350_/S _21219_/A vssd1 vssd1 vccd1 vccd1 _17703_/X sky130_fd_sc_hd__and2_1
XFILLER_76_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput272 partID[2] vssd1 vssd1 vccd1 vccd1 _22166_/A sky130_fd_sc_hd__clkbuf_1
XTAP_5483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14915_ _14913_/X _14914_/X _15004_/S vssd1 vssd1 vccd1 vccd1 _14915_/X sky130_fd_sc_hd__mux2_1
Xinput283 versionID[3] vssd1 vssd1 vccd1 vccd1 input283/X sky130_fd_sc_hd__buf_2
XTAP_5494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18683_ _18683_/A _18683_/B vssd1 vssd1 vccd1 vccd1 _18683_/X sky130_fd_sc_hd__or2_1
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15895_ _26921_/Q _26405_/Q _15895_/S vssd1 vssd1 vccd1 vccd1 _15895_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17634_ _17634_/A vssd1 vssd1 vccd1 vccd1 _17650_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_251_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14846_ _26937_/Q _14846_/B vssd1 vssd1 vccd1 vccd1 _14846_/X sky130_fd_sc_hd__or2_1
XFILLER_1_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17565_ _25910_/Q _17517_/X _13748_/B _17525_/X vssd1 vssd1 vccd1 vccd1 _17565_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_14777_ _14777_/A vssd1 vssd1 vccd1 vccd1 _14778_/A sky130_fd_sc_hd__buf_6
XFILLER_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19304_ _27063_/Q _18811_/X _19301_/X _19303_/X _18823_/X vssd1 vssd1 vccd1 vccd1
+ _19304_/X sky130_fd_sc_hd__o221a_2
X_16516_ _16517_/A _16512_/X _16515_/X _12758_/A vssd1 vssd1 vccd1 vccd1 _16521_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_220_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13728_ _26916_/Q _26400_/Q _15464_/B vssd1 vssd1 vccd1 vccd1 _13728_/X sky130_fd_sc_hd__mux2_1
XFILLER_210_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17496_ _17704_/S vssd1 vssd1 vccd1 vccd1 _24350_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_165_wb_clk_i clkbuf_opt_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26282_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_231_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19235_ _19252_/B _19235_/B vssd1 vssd1 vccd1 vccd1 _19235_/Y sky130_fd_sc_hd__nand2_1
X_16447_ _16280_/S _16439_/X _16446_/X _14723_/A vssd1 vssd1 vccd1 vccd1 _16447_/X
+ sky130_fd_sc_hd__a31o_1
X_13659_ _13252_/A _25767_/Q _16020_/S _26853_/Q _13344_/A vssd1 vssd1 vccd1 vccd1
+ _13659_/X sky130_fd_sc_hd__o221a_1
XFILLER_177_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19166_ _27155_/Q _19302_/B vssd1 vssd1 vccd1 vccd1 _19166_/X sky130_fd_sc_hd__or2_1
X_16378_ _16376_/X _16377_/X _16378_/S vssd1 vssd1 vccd1 vccd1 _16378_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18117_ _18119_/A _18119_/B vssd1 vssd1 vccd1 vccd1 _18121_/A sky130_fd_sc_hd__or2_1
X_15329_ _15327_/X _15328_/X _16278_/S vssd1 vssd1 vccd1 vccd1 _15329_/X sky130_fd_sc_hd__mux2_1
X_19097_ _25553_/Q _18459_/A _19096_/X _17688_/A _18466_/A vssd1 vssd1 vccd1 vccd1
+ _19097_/X sky130_fd_sc_hd__a221o_1
XFILLER_172_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18048_ _17899_/X _17909_/X _18062_/S vssd1 vssd1 vccd1 vccd1 _18048_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20010_ _25737_/Q vssd1 vssd1 vccd1 vccd1 _20656_/A sky130_fd_sc_hd__buf_8
XFILLER_235_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19999_ _19999_/A _19999_/B _19999_/C vssd1 vssd1 vccd1 vccd1 _19999_/Y sky130_fd_sc_hd__nor3_1
XFILLER_274_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21961_ _24004_/B _23139_/A vssd1 vssd1 vccd1 vccd1 _22018_/A sky130_fd_sc_hd__nor2_4
XFILLER_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23700_ _23699_/X _26752_/Q _23700_/S vssd1 vssd1 vccd1 vccd1 _23701_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20912_ _20912_/A vssd1 vssd1 vccd1 vccd1 _25841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_255_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21892_ _20484_/X _26064_/Q _21900_/S vssd1 vssd1 vccd1 vccd1 _21893_/A sky130_fd_sc_hd__mux2_1
X_24680_ _24701_/A vssd1 vssd1 vccd1 vccd1 _24680_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_270_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23631_ _23631_/A vssd1 vssd1 vccd1 vccd1 _26723_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20843_ _20843_/A vssd1 vssd1 vccd1 vccd1 _25817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26350_ _26610_/CLK _26350_/D vssd1 vssd1 vccd1 vccd1 _26350_/Q sky130_fd_sc_hd__dfxtp_1
X_20774_ _20774_/A vssd1 vssd1 vccd1 vccd1 _20783_/S sky130_fd_sc_hd__clkbuf_4
X_23562_ _23562_/A vssd1 vssd1 vccd1 vccd1 _23562_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_223_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_380 _17000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25301_ _25301_/A vssd1 vssd1 vccd1 vccd1 _27253_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_391 _17031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22513_ _22513_/A _22513_/B vssd1 vssd1 vccd1 vccd1 _22514_/A sky130_fd_sc_hd__and2_1
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26281_ _26286_/CLK _26281_/D vssd1 vssd1 vccd1 vccd1 _26281_/Q sky130_fd_sc_hd__dfxtp_1
X_23493_ _23493_/A vssd1 vssd1 vccd1 vccd1 _23502_/S sky130_fd_sc_hd__buf_6
XFILLER_195_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22444_ _26250_/Q _22444_/B vssd1 vssd1 vccd1 vccd1 _22444_/X sky130_fd_sc_hd__or2_1
XFILLER_210_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25232_ _27222_/Q _25217_/X _25231_/X _25221_/X vssd1 vssd1 vccd1 vccd1 _27222_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22375_ _22375_/A vssd1 vssd1 vccd1 vccd1 _26235_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25163_ _25754_/Q _25138_/A _25162_/X vssd1 vssd1 vccd1 vccd1 _25163_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21326_ _21276_/X _21325_/X _21227_/X vssd1 vssd1 vccd1 vccd1 _21326_/Y sky130_fd_sc_hd__o21ai_1
X_24114_ _26924_/Q _23562_/X _24120_/S vssd1 vssd1 vccd1 vccd1 _24115_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25094_ _20666_/A _25086_/X _25093_/X vssd1 vssd1 vccd1 vccd1 _25094_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_124_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24045_ _24045_/A vssd1 vssd1 vccd1 vccd1 _26893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21257_ input54/X input69/X _21356_/S vssd1 vssd1 vccd1 vccd1 _21258_/B sky130_fd_sc_hd__mux2_8
XFILLER_278_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20208_ _20208_/A _20260_/B vssd1 vssd1 vccd1 vccd1 _20208_/Y sky130_fd_sc_hd__nor2_1
XFILLER_277_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21188_ _21188_/A _21188_/B vssd1 vssd1 vccd1 vccd1 _21189_/A sky130_fd_sc_hd__or2_1
X_20139_ _22507_/A _20078_/X _20130_/X _20138_/X _20076_/X vssd1 vssd1 vccd1 vccd1
+ _25677_/D sky130_fd_sc_hd__o221a_1
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25996_ _27227_/CLK _25996_/D vssd1 vssd1 vccd1 vccd1 _25996_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24947_ _27148_/Q _24927_/X _24946_/Y vssd1 vssd1 vccd1 vccd1 _27148_/D sky130_fd_sc_hd__o21a_1
X_12961_ _12961_/A _20485_/A _21887_/B _21888_/B vssd1 vssd1 vccd1 vccd1 _12963_/C
+ sky130_fd_sc_hd__or4_1
XINSDIODE2_40 _19441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_51 _20637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_62 _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14700_ _14698_/X _14699_/X _14700_/S vssd1 vssd1 vccd1 vccd1 _14700_/X sky130_fd_sc_hd__mux2_1
XFILLER_234_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_73 _20681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_84 _23712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _26796_/Q _26440_/Q _16271_/S vssd1 vssd1 vccd1 vccd1 _15680_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_95 _21305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12892_ _12892_/A vssd1 vssd1 vccd1 vccd1 _13911_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_24878_ _27126_/Q _24890_/B vssd1 vssd1 vccd1 vccd1 _24878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _15548_/S vssd1 vssd1 vccd1 vccd1 _16305_/A sky130_fd_sc_hd__buf_4
X_26617_ _27321_/CLK _26617_/D vssd1 vssd1 vccd1 vccd1 _26617_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23829_ _23829_/A vssd1 vssd1 vccd1 vccd1 _26797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17350_ _17347_/X _17351_/C _25536_/Q vssd1 vssd1 vccd1 vccd1 _17352_/B sky130_fd_sc_hd__a21oi_1
XFILLER_14_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14562_ _14562_/A _14562_/B vssd1 vssd1 vccd1 vccd1 _14562_/X sky130_fd_sc_hd__and2_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26548_ _26744_/CLK _26548_/D vssd1 vssd1 vccd1 vccd1 _26548_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _26869_/Q _25783_/Q _16301_/S vssd1 vssd1 vccd1 vccd1 _16301_/X sky130_fd_sc_hd__mux2_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13513_ _13510_/X _13511_/X _15606_/A vssd1 vssd1 vccd1 vccd1 _13513_/X sky130_fd_sc_hd__mux2_1
X_17281_ _17278_/X _17282_/C _25515_/Q vssd1 vssd1 vccd1 vccd1 _17283_/B sky130_fd_sc_hd__a21oi_1
XFILLER_201_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _13578_/A _14492_/X _14486_/A vssd1 vssd1 vccd1 vccd1 _14528_/B sky130_fd_sc_hd__o21ai_1
X_26479_ _27287_/CLK _26479_/D vssd1 vssd1 vccd1 vccd1 _26479_/Q sky130_fd_sc_hd__dfxtp_1
X_19020_ _25519_/Q _18807_/X _18808_/X _25551_/Q vssd1 vssd1 vccd1 vccd1 _19020_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16232_ _26931_/Q _16301_/S vssd1 vssd1 vccd1 vccd1 _16232_/X sky130_fd_sc_hd__or2_1
X_13444_ _13439_/X _13443_/X _13711_/A vssd1 vssd1 vccd1 vccd1 _13444_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16163_ _26673_/Q _25713_/Q _16163_/S vssd1 vssd1 vccd1 vccd1 _16163_/X sky130_fd_sc_hd__mux2_1
X_13375_ _14317_/B vssd1 vssd1 vccd1 vccd1 _16581_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15114_ _26806_/Q _26450_/Q _15119_/S vssd1 vssd1 vccd1 vccd1 _15114_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16094_ _26083_/Q _25888_/Q _16271_/S vssd1 vssd1 vccd1 vccd1 _16094_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15045_ _26678_/Q _25718_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _15045_/X sky130_fd_sc_hd__mux2_1
X_19922_ _19980_/C _19923_/A _19976_/C vssd1 vssd1 vccd1 vccd1 _19951_/B sky130_fd_sc_hd__or3b_1
XFILLER_107_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19853_ _19853_/A _19853_/B _19808_/A _19830_/C vssd1 vssd1 vccd1 vccd1 _19853_/X
+ sky130_fd_sc_hd__or4bb_1
XFILLER_269_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18804_ _18792_/X _18796_/X _18803_/X vssd1 vssd1 vccd1 vccd1 _18804_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16996_ _16996_/A vssd1 vssd1 vccd1 vccd1 _16996_/X sky130_fd_sc_hd__clkbuf_2
X_19784_ _19790_/A _27072_/Q vssd1 vssd1 vccd1 vccd1 _19784_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_95_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15947_ _13638_/X _23552_/A _15946_/Y _13214_/A vssd1 vssd1 vccd1 vccd1 _20008_/A
+ sky130_fd_sc_hd__o211ai_4
X_18735_ _18734_/X _18643_/A _18735_/S vssd1 vssd1 vccd1 vccd1 _18735_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18666_ _18666_/A _18666_/B vssd1 vssd1 vccd1 vccd1 _18666_/Y sky130_fd_sc_hd__nor2_1
XFILLER_252_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ _25611_/Q _14594_/A _15877_/X _12977_/A vssd1 vssd1 vccd1 vccd1 _15913_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_236_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17617_ _17560_/X _17623_/B _14026_/X _17554_/X _25923_/Q vssd1 vssd1 vccd1 vccd1
+ _17617_/Y sky130_fd_sc_hd__o32ai_1
XFILLER_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14829_ _20701_/A _19442_/A _15012_/S vssd1 vssd1 vccd1 vccd1 _17779_/A sky130_fd_sc_hd__mux2_2
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18597_ _18597_/A vssd1 vssd1 vccd1 vccd1 _18597_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_240_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17548_ _17548_/A _17548_/B vssd1 vssd1 vccd1 vccd1 _25570_/D sky130_fd_sc_hd__nor2_1
XFILLER_177_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17479_ _16673_/C _17459_/A _17478_/X _17458_/B vssd1 vssd1 vccd1 vccd1 _21209_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_177_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19218_ _19218_/A vssd1 vssd1 vccd1 vccd1 _19218_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20490_ _24004_/A _25249_/C vssd1 vssd1 vccd1 vccd1 _20597_/A sky130_fd_sc_hd__or2_4
XFILLER_192_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19149_ _18976_/X _19145_/X _19148_/X _19003_/X vssd1 vssd1 vccd1 vccd1 _19149_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22160_ _22179_/A vssd1 vssd1 vccd1 vccd1 _22160_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21111_ _21111_/A vssd1 vssd1 vccd1 vccd1 _25911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_62_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27307_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_172_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22091_ _26153_/Q _20951_/X _22099_/S vssd1 vssd1 vccd1 vccd1 _22092_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21042_ _25890_/Q _20939_/X _21048_/S vssd1 vssd1 vccd1 vccd1 _21043_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25850_ _27284_/CLK _25850_/D vssd1 vssd1 vccd1 vccd1 _25850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24801_ _24801_/A vssd1 vssd1 vccd1 vccd1 _24877_/A sky130_fd_sc_hd__buf_2
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25781_ _26611_/CLK _25781_/D vssd1 vssd1 vccd1 vccd1 _25781_/Q sky130_fd_sc_hd__dfxtp_1
X_22993_ _26469_/Q _22685_/X _22995_/S vssd1 vssd1 vccd1 vccd1 _22994_/A sky130_fd_sc_hd__mux2_1
XFILLER_274_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24732_ _24739_/A _24732_/B vssd1 vssd1 vccd1 vccd1 _24732_/Y sky130_fd_sc_hd__nand2_4
XFILLER_215_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21944_ _20592_/X _26088_/Q _21944_/S vssd1 vssd1 vccd1 vccd1 _21945_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24663_ _24920_/A vssd1 vssd1 vccd1 vccd1 _24664_/B sky130_fd_sc_hd__inv_2
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21875_ _21867_/Y _21872_/X _21874_/X _20697_/X vssd1 vssd1 vccd1 vccd1 _26061_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_257_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26402_ _27277_/CLK _26402_/D vssd1 vssd1 vccd1 vccd1 _26402_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_199_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23614_ _23682_/S vssd1 vssd1 vccd1 vccd1 _23623_/S sky130_fd_sc_hd__clkbuf_4
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20826_ _25809_/Q vssd1 vssd1 vccd1 vccd1 _20827_/A sky130_fd_sc_hd__clkbuf_1
X_24594_ _27053_/Q _24589_/X _24592_/Y _24593_/X vssd1 vssd1 vccd1 vccd1 _27053_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_70_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26333_ _26462_/CLK _26333_/D vssd1 vssd1 vccd1 vccd1 _26333_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_24_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23545_ _23545_/A vssd1 vssd1 vccd1 vccd1 _26694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20757_ _20563_/X _25775_/Q _20761_/S vssd1 vssd1 vccd1 vccd1 _20758_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26264_ _26264_/CLK _26264_/D vssd1 vssd1 vccd1 vccd1 _26264_/Q sky130_fd_sc_hd__dfxtp_1
X_23476_ _26669_/Q _23092_/X _23480_/S vssd1 vssd1 vccd1 vccd1 _23477_/A sky130_fd_sc_hd__mux2_1
X_20688_ _26285_/Q _20686_/X _20687_/Y _20684_/X vssd1 vssd1 vccd1 vccd1 _25748_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25215_ _27055_/Q _21874_/A input179/X _25214_/X _25199_/A vssd1 vssd1 vccd1 vccd1
+ _25215_/X sky130_fd_sc_hd__a41o_1
X_22427_ _26244_/Q _22430_/B vssd1 vssd1 vccd1 vccd1 _22427_/X sky130_fd_sc_hd__or2_1
XFILLER_40_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26195_ _26250_/CLK _26195_/D vssd1 vssd1 vccd1 vccd1 _26195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13160_ _15174_/A _13154_/X _13158_/X _15039_/A vssd1 vssd1 vccd1 vccd1 _13160_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_152_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25146_ _19315_/A _25138_/X _25145_/X vssd1 vssd1 vccd1 vccd1 _25146_/X sky130_fd_sc_hd__o21a_1
X_22358_ _22361_/A _22361_/B vssd1 vssd1 vccd1 vccd1 _22381_/A sky130_fd_sc_hd__nand2_1
XFILLER_151_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21309_ _21309_/A vssd1 vssd1 vccd1 vccd1 _21573_/A sky130_fd_sc_hd__clkbuf_4
X_13091_ _15630_/A vssd1 vssd1 vccd1 vccd1 _15653_/S sky130_fd_sc_hd__clkbuf_4
X_22289_ _26208_/Q _22284_/X _22287_/X _22288_/X vssd1 vssd1 vccd1 vccd1 _26208_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25077_ _24696_/Y _25070_/X _25076_/Y _25055_/X vssd1 vssd1 vccd1 vccd1 _25077_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24028_ _24074_/S vssd1 vssd1 vccd1 vccd1 _24037_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16850_ _16864_/A _16850_/B vssd1 vssd1 vccd1 vccd1 _16851_/A sky130_fd_sc_hd__and2_1
XFILLER_278_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15801_ _27245_/Q _15820_/B vssd1 vssd1 vccd1 vccd1 _15801_/X sky130_fd_sc_hd__or2_1
XFILLER_266_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16781_ _22528_/A _16769_/X _16770_/X _16575_/B vssd1 vssd1 vccd1 vccd1 _16781_/X
+ sky130_fd_sc_hd__a22o_4
X_25979_ _27022_/CLK _25979_/D vssd1 vssd1 vccd1 vccd1 _25979_/Q sky130_fd_sc_hd__dfxtp_4
X_13993_ _13993_/A vssd1 vssd1 vccd1 vccd1 _14520_/S sky130_fd_sc_hd__buf_2
XFILLER_59_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18520_ _27044_/Q _18503_/X _18512_/X _18518_/X _18519_/X vssd1 vssd1 vccd1 vccd1
+ _18520_/X sky130_fd_sc_hd__o221a_1
XFILLER_281_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15732_ _13585_/X _26407_/Q _15727_/S _15731_/X vssd1 vssd1 vccd1 vccd1 _15732_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12944_ _12860_/B _12878_/Y _12941_/A _12872_/A vssd1 vssd1 vccd1 vccd1 _12944_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18451_ _27011_/Q _18116_/B _18161_/C _17742_/Y vssd1 vssd1 vccd1 vccd1 _18451_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ _16088_/A _15663_/B vssd1 vssd1 vccd1 vccd1 _15663_/X sky130_fd_sc_hd__or2_1
XFILLER_283_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12875_ _14411_/A vssd1 vssd1 vccd1 vccd1 _15954_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _17430_/A _17408_/C vssd1 vssd1 vccd1 vccd1 _17402_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _25660_/Q _24351_/B _14613_/X vssd1 vssd1 vccd1 vccd1 _14614_/X sky130_fd_sc_hd__a21o_1
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _18382_/A vssd1 vssd1 vccd1 vccd1 _18382_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _15587_/X _15593_/X _13314_/A vssd1 vssd1 vccd1 vccd1 _15594_/Y sky130_fd_sc_hd__o21ai_2
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _25531_/Q _17333_/B vssd1 vssd1 vccd1 vccd1 _17341_/C sky130_fd_sc_hd__and2_2
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14543_/X _14544_/X _14552_/S vssd1 vssd1 vccd1 vccd1 _14545_/X sky130_fd_sc_hd__mux2_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17264_ _17283_/A _17264_/B _17265_/B vssd1 vssd1 vccd1 vccd1 _25509_/D sky130_fd_sc_hd__nor3_1
X_14476_ _14468_/A _14474_/X _14475_/X _14067_/X vssd1 vssd1 vccd1 vccd1 _14476_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_197_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19003_ _19003_/A vssd1 vssd1 vccd1 vccd1 _19003_/X sky130_fd_sc_hd__clkbuf_2
X_16215_ _26675_/Q _25715_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _16215_/X sky130_fd_sc_hd__mux2_1
X_13427_ _15806_/S vssd1 vssd1 vccd1 vccd1 _15473_/S sky130_fd_sc_hd__buf_2
XFILLER_220_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17195_ _17195_/A _17195_/B vssd1 vssd1 vccd1 vccd1 _17195_/Y sky130_fd_sc_hd__nand2_1
X_16146_ _25890_/Q _16310_/B vssd1 vssd1 vccd1 vccd1 _16146_/X sky130_fd_sc_hd__or2_1
X_13358_ _13358_/A vssd1 vssd1 vccd1 vccd1 _13359_/A sky130_fd_sc_hd__buf_2
XFILLER_143_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16077_ _26539_/Q _26147_/Q _16078_/S vssd1 vssd1 vccd1 vccd1 _16077_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13289_ _26499_/Q _26371_/Q _16087_/S vssd1 vssd1 vccd1 vccd1 _13290_/B sky130_fd_sc_hd__mux2_1
XFILLER_142_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15028_ _14877_/S _15025_/X _15027_/X _14661_/A vssd1 vssd1 vccd1 vccd1 _15028_/X
+ sky130_fd_sc_hd__a211o_1
X_19905_ _19905_/A vssd1 vssd1 vccd1 vccd1 _19905_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19836_ _19833_/X _19845_/B _19835_/Y _20248_/A vssd1 vssd1 vccd1 vccd1 _19837_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_110_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19767_ _20034_/B vssd1 vssd1 vccd1 vccd1 _19824_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_110_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput3 coreIndex[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_84_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16979_ _16878_/X _16954_/X _16956_/X _16877_/X _16978_/X vssd1 vssd1 vccd1 vccd1
+ _16980_/C sky130_fd_sc_hd__a221o_1
XFILLER_284_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18718_ _19287_/B vssd1 vssd1 vccd1 vccd1 _18719_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19698_ _19771_/A vssd1 vssd1 vccd1 vccd1 _19698_/X sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_180_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26744_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_149_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18649_ _25734_/Q _18650_/B vssd1 vssd1 vccd1 vccd1 _18843_/D sky130_fd_sc_hd__and2_2
XFILLER_37_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21660_ _25971_/Q input206/X _21662_/S vssd1 vssd1 vccd1 vccd1 _21661_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20611_ _20611_/A vssd1 vssd1 vccd1 vccd1 _25720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21591_ _19315_/A _21545_/X _21563_/X _21590_/X vssd1 vssd1 vccd1 vccd1 _21591_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_177_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20542_ _23725_/A vssd1 vssd1 vccd1 vccd1 _20542_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23330_ _23330_/A vssd1 vssd1 vccd1 vccd1 _26604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_257_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20473_ _19766_/A _20471_/Y _20472_/X _20015_/A vssd1 vssd1 vccd1 vccd1 _20473_/X
+ sky130_fd_sc_hd__a31o_1
X_23261_ _23261_/A vssd1 vssd1 vccd1 vccd1 _26573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25000_ _25159_/B vssd1 vssd1 vccd1 vccd1 _25000_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22212_ _26186_/Q _22201_/X _22206_/X _22211_/X _22203_/X vssd1 vssd1 vccd1 vccd1
+ _22212_/X sky130_fd_sc_hd__a221o_1
X_23192_ _26543_/Q _23111_/X _23194_/S vssd1 vssd1 vccd1 vccd1 _23193_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22143_ _26166_/Q _22122_/A _22140_/X input260/X _22137_/X vssd1 vssd1 vccd1 vccd1
+ _22143_/X sky130_fd_sc_hd__a221o_1
XFILLER_279_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput340 _16886_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[15] sky130_fd_sc_hd__buf_2
Xoutput351 _16950_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[25] sky130_fd_sc_hd__buf_2
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput362 _16832_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[6] sky130_fd_sc_hd__buf_2
X_26951_ _26987_/CLK _26951_/D vssd1 vssd1 vccd1 vccd1 _26951_/Q sky130_fd_sc_hd__dfxtp_1
X_22074_ _22074_/A vssd1 vssd1 vccd1 vccd1 _26145_/D sky130_fd_sc_hd__clkbuf_1
Xoutput373 _16682_/X vssd1 vssd1 vccd1 vccd1 csb0[1] sky130_fd_sc_hd__buf_2
XFILLER_121_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput384 _17031_/X vssd1 vssd1 vccd1 vccd1 din0[17] sky130_fd_sc_hd__buf_2
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput395 _17045_/X vssd1 vssd1 vccd1 vccd1 din0[27] sky130_fd_sc_hd__buf_2
X_21025_ _21025_/A vssd1 vssd1 vccd1 vccd1 _25882_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25902_ _26278_/CLK _25902_/D vssd1 vssd1 vccd1 vccd1 _25902_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_86_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26882_ _26917_/CLK _26882_/D vssd1 vssd1 vccd1 vccd1 _26882_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_259_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25833_ _26462_/CLK _25833_/D vssd1 vssd1 vccd1 vccd1 _25833_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25764_ _27269_/CLK _25764_/D vssd1 vssd1 vccd1 vccd1 _25764_/Q sky130_fd_sc_hd__dfxtp_1
X_22976_ _26461_/Q _22659_/X _22984_/S vssd1 vssd1 vccd1 vccd1 _22977_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24715_ _24725_/A _24715_/B vssd1 vssd1 vccd1 vccd1 _24715_/Y sky130_fd_sc_hd__nand2_2
XFILLER_204_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21927_ _20559_/X _26080_/Q _21933_/S vssd1 vssd1 vccd1 vccd1 _21928_/A sky130_fd_sc_hd__mux2_1
X_25695_ _26593_/CLK _25695_/D vssd1 vssd1 vccd1 vccd1 _25695_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24646_ _19640_/A _19634_/B _24636_/A _24645_/Y vssd1 vssd1 vccd1 vccd1 _24646_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_163_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21858_ _26057_/Q _20961_/X _21860_/S vssd1 vssd1 vccd1 vccd1 _21859_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20809_ _20809_/A vssd1 vssd1 vccd1 vccd1 _25800_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24577_ _24577_/A _24582_/B vssd1 vssd1 vccd1 vccd1 _24577_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21789_ _20617_/X _26027_/Q _21791_/S vssd1 vssd1 vccd1 vccd1 _21790_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26316_ _26319_/CLK _26316_/D vssd1 vssd1 vccd1 vccd1 _26316_/Q sky130_fd_sc_hd__dfxtp_2
X_14330_ _14330_/A _14330_/B _14330_/C vssd1 vssd1 vccd1 vccd1 _14330_/X sky130_fd_sc_hd__or3_1
XFILLER_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23528_ _26689_/Q _23526_/X _23540_/S vssd1 vssd1 vccd1 vccd1 _23529_/A sky130_fd_sc_hd__mux2_1
X_27296_ _27297_/CLK _27296_/D vssd1 vssd1 vccd1 vccd1 _27296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14261_ _13857_/X _14254_/X _14260_/X _13163_/A vssd1 vssd1 vccd1 vccd1 _14261_/X
+ sky130_fd_sc_hd__o211a_1
X_26247_ _26248_/CLK _26247_/D vssd1 vssd1 vccd1 vccd1 _26247_/Q sky130_fd_sc_hd__dfxtp_1
X_23459_ _23459_/A vssd1 vssd1 vccd1 vccd1 _26661_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16000_ _15509_/A _15997_/X _15999_/X _15311_/A vssd1 vssd1 vccd1 vccd1 _16000_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13212_ _13212_/A vssd1 vssd1 vccd1 vccd1 _13683_/A sky130_fd_sc_hd__buf_2
X_26178_ _26186_/CLK _26178_/D vssd1 vssd1 vccd1 vccd1 _26178_/Q sky130_fd_sc_hd__dfxtp_1
X_14192_ _25576_/Q _14187_/A _14187_/Y _14193_/B vssd1 vssd1 vccd1 vccd1 _14192_/X
+ sky130_fd_sc_hd__o211a_1
X_13143_ _13159_/A vssd1 vssd1 vccd1 vccd1 _13144_/A sky130_fd_sc_hd__buf_2
X_25129_ _22520_/A _25119_/X _25114_/X _16606_/Y _25106_/X vssd1 vssd1 vccd1 vccd1
+ _25129_/X sky130_fd_sc_hd__a221o_1
XFILLER_125_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13074_ _13590_/A vssd1 vssd1 vccd1 vccd1 _14109_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_152_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17951_ _17949_/X _17950_/X _18067_/S vssd1 vssd1 vccd1 vccd1 _17951_/X sky130_fd_sc_hd__mux2_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16902_ _16955_/B _16818_/C _16852_/X _16868_/A _16939_/B vssd1 vssd1 vccd1 vccd1
+ _16902_/X sky130_fd_sc_hd__o221a_1
XFILLER_239_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17882_ _17957_/S vssd1 vssd1 vccd1 vccd1 _17990_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19621_ _27061_/Q _19617_/B input185/X _19620_/X vssd1 vssd1 vccd1 vccd1 _19621_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_76_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16833_ _16833_/A _16833_/B vssd1 vssd1 vccd1 vccd1 _16883_/B sky130_fd_sc_hd__and2_2
XFILLER_226_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19552_ _19552_/A vssd1 vssd1 vccd1 vccd1 _19563_/B sky130_fd_sc_hd__clkbuf_1
X_16764_ _25681_/Q vssd1 vssd1 vccd1 vccd1 _22516_/A sky130_fd_sc_hd__buf_2
XFILLER_19_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13976_ _13976_/A vssd1 vssd1 vccd1 vccd1 _13976_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_207_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15715_ _26635_/Q _26731_/Q _15988_/S vssd1 vssd1 vccd1 vccd1 _15715_/X sky130_fd_sc_hd__mux2_1
X_18503_ _18503_/A vssd1 vssd1 vccd1 vccd1 _18503_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12927_ _13569_/A vssd1 vssd1 vccd1 vccd1 _14237_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_206_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19483_ _19551_/A vssd1 vssd1 vccd1 vccd1 _19512_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16695_ _14562_/X _16706_/A vssd1 vssd1 vccd1 vccd1 _18184_/A sky130_fd_sc_hd__and2b_2
XFILLER_206_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15646_ _15646_/A vssd1 vssd1 vccd1 vccd1 _15647_/S sky130_fd_sc_hd__clkbuf_4
X_18434_ _18530_/B _18434_/B vssd1 vssd1 vccd1 vccd1 _18434_/Y sky130_fd_sc_hd__nor2_1
XFILLER_221_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12858_ _25500_/Q _25480_/Q vssd1 vssd1 vccd1 vccd1 _12878_/B sky130_fd_sc_hd__and2b_1
XFILLER_22_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18365_ _18362_/X _18363_/X _18364_/X vssd1 vssd1 vccd1 vccd1 _18365_/Y sky130_fd_sc_hd__o21ai_4
X_15577_ _13321_/A _15574_/X _15576_/X _13291_/A vssd1 vssd1 vccd1 vccd1 _15581_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12789_ _13269_/A _25595_/Q vssd1 vssd1 vccd1 vccd1 _17218_/A sky130_fd_sc_hd__nand2_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _25525_/Q _17314_/B _17315_/Y vssd1 vssd1 vccd1 vccd1 _25525_/D sky130_fd_sc_hd__o21a_1
XFILLER_187_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14528_ _14528_/A _14528_/B vssd1 vssd1 vccd1 vccd1 _23508_/A sky130_fd_sc_hd__and2_2
XFILLER_30_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18296_ _27137_/Q _18757_/A vssd1 vssd1 vccd1 vccd1 _18296_/X sky130_fd_sc_hd__or2_1
X_17247_ _17285_/A _17253_/C vssd1 vssd1 vccd1 vccd1 _17247_/Y sky130_fd_sc_hd__nor2_1
X_14459_ _25798_/Q _27232_/Q _14459_/S vssd1 vssd1 vccd1 vccd1 _14459_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17178_ _14804_/X _17170_/X _17177_/X _17175_/X vssd1 vssd1 vccd1 vccd1 _25485_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16129_ _15245_/A _15871_/Y _14603_/A vssd1 vssd1 vccd1 vccd1 _16129_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19819_ _19819_/A _19819_/B vssd1 vssd1 vccd1 vccd1 _19819_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_243_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22830_ _22830_/A vssd1 vssd1 vccd1 vccd1 _26396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22761_ _26366_/Q _22663_/X _22767_/S vssd1 vssd1 vccd1 vccd1 _22762_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24500_ _27028_/Q _24480_/X _24498_/Y _24499_/X vssd1 vssd1 vccd1 vccd1 _27028_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_225_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21712_ _16668_/B _21652_/X _20977_/A vssd1 vssd1 vccd1 vccd1 _21713_/C sky130_fd_sc_hd__o21ai_1
XFILLER_25_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25480_ _26881_/CLK _25480_/D vssd1 vssd1 vccd1 vccd1 _25480_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22692_ _22724_/A vssd1 vssd1 vccd1 vccd1 _22705_/S sky130_fd_sc_hd__buf_4
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24431_ _26305_/Q _24382_/X _24383_/X input218/X _24404_/X vssd1 vssd1 vccd1 vccd1
+ _24431_/X sky130_fd_sc_hd__a221o_1
X_21643_ _21641_/Y _21642_/X _21290_/A vssd1 vssd1 vccd1 vccd1 _21643_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27150_ _27227_/CLK _27150_/D vssd1 vssd1 vccd1 vccd1 _27150_/Q sky130_fd_sc_hd__dfxtp_4
X_24362_ _24781_/B vssd1 vssd1 vccd1 vccd1 _24548_/A sky130_fd_sc_hd__inv_2
X_21574_ _25493_/Q _21574_/B vssd1 vssd1 vccd1 vccd1 _21574_/X sky130_fd_sc_hd__or2_1
XFILLER_268_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26101_ _27266_/CLK _26101_/D vssd1 vssd1 vccd1 vccd1 _26101_/Q sky130_fd_sc_hd__dfxtp_2
X_23313_ _20529_/X _26597_/Q _23313_/S vssd1 vssd1 vccd1 vccd1 _23314_/A sky130_fd_sc_hd__mux2_1
X_20525_ _23712_/A vssd1 vssd1 vccd1 vccd1 _20525_/X sky130_fd_sc_hd__clkbuf_1
X_27081_ _27196_/CLK _27081_/D vssd1 vssd1 vccd1 vccd1 _27081_/Q sky130_fd_sc_hd__dfxtp_1
X_24293_ _26988_/Q _26987_/Q _24293_/C vssd1 vssd1 vccd1 vccd1 _24295_/B sky130_fd_sc_hd__and3_1
XFILLER_122_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26032_ _27267_/CLK _26032_/D vssd1 vssd1 vccd1 vccd1 _26032_/Q sky130_fd_sc_hd__dfxtp_1
X_23244_ _26566_/Q _23082_/X _23244_/S vssd1 vssd1 vccd1 vccd1 _23245_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20456_ _27163_/Q _27097_/Q vssd1 vssd1 vccd1 vccd1 _20457_/B sky130_fd_sc_hd__or2_1
XFILLER_192_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23175_ _26535_/Q _23085_/X _23183_/S vssd1 vssd1 vccd1 vccd1 _23176_/A sky130_fd_sc_hd__mux2_1
X_20387_ _27160_/Q _27094_/Q vssd1 vssd1 vccd1 vccd1 _20389_/A sky130_fd_sc_hd__or2_1
X_22126_ _26161_/Q _22110_/X _22125_/X _21878_/X vssd1 vssd1 vccd1 vccd1 _26161_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26934_ _27321_/CLK _26934_/D vssd1 vssd1 vccd1 vccd1 _26934_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22057_ _22103_/S vssd1 vssd1 vccd1 vccd1 _22066_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_102_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21008_ _21008_/A vssd1 vssd1 vccd1 vccd1 _25874_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26865_ _26929_/CLK _26865_/D vssd1 vssd1 vccd1 vccd1 _26865_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13830_ _25804_/Q _27238_/Q _16020_/S vssd1 vssd1 vccd1 vccd1 _13831_/B sky130_fd_sc_hd__mux2_1
X_25816_ _26917_/CLK _25816_/D vssd1 vssd1 vccd1 vccd1 _25816_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_247_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26796_ _26796_/CLK _26796_/D vssd1 vssd1 vccd1 vccd1 _26796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_251_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13761_ _15300_/A _13758_/X _13760_/X _15317_/A vssd1 vssd1 vccd1 vccd1 _13761_/X
+ sky130_fd_sc_hd__a211o_1
X_25747_ _26286_/CLK _25747_/D vssd1 vssd1 vccd1 vccd1 _25747_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22959_ _22959_/A vssd1 vssd1 vccd1 vccd1 _26454_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_209 _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15500_ _15515_/S vssd1 vssd1 vccd1 vccd1 _15501_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12712_ _15983_/S vssd1 vssd1 vccd1 vccd1 _13711_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_204_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16480_ _16477_/X _16478_/X _16480_/S vssd1 vssd1 vccd1 vccd1 _16481_/B sky130_fd_sc_hd__mux2_1
X_13692_ _15630_/A vssd1 vssd1 vccd1 vccd1 _16060_/S sky130_fd_sc_hd__buf_4
X_25678_ _26278_/CLK _25678_/D vssd1 vssd1 vccd1 vccd1 _25678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15431_ _15418_/X _15421_/X _15430_/Y vssd1 vssd1 vccd1 vccd1 _15431_/Y sky130_fd_sc_hd__o21bai_1
X_24629_ _24629_/A _24629_/B vssd1 vssd1 vccd1 vccd1 _24629_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18150_ _19709_/A _18227_/C vssd1 vssd1 vccd1 vccd1 _18150_/X sky130_fd_sc_hd__xor2_2
XFILLER_8_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15362_ _26348_/Q _26608_/Q _15374_/S vssd1 vssd1 vccd1 vccd1 _15362_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17101_ _25208_/B vssd1 vssd1 vccd1 vccd1 _20978_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14313_ _15516_/A _14309_/X _14312_/X _13311_/A vssd1 vssd1 vccd1 vccd1 _14313_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_196_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18081_ _18271_/B _17889_/X _18197_/S vssd1 vssd1 vccd1 vccd1 _18081_/X sky130_fd_sc_hd__mux2_1
X_15293_ _15596_/S vssd1 vssd1 vccd1 vccd1 _15834_/S sky130_fd_sc_hd__buf_6
XFILLER_157_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27279_ _27282_/CLK _27279_/D vssd1 vssd1 vccd1 vccd1 _27279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17032_ _17039_/A vssd1 vssd1 vccd1 vccd1 _17032_/X sky130_fd_sc_hd__buf_2
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14244_ _25800_/Q _27234_/Q _14245_/S vssd1 vssd1 vccd1 vccd1 _14244_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14175_ _13409_/A _14172_/X _14174_/X _13141_/A vssd1 vssd1 vccd1 vccd1 _14175_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13126_ _13126_/A vssd1 vssd1 vccd1 vccd1 _15538_/A sky130_fd_sc_hd__buf_2
XFILLER_112_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ _17772_/B _18978_/A _18981_/Y _18982_/X vssd1 vssd1 vccd1 vccd1 _18983_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_258_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_119_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25992_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13057_ _15895_/S vssd1 vssd1 vccd1 vccd1 _14001_/B sky130_fd_sc_hd__clkbuf_4
X_17934_ _17797_/B _17782_/B _17949_/S vssd1 vssd1 vccd1 vccd1 _17934_/X sky130_fd_sc_hd__mux2_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17865_ _18859_/A vssd1 vssd1 vccd1 vccd1 _18683_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19604_ _19943_/B vssd1 vssd1 vccd1 vccd1 _19604_/X sky130_fd_sc_hd__clkbuf_2
X_16816_ _16838_/A _16816_/B vssd1 vssd1 vccd1 vccd1 _16855_/B sky130_fd_sc_hd__or2_2
XFILLER_94_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17796_ _16289_/A _17794_/X _17795_/X vssd1 vssd1 vccd1 vccd1 _19237_/B sky130_fd_sc_hd__o21a_1
XFILLER_54_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19535_ _19525_/X _19030_/X _19534_/X _19528_/X vssd1 vssd1 vccd1 vccd1 _25648_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13959_ _26914_/Q _26398_/Q _16005_/S vssd1 vssd1 vccd1 vccd1 _13959_/X sky130_fd_sc_hd__mux2_1
X_16747_ _25675_/Q vssd1 vssd1 vccd1 vccd1 _22502_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19466_ _27036_/Q _18756_/X _19465_/X _18759_/X vssd1 vssd1 vccd1 vccd1 _19466_/X
+ sky130_fd_sc_hd__a22o_1
X_16678_ _20978_/B _16679_/B _17042_/A vssd1 vssd1 vccd1 vccd1 _16678_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_234_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18417_ _18201_/X _18196_/X _18489_/S vssd1 vssd1 vccd1 vccd1 _18417_/X sky130_fd_sc_hd__mux2_1
X_15629_ _15142_/A _15626_/X _15628_/X _15040_/A vssd1 vssd1 vccd1 vccd1 _15629_/X
+ sky130_fd_sc_hd__a211o_1
X_19397_ _25530_/Q _18743_/X _18744_/X _25562_/Q vssd1 vssd1 vccd1 vccd1 _19397_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_195_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18348_ _18071_/X _18061_/Y _18348_/S vssd1 vssd1 vccd1 vccd1 _18348_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18279_ _19078_/A _18230_/Y _18250_/X _18278_/X _18220_/X vssd1 vssd1 vccd1 vccd1
+ _18279_/X sky130_fd_sc_hd__a32o_1
XFILLER_147_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20310_ _20359_/A _20353_/A vssd1 vssd1 vccd1 vccd1 _20351_/A sky130_fd_sc_hd__xnor2_1
XFILLER_163_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21290_ _21290_/A vssd1 vssd1 vccd1 vccd1 _21290_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput50 dout0[16] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_2
Xinput61 dout0[26] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_2
Xinput72 dout0[36] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput83 dout0[46] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__clkbuf_1
X_20241_ _27154_/Q _27088_/Q vssd1 vssd1 vccd1 vccd1 _20241_/X sky130_fd_sc_hd__or2_1
XFILLER_192_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput94 dout0[56] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20172_ _17444_/D _18016_/A _20125_/A _20125_/B vssd1 vssd1 vccd1 vccd1 _20173_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_192_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24980_ _24625_/A _24902_/A _24966_/X vssd1 vssd1 vccd1 vccd1 _24980_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_269_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23931_ _23931_/A vssd1 vssd1 vccd1 vccd1 _26843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26650_ _27259_/CLK _26650_/D vssd1 vssd1 vccd1 vccd1 _26650_/Q sky130_fd_sc_hd__dfxtp_1
X_23862_ _23930_/S vssd1 vssd1 vccd1 vccd1 _23871_/S sky130_fd_sc_hd__clkbuf_4
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25601_ _25607_/CLK _25601_/D vssd1 vssd1 vccd1 vccd1 _25601_/Q sky130_fd_sc_hd__dfxtp_4
X_22813_ _26390_/Q _22739_/X _22815_/S vssd1 vssd1 vccd1 vccd1 _22814_/A sky130_fd_sc_hd__mux2_1
X_26581_ _27321_/CLK _26581_/D vssd1 vssd1 vccd1 vccd1 _26581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_272_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23793_ _23690_/X _26781_/Q _23799_/S vssd1 vssd1 vccd1 vccd1 _23794_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25532_ _26257_/CLK _25532_/D vssd1 vssd1 vccd1 vccd1 _25532_/Q sky130_fd_sc_hd__dfxtp_1
X_22744_ _22744_/A vssd1 vssd1 vccd1 vccd1 _26359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25463_ _23785_/X _27326_/Q _25463_/S vssd1 vssd1 vccd1 vccd1 _25464_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22675_ _23718_/A vssd1 vssd1 vccd1 vccd1 _22675_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_179_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27202_ _27230_/CLK _27202_/D vssd1 vssd1 vccd1 vccd1 _27202_/Q sky130_fd_sc_hd__dfxtp_1
X_24414_ _24434_/A _24572_/A vssd1 vssd1 vccd1 vccd1 _24414_/Y sky130_fd_sc_hd__nand2_1
XFILLER_157_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21626_ _21626_/A vssd1 vssd1 vccd1 vccd1 _21626_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25394_ _25450_/A vssd1 vssd1 vccd1 vccd1 _25463_/S sky130_fd_sc_hd__buf_4
XFILLER_139_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27133_ _27133_/CLK _27133_/D vssd1 vssd1 vccd1 vccd1 _27133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24345_ _21203_/A _25495_/Q _17694_/Y vssd1 vssd1 vccd1 vccd1 _24347_/C sky130_fd_sc_hd__a21o_1
XFILLER_139_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21557_ _21551_/Y _21555_/X _21556_/X vssd1 vssd1 vccd1 vccd1 _21557_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20508_ _23699_/A vssd1 vssd1 vccd1 vccd1 _20508_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_27064_ _27160_/CLK _27064_/D vssd1 vssd1 vccd1 vccd1 _27064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24276_ _24285_/A _24276_/B _24278_/B vssd1 vssd1 vccd1 vccd1 _26982_/D sky130_fd_sc_hd__nor3_1
X_21488_ _21552_/A vssd1 vssd1 vccd1 vccd1 _21488_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26015_ _26531_/CLK _26015_/D vssd1 vssd1 vccd1 vccd1 _26015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23227_ _26558_/Q _23057_/X _23233_/S vssd1 vssd1 vccd1 vccd1 _23228_/A sky130_fd_sc_hd__mux2_1
X_20439_ _20429_/Y _20430_/X _20438_/X _20712_/A _19651_/X vssd1 vssd1 vccd1 vccd1
+ _20439_/X sky130_fd_sc_hd__a221o_1
XFILLER_134_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23158_ _23158_/A vssd1 vssd1 vccd1 vccd1 _26527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22109_ _22200_/A vssd1 vssd1 vccd1 vccd1 _22152_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15980_ _26632_/Q _26728_/Q _15980_/S vssd1 vssd1 vccd1 vccd1 _15980_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23089_ _23562_/A vssd1 vssd1 vccd1 vccd1 _23089_/X sky130_fd_sc_hd__buf_2
XFILLER_103_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14931_ _19408_/A vssd1 vssd1 vccd1 vccd1 _14931_/Y sky130_fd_sc_hd__inv_2
XTAP_5654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26917_ _26917_/CLK _26917_/D vssd1 vssd1 vccd1 vccd1 _26917_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14862_ _14948_/S _14857_/X _14861_/X _14662_/A vssd1 vssd1 vccd1 vccd1 _14862_/X
+ sky130_fd_sc_hd__a211o_1
X_17650_ _17650_/A _17650_/B vssd1 vssd1 vccd1 vccd1 _25595_/D sky130_fd_sc_hd__nor2_1
XFILLER_275_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26848_ _26880_/CLK _26848_/D vssd1 vssd1 vccd1 vccd1 _26848_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13813_ _13835_/A vssd1 vssd1 vccd1 vccd1 _13813_/X sky130_fd_sc_hd__clkbuf_2
X_16601_ _20798_/B _16604_/A _16639_/B vssd1 vssd1 vccd1 vccd1 _16989_/A sky130_fd_sc_hd__and3_2
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17581_ _17534_/X _17592_/B _14136_/X _17536_/X _25914_/Q vssd1 vssd1 vccd1 vccd1
+ _17581_/Y sky130_fd_sc_hd__o32ai_4
XFILLER_217_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26779_ _26843_/CLK _26779_/D vssd1 vssd1 vccd1 vccd1 _26779_/Q sky130_fd_sc_hd__dfxtp_1
X_14793_ _14793_/A vssd1 vssd1 vccd1 vccd1 _14794_/A sky130_fd_sc_hd__buf_2
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19320_ _25624_/Q _19153_/X _19319_/X _19185_/X vssd1 vssd1 vccd1 vccd1 _25624_/D
+ sky130_fd_sc_hd__o211a_1
X_16532_ _16530_/X _16531_/X _16540_/S vssd1 vssd1 vccd1 vccd1 _16532_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13744_ _14025_/A _13923_/B _14025_/B _13744_/D vssd1 vssd1 vccd1 vccd1 _13744_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_232_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19251_ _19317_/A _19251_/B vssd1 vssd1 vccd1 vccd1 _19251_/Y sky130_fd_sc_hd__nand2_1
X_16463_ _16463_/A vssd1 vssd1 vccd1 vccd1 _16463_/X sky130_fd_sc_hd__clkbuf_4
X_13675_ _26529_/Q _26137_/Q _13675_/S vssd1 vssd1 vccd1 vccd1 _13675_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18202_ _18202_/A vssd1 vssd1 vccd1 vccd1 _18345_/S sky130_fd_sc_hd__clkbuf_2
X_15414_ _15414_/A vssd1 vssd1 vccd1 vccd1 _16361_/S sky130_fd_sc_hd__clkbuf_4
XPHY_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19182_ _19317_/A _19182_/B vssd1 vssd1 vccd1 vccd1 _19182_/Y sky130_fd_sc_hd__nand2_1
XPHY_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16394_ _15044_/X _16392_/X _16393_/X vssd1 vssd1 vccd1 vccd1 _16394_/X sky130_fd_sc_hd__o21a_1
XFILLER_85_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18133_ _18555_/A _18100_/X _18132_/X vssd1 vssd1 vccd1 vccd1 _18133_/X sky130_fd_sc_hd__a21o_4
X_15345_ _15345_/A _15345_/B vssd1 vssd1 vccd1 vccd1 _15345_/X sky130_fd_sc_hd__or2_1
XFILLER_184_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18064_ _18062_/X _18063_/X _18254_/A vssd1 vssd1 vccd1 vccd1 _18064_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15276_ _26118_/Q _26019_/Q _15276_/S vssd1 vssd1 vccd1 vccd1 _15276_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17015_ _17042_/A vssd1 vssd1 vccd1 vccd1 _17015_/X sky130_fd_sc_hd__clkbuf_4
X_14227_ _13806_/X _14223_/X _14226_/X _13543_/A vssd1 vssd1 vccd1 vccd1 _14227_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_208_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14158_ _14176_/S vssd1 vssd1 vccd1 vccd1 _15902_/S sky130_fd_sc_hd__buf_4
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13109_ _13717_/A vssd1 vssd1 vccd1 vccd1 _14708_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_140_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14089_ _14084_/X _14088_/X _14089_/S vssd1 vssd1 vccd1 vccd1 _14089_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18966_ _18723_/X _18962_/X _18965_/X _18884_/X vssd1 vssd1 vccd1 vccd1 _18967_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_224_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17917_ _18349_/S vssd1 vssd1 vccd1 vccd1 _18492_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_255_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18897_ _17920_/X _18492_/B _18896_/X _18547_/S vssd1 vssd1 vccd1 vccd1 _18936_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_239_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17848_ _19355_/A _19355_/B _19355_/C _19356_/A vssd1 vssd1 vccd1 vccd1 _19389_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_27_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_87_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25598_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17779_ _17779_/A vssd1 vssd1 vccd1 vccd1 _17779_/Y sky130_fd_sc_hd__inv_2
XFILLER_282_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19518_ _19512_/X _18702_/X _19517_/X _19515_/X vssd1 vssd1 vccd1 vccd1 _25641_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_223_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20790_ _22472_/B _20973_/B _20790_/C vssd1 vssd1 vccd1 vccd1 _20791_/A sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_16_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27282_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_223_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_540 _25737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_551 _25925_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19449_ _19449_/A _25161_/A vssd1 vssd1 vccd1 vccd1 _19449_/Y sky130_fd_sc_hd__nand2_1
XFILLER_250_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22460_ _22460_/A vssd1 vssd1 vccd1 vccd1 _22470_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_194_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21411_ _21354_/X _21355_/X _21410_/Y _21386_/X vssd1 vssd1 vccd1 vccd1 _21411_/X
+ sky130_fd_sc_hd__a31o_1
X_22391_ _22387_/B _22362_/B _22381_/X _22385_/X _22390_/Y vssd1 vssd1 vccd1 vccd1
+ _22391_/X sky130_fd_sc_hd__o221a_1
XFILLER_120_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24130_ _24130_/A vssd1 vssd1 vccd1 vccd1 _26931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21342_ _21544_/A vssd1 vssd1 vccd1 vccd1 _21342_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24061_ _24061_/A vssd1 vssd1 vccd1 vccd1 _24070_/S sky130_fd_sc_hd__buf_6
X_21273_ _21273_/A _21273_/B vssd1 vssd1 vccd1 vccd1 _21273_/Y sky130_fd_sc_hd__nor2_2
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23012_ _23012_/A vssd1 vssd1 vccd1 vccd1 _26477_/D sky130_fd_sc_hd__clkbuf_1
X_20224_ _22513_/A _20078_/X _20213_/X _20221_/Y _20223_/X vssd1 vssd1 vccd1 vccd1
+ _25680_/D sky130_fd_sc_hd__o221a_1
XFILLER_270_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20155_ _27119_/Q _20079_/X _20112_/X _20154_/Y vssd1 vssd1 vccd1 vccd1 _20155_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24963_ _27154_/Q _24957_/X _24962_/Y vssd1 vssd1 vccd1 vccd1 _27154_/D sky130_fd_sc_hd__o21a_1
X_20086_ _20040_/X _20082_/Y _20085_/X vssd1 vssd1 vccd1 vccd1 _20086_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26702_ _27308_/CLK _26702_/D vssd1 vssd1 vccd1 vccd1 _26702_/Q sky130_fd_sc_hd__dfxtp_2
X_23914_ _23914_/A vssd1 vssd1 vccd1 vccd1 _26835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24894_ _20701_/A _19724_/X _24768_/Y _24782_/X vssd1 vssd1 vccd1 vccd1 _24894_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26633_ _27304_/CLK _26633_/D vssd1 vssd1 vccd1 vccd1 _26633_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23845_ _23845_/A vssd1 vssd1 vccd1 vccd1 _23854_/S sky130_fd_sc_hd__buf_6
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26564_ _26920_/CLK _26564_/D vssd1 vssd1 vccd1 vccd1 _26564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23776_ _23776_/A vssd1 vssd1 vccd1 vccd1 _23776_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20988_ _16681_/Y _25867_/D vssd1 vssd1 vccd1 vccd1 _20989_/A sky130_fd_sc_hd__and2b_1
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25515_ _25518_/CLK _25515_/D vssd1 vssd1 vccd1 vccd1 _25515_/Q sky130_fd_sc_hd__dfxtp_1
X_22727_ _23770_/A vssd1 vssd1 vccd1 vccd1 _22727_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26495_ _27272_/CLK _26495_/D vssd1 vssd1 vccd1 vccd1 _26495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25446_ _23760_/X _27318_/Q _25448_/S vssd1 vssd1 vccd1 vccd1 _25447_/A sky130_fd_sc_hd__mux2_1
X_13460_ _14560_/S vssd1 vssd1 vccd1 vccd1 _16031_/S sky130_fd_sc_hd__buf_2
X_22658_ _22658_/A vssd1 vssd1 vccd1 vccd1 _26332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21609_ _25963_/Q _21573_/X _21608_/Y _21597_/X vssd1 vssd1 vccd1 vccd1 _25963_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_199_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13391_ _13916_/A _13923_/B _13397_/B _13391_/D vssd1 vssd1 vccd1 vccd1 _13391_/X
+ sky130_fd_sc_hd__or4_2
X_25377_ _25377_/A vssd1 vssd1 vccd1 vccd1 _27287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_279_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22589_ _26311_/Q _22591_/B vssd1 vssd1 vccd1 vccd1 _22589_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15130_ _17787_/A _17786_/A vssd1 vssd1 vccd1 vccd1 _19294_/S sky130_fd_sc_hd__nor2_2
X_27116_ _27117_/CLK _27116_/D vssd1 vssd1 vccd1 vccd1 _27116_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24328_ _27001_/Q _24331_/C vssd1 vssd1 vccd1 vccd1 _24329_/B sky130_fd_sc_hd__and2_1
XFILLER_182_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27047_ _27062_/CLK _27047_/D vssd1 vssd1 vccd1 vccd1 _27047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15061_ _16328_/A vssd1 vssd1 vccd1 vccd1 _16405_/A sky130_fd_sc_hd__clkbuf_2
X_24259_ _24285_/A _24259_/B _24260_/B vssd1 vssd1 vccd1 vccd1 _26976_/D sky130_fd_sc_hd__nor3_1
XFILLER_107_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14012_ _25875_/Q _14173_/B vssd1 vssd1 vccd1 vccd1 _14012_/X sky130_fd_sc_hd__or2_1
XFILLER_49_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18820_ _27146_/Q _19367_/B vssd1 vssd1 vccd1 vccd1 _18820_/X sky130_fd_sc_hd__or2_1
XFILLER_122_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18751_ _18815_/A vssd1 vssd1 vccd1 vccd1 _18751_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15963_ _13402_/A _15960_/X _15962_/X _13126_/A vssd1 vssd1 vccd1 vccd1 _15963_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput240 localMemory_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input240/X sky130_fd_sc_hd__buf_6
XTAP_5462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput251 localMemory_wb_stb_i vssd1 vssd1 vccd1 vccd1 _21654_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17702_ _17691_/A _17443_/A _17701_/X vssd1 vssd1 vccd1 vccd1 _17736_/C sky130_fd_sc_hd__a21oi_1
Xinput262 manufacturerID[8] vssd1 vssd1 vccd1 vccd1 input262/X sky130_fd_sc_hd__clkbuf_2
X_14914_ _26937_/Q _26421_/Q _14996_/S vssd1 vssd1 vccd1 vccd1 _14914_/X sky130_fd_sc_hd__mux2_1
Xinput273 partID[3] vssd1 vssd1 vccd1 vccd1 input273/X sky130_fd_sc_hd__clkbuf_1
XTAP_5484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15894_ _27308_/Q _26565_/Q _15895_/S vssd1 vssd1 vccd1 vccd1 _15894_/X sky130_fd_sc_hd__mux2_1
X_18682_ _18682_/A vssd1 vssd1 vccd1 vccd1 _18682_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput284 wb_rst_i vssd1 vssd1 vccd1 vccd1 _20487_/B sky130_fd_sc_hd__buf_12
XFILLER_91_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ _17633_/A _17633_/B vssd1 vssd1 vccd1 vccd1 _25590_/D sky130_fd_sc_hd__nor2_1
XFILLER_263_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14845_ _27324_/Q _26581_/Q _14960_/B vssd1 vssd1 vccd1 vccd1 _14845_/X sky130_fd_sc_hd__mux2_1
XFILLER_252_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14776_ _16521_/A _14776_/B _14776_/C vssd1 vssd1 vccd1 vccd1 _14776_/Y sky130_fd_sc_hd__nor3_1
X_17564_ _17635_/A vssd1 vssd1 vccd1 vccd1 _17564_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_189_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19303_ _27031_/Q _18449_/X _19302_/X _18821_/X vssd1 vssd1 vccd1 vccd1 _19303_/X
+ sky130_fd_sc_hd__a22o_1
X_13727_ _27303_/Q _26560_/Q _15464_/B vssd1 vssd1 vccd1 vccd1 _13727_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16515_ _16513_/X _26715_/Q _26843_/Q _16526_/S _14773_/X vssd1 vssd1 vccd1 vccd1
+ _16515_/X sky130_fd_sc_hd__a221o_1
XFILLER_32_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17495_ _17706_/A vssd1 vssd1 vccd1 vccd1 _17704_/S sky130_fd_sc_hd__buf_2
XFILLER_177_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19234_ _19234_/A _19234_/B _19234_/C vssd1 vssd1 vccd1 vccd1 _19234_/X sky130_fd_sc_hd__or3_4
X_13658_ _16021_/S vssd1 vssd1 vccd1 vccd1 _16020_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_31_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16446_ _14759_/A _16442_/X _16445_/X _14779_/A vssd1 vssd1 vccd1 vccd1 _16446_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_223_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16377_ _26871_/Q _25785_/Q _16377_/S vssd1 vssd1 vccd1 vccd1 _16377_/X sky130_fd_sc_hd__mux2_1
X_19165_ _27123_/Q _18812_/X _19163_/X _19164_/X vssd1 vssd1 vccd1 vccd1 _19165_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_219_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13589_ _27272_/Q _26465_/Q _13589_/S vssd1 vssd1 vccd1 vccd1 _13589_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18116_ _18116_/A _18116_/B vssd1 vssd1 vccd1 vccd1 _18119_/B sky130_fd_sc_hd__or2_1
X_15328_ _27285_/Q _26478_/Q _15414_/A vssd1 vssd1 vccd1 vccd1 _15328_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19096_ _26961_/Q _18461_/A _18463_/A _26993_/Q vssd1 vssd1 vccd1 vccd1 _19096_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_145_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_134_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27166_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18047_ _18058_/S vssd1 vssd1 vccd1 vccd1 _18062_/S sky130_fd_sc_hd__clkbuf_2
X_15259_ _25819_/Q _16387_/S _16401_/S _15258_/X vssd1 vssd1 vccd1 vccd1 _15259_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19998_ _19999_/A _19999_/B _19999_/C vssd1 vssd1 vccd1 vccd1 _19998_/X sky130_fd_sc_hd__o21a_1
XFILLER_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18949_ _27215_/Q _18949_/B vssd1 vssd1 vccd1 vccd1 _18949_/X sky130_fd_sc_hd__and2_1
XFILLER_255_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21960_ _21960_/A vssd1 vssd1 vccd1 vccd1 _26095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20911_ _25841_/Q _20910_/X _20917_/S vssd1 vssd1 vccd1 vccd1 _20912_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21891_ _21959_/S vssd1 vssd1 vccd1 vccd1 _21900_/S sky130_fd_sc_hd__buf_2
XFILLER_282_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23630_ _26723_/Q _23533_/X _23634_/S vssd1 vssd1 vccd1 vccd1 _23631_/A sky130_fd_sc_hd__mux2_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20842_ _25817_/Q vssd1 vssd1 vccd1 vccd1 _20843_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_42_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23561_ _23561_/A vssd1 vssd1 vccd1 vccd1 _26699_/D sky130_fd_sc_hd__clkbuf_1
X_20773_ _20773_/A vssd1 vssd1 vccd1 vccd1 _25782_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_370 _17062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25300_ _23757_/X _27253_/Q _25304_/S vssd1 vssd1 vccd1 vccd1 _25301_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22512_ _22512_/A vssd1 vssd1 vccd1 vccd1 _26280_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_381 _16774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26280_ _26282_/CLK _26280_/D vssd1 vssd1 vccd1 vccd1 _26280_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_392 _17033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23492_ _23492_/A vssd1 vssd1 vccd1 vccd1 _26676_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25231_ _24988_/X _19623_/X _24771_/X _24739_/B _25219_/X vssd1 vssd1 vccd1 vccd1
+ _25231_/X sky130_fd_sc_hd__a221o_1
XFILLER_50_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22443_ _26201_/Q _22432_/X _22440_/X _22442_/X vssd1 vssd1 vccd1 vccd1 _26249_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_210_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25162_ _22533_/A _25119_/X _25139_/A _25161_/Y _25024_/A vssd1 vssd1 vccd1 vccd1
+ _25162_/X sky130_fd_sc_hd__a221o_1
X_22374_ _22377_/A _22374_/B vssd1 vssd1 vccd1 vccd1 _22375_/A sky130_fd_sc_hd__and2_1
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24113_ _24113_/A vssd1 vssd1 vccd1 vccd1 _26923_/D sky130_fd_sc_hd__clkbuf_1
X_21325_ _20639_/A _21278_/X _21279_/X _21324_/X vssd1 vssd1 vccd1 vccd1 _21325_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25093_ _22505_/A _25092_/X _25087_/X _18968_/B _25079_/X vssd1 vssd1 vccd1 vccd1
+ _25093_/X sky130_fd_sc_hd__a221o_1
XFILLER_191_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24044_ _26893_/Q _23565_/X _24048_/S vssd1 vssd1 vccd1 vccd1 _24045_/A sky130_fd_sc_hd__mux2_1
X_21256_ _26062_/Q _17482_/B _21866_/B _21544_/A _21255_/X vssd1 vssd1 vccd1 vccd1
+ _21256_/X sky130_fd_sc_hd__a311o_1
XFILLER_104_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20207_ _20206_/B _20206_/C _20206_/A vssd1 vssd1 vccd1 vccd1 _20260_/B sky130_fd_sc_hd__o21a_1
X_21187_ _25933_/Q _21112_/A _21113_/A input34/X vssd1 vssd1 vccd1 vccd1 _21188_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_145_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20138_ _19894_/X _20137_/X _19902_/X vssd1 vssd1 vccd1 vccd1 _20138_/X sky130_fd_sc_hd__a21o_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25995_ _27156_/CLK _25995_/D vssd1 vssd1 vccd1 vccd1 _25995_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24946_ _24590_/A _24941_/X _24938_/X vssd1 vssd1 vccd1 vccd1 _24946_/Y sky130_fd_sc_hd__a21oi_1
X_12960_ _20868_/A _12996_/A vssd1 vssd1 vccd1 vccd1 _21888_/B sky130_fd_sc_hd__or2b_1
X_20069_ _27148_/Q _27082_/Q vssd1 vssd1 vccd1 vccd1 _20069_/Y sky130_fd_sc_hd__nand2_1
XINSDIODE2_30 _19285_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_41 _19441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_52 _20641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_63 _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_74 _20681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _12891_/A vssd1 vssd1 vccd1 vccd1 _12892_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_24877_ _24877_/A vssd1 vssd1 vccd1 vccd1 _24890_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_85 _23712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_96 _21385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14700_/S vssd1 vssd1 vccd1 vccd1 _16499_/S sky130_fd_sc_hd__clkbuf_2
X_23828_ _23741_/X _26797_/Q _23832_/S vssd1 vssd1 vccd1 vccd1 _23829_/A sky130_fd_sc_hd__mux2_1
X_26616_ _27324_/CLK _26616_/D vssd1 vssd1 vccd1 vccd1 _26616_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26547_ _26903_/CLK _26547_/D vssd1 vssd1 vccd1 vccd1 _26547_/Q sky130_fd_sc_hd__dfxtp_1
X_14561_ _15615_/S _16581_/B _17807_/A vssd1 vssd1 vccd1 vccd1 _16580_/A sky130_fd_sc_hd__and3_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23759_ _23759_/A vssd1 vssd1 vccd1 vccd1 _26770_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _13512_/A vssd1 vssd1 vccd1 vccd1 _15606_/A sky130_fd_sc_hd__buf_4
X_16300_ _16386_/S _16297_/X _16299_/X _15020_/A vssd1 vssd1 vccd1 vccd1 _16300_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17280_ _17278_/X _17282_/C _17279_/Y vssd1 vssd1 vccd1 vccd1 _25514_/D sky130_fd_sc_hd__o21a_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14407_/X _14490_/X _14491_/X _13557_/A vssd1 vssd1 vccd1 vccd1 _14492_/X
+ sky130_fd_sc_hd__o211a_1
X_26478_ _26611_/CLK _26478_/D vssd1 vssd1 vccd1 vccd1 _26478_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16231_ _27318_/Q _26575_/Q _16235_/S vssd1 vssd1 vccd1 vccd1 _16231_/X sky130_fd_sc_hd__mux2_1
X_13443_ _12745_/A _13441_/X _13442_/X vssd1 vssd1 vccd1 vccd1 _13443_/X sky130_fd_sc_hd__o21a_1
X_25429_ _23734_/X _27310_/Q _25437_/S vssd1 vssd1 vccd1 vccd1 _25430_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16162_ _15265_/X _16161_/X _14694_/A _12703_/A vssd1 vssd1 vccd1 vccd1 _16162_/X
+ sky130_fd_sc_hd__o211a_1
X_13374_ _14481_/B vssd1 vssd1 vccd1 vccd1 _14317_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15113_ _14764_/A _15108_/X _15112_/X _12756_/A vssd1 vssd1 vccd1 vccd1 _15117_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16093_ _16093_/A _16093_/B vssd1 vssd1 vccd1 vccd1 _16093_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15044_ _15044_/A vssd1 vssd1 vccd1 vccd1 _15044_/X sky130_fd_sc_hd__buf_2
X_19921_ _19887_/A _19779_/A _19883_/X _20119_/B _19885_/Y vssd1 vssd1 vccd1 vccd1
+ _19976_/C sky130_fd_sc_hd__o221ai_4
XFILLER_269_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_19852_ _19852_/A _19976_/B vssd1 vssd1 vccd1 vccd1 _19980_/A sky130_fd_sc_hd__xor2_1
XFILLER_214_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18803_ _19583_/A _18803_/B _18803_/C _18803_/D vssd1 vssd1 vccd1 vccd1 _18803_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_110_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19783_ _27106_/Q _19722_/X _19761_/X _19782_/Y vssd1 vssd1 vccd1 vccd1 _19783_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_284_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16995_ _22483_/A _16988_/X _16990_/X _18424_/A vssd1 vssd1 vccd1 vccd1 _16995_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_95_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18734_ _18734_/A vssd1 vssd1 vccd1 vccd1 _18734_/X sky130_fd_sc_hd__buf_2
XTAP_5270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15946_ _15921_/Y _15929_/Y _13466_/A _15945_/Y vssd1 vssd1 vccd1 vccd1 _15946_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_5281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18665_ _18435_/X _18663_/X _18666_/B vssd1 vssd1 vccd1 vccd1 _18665_/X sky130_fd_sc_hd__a21o_1
XFILLER_237_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ _12951_/X _15875_/X _15876_/X vssd1 vssd1 vccd1 vccd1 _15877_/X sky130_fd_sc_hd__o21a_1
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17616_ _17634_/A vssd1 vssd1 vccd1 vccd1 _17633_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14828_ _14724_/X _14620_/Y _14824_/X _14827_/X vssd1 vssd1 vccd1 vccd1 _19442_/A
+ sky130_fd_sc_hd__a211o_4
X_18596_ _16732_/X _19354_/B _18595_/X vssd1 vssd1 vccd1 vccd1 _18596_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_224_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17547_ _25570_/Q _17529_/X _17540_/X _17546_/Y vssd1 vssd1 vccd1 vccd1 _17548_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14759_ _14759_/A vssd1 vssd1 vccd1 vccd1 _14760_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_189_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17478_ _26260_/Q _26259_/Q _26258_/Q vssd1 vssd1 vccd1 vccd1 _17478_/X sky130_fd_sc_hd__or3_2
XFILLER_220_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19217_ _25621_/Q _19153_/X _19216_/X _19185_/X vssd1 vssd1 vccd1 vccd1 _25621_/D
+ sky130_fd_sc_hd__o211a_1
X_16429_ _14743_/A _25785_/Q _15228_/S _26871_/Q _16360_/S vssd1 vssd1 vccd1 vccd1
+ _16429_/X sky130_fd_sc_hd__o221a_1
XFILLER_9_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19148_ _19179_/B _19148_/B vssd1 vssd1 vccd1 vccd1 _19148_/X sky130_fd_sc_hd__or2_2
XFILLER_117_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19079_ _18716_/X _19053_/X _19077_/X _19078_/X vssd1 vssd1 vccd1 vccd1 _19079_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_145_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21110_ _21118_/A _21110_/B vssd1 vssd1 vccd1 vccd1 _21111_/A sky130_fd_sc_hd__or2_1
XFILLER_117_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22090_ _22090_/A vssd1 vssd1 vccd1 vccd1 _22099_/S sky130_fd_sc_hd__buf_6
XFILLER_114_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21041_ _21041_/A vssd1 vssd1 vccd1 vccd1 _25889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24800_ _24798_/Y _24799_/X _24796_/X vssd1 vssd1 vccd1 vccd1 _27105_/D sky130_fd_sc_hd__a21oi_1
X_25780_ _26610_/CLK _25780_/D vssd1 vssd1 vccd1 vccd1 _25780_/Q sky130_fd_sc_hd__dfxtp_1
X_22992_ _22992_/A vssd1 vssd1 vccd1 vccd1 _26468_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26880_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24731_ _24742_/A _24731_/B vssd1 vssd1 vccd1 vccd1 _27089_/D sky130_fd_sc_hd__nor2_1
X_21943_ _21943_/A vssd1 vssd1 vccd1 vccd1 _26087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24662_ _24678_/A _24662_/B vssd1 vssd1 vccd1 vccd1 _27073_/D sky130_fd_sc_hd__nor2_1
X_21874_ _21874_/A _21885_/B vssd1 vssd1 vccd1 vccd1 _21874_/X sky130_fd_sc_hd__or2_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26401_ _26433_/CLK _26401_/D vssd1 vssd1 vccd1 vccd1 _26401_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23613_ _23669_/A vssd1 vssd1 vccd1 vccd1 _23682_/S sky130_fd_sc_hd__buf_4
X_20825_ _20825_/A vssd1 vssd1 vccd1 vccd1 _25808_/D sky130_fd_sc_hd__clkbuf_1
X_24593_ _24619_/A vssd1 vssd1 vccd1 vccd1 _24593_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26332_ _26462_/CLK _26332_/D vssd1 vssd1 vccd1 vccd1 _26332_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_168_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23544_ _26694_/Q _23542_/X _23556_/S vssd1 vssd1 vccd1 vccd1 _23545_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20756_ _20756_/A vssd1 vssd1 vccd1 vccd1 _25774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26263_ _26264_/CLK _26263_/D vssd1 vssd1 vccd1 vccd1 _26263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23475_ _23475_/A vssd1 vssd1 vccd1 vccd1 _26668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20687_ _20687_/A _20687_/B vssd1 vssd1 vccd1 vccd1 _20687_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25214_ _25214_/A vssd1 vssd1 vccd1 vccd1 _25214_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22426_ _26195_/Q _22418_/X _22425_/X _22348_/X vssd1 vssd1 vccd1 vccd1 _26243_/D
+ sky130_fd_sc_hd__o211a_1
X_26194_ _26297_/CLK _26194_/D vssd1 vssd1 vccd1 vccd1 _26194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25145_ _22526_/A _24639_/A _25139_/X _16575_/C _12781_/X vssd1 vssd1 vccd1 vccd1
+ _25145_/X sky130_fd_sc_hd__a221o_1
XFILLER_109_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22357_ _22357_/A vssd1 vssd1 vccd1 vccd1 _26231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_276_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21308_ _25940_/Q _21202_/X _21307_/Y _21262_/X vssd1 vssd1 vccd1 vccd1 _25940_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_151_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13090_ _13616_/S vssd1 vssd1 vccd1 vccd1 _15630_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_191_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25076_ _20656_/A _25059_/X _25075_/X vssd1 vssd1 vccd1 vccd1 _25076_/Y sky130_fd_sc_hd__o21ai_1
X_22288_ _22288_/A vssd1 vssd1 vccd1 vccd1 _22288_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24027_ _24027_/A vssd1 vssd1 vccd1 vccd1 _26885_/D sky130_fd_sc_hd__clkbuf_1
X_21239_ _21309_/A vssd1 vssd1 vccd1 vccd1 _21273_/A sky130_fd_sc_hd__buf_6
XFILLER_277_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15800_ _26858_/Q _25772_/Q _15800_/S vssd1 vssd1 vccd1 vccd1 _15800_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13992_ _13884_/S _13990_/X _13991_/X vssd1 vssd1 vccd1 vccd1 _13992_/X sky130_fd_sc_hd__o21a_1
X_16780_ _25687_/Q vssd1 vssd1 vccd1 vccd1 _22528_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25978_ _27022_/CLK _25978_/D vssd1 vssd1 vccd1 vccd1 _25978_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_120_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15731_ _26923_/Q _15805_/S vssd1 vssd1 vccd1 vccd1 _15731_/X sky130_fd_sc_hd__or2_1
X_12943_ _12868_/Y _12941_/Y _14325_/S vssd1 vssd1 vccd1 vccd1 _12943_/Y sky130_fd_sc_hd__a21oi_2
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24929_ _19870_/A _24927_/X _24928_/Y vssd1 vssd1 vccd1 vccd1 _27141_/D sky130_fd_sc_hd__o21a_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18450_ _18445_/X _18448_/X _18449_/X vssd1 vssd1 vccd1 vccd1 _18450_/X sky130_fd_sc_hd__a21o_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12874_ _14407_/A _14486_/A vssd1 vssd1 vccd1 vccd1 _14411_/A sky130_fd_sc_hd__nand2_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _26636_/Q _26732_/Q _15662_/S vssd1 vssd1 vccd1 vccd1 _15663_/B sky130_fd_sc_hd__mux2_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _25552_/Q _17401_/B vssd1 vssd1 vccd1 vccd1 _17408_/C sky130_fd_sc_hd__and2_1
XFILLER_27_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _15135_/A vssd1 vssd1 vccd1 vccd1 _14613_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_261_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15593_ _16195_/S _15590_/X _15592_/X _13305_/A vssd1 vssd1 vccd1 vccd1 _15593_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18381_ _18381_/A vssd1 vssd1 vccd1 vccd1 _18382_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17332_ _17332_/A _17332_/B _17333_/B vssd1 vssd1 vccd1 vccd1 _25530_/D sky130_fd_sc_hd__nor3_1
X_14544_ _26908_/Q _26392_/Q _14544_/S vssd1 vssd1 vccd1 vccd1 _14544_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17263_ _25508_/Q _25509_/Q _17263_/C vssd1 vssd1 vccd1 vccd1 _17265_/B sky130_fd_sc_hd__and3_1
X_14475_ _13250_/A _26877_/Q _26749_/Q _13657_/A _12731_/A vssd1 vssd1 vccd1 vccd1
+ _14475_/X sky130_fd_sc_hd__a221o_1
XFILLER_201_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19002_ _25741_/Q _19037_/C vssd1 vssd1 vccd1 vccd1 _19002_/Y sky130_fd_sc_hd__xnor2_2
X_13426_ _13420_/X _13421_/X _13698_/A vssd1 vssd1 vccd1 vccd1 _13426_/X sky130_fd_sc_hd__mux2_1
X_16214_ _25621_/Q _14597_/A _16213_/X _14618_/A vssd1 vssd1 vccd1 vccd1 _23584_/A
+ sky130_fd_sc_hd__o22a_4
X_17194_ _14662_/X _17190_/X _17193_/X _17188_/X vssd1 vssd1 vccd1 vccd1 _25490_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16145_ _27284_/Q _26477_/Q _16163_/S vssd1 vssd1 vccd1 vccd1 _16145_/X sky130_fd_sc_hd__mux2_1
X_13357_ _15484_/S vssd1 vssd1 vccd1 vccd1 _15299_/S sky130_fd_sc_hd__buf_6
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16076_ _15645_/S _16075_/X _13703_/A vssd1 vssd1 vccd1 vccd1 _16076_/X sky130_fd_sc_hd__a21o_1
X_13288_ _15582_/A vssd1 vssd1 vccd1 vccd1 _16087_/S sky130_fd_sc_hd__buf_6
XFILLER_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19904_ _22489_/A _19876_/X _19893_/X _19903_/X _19874_/X vssd1 vssd1 vccd1 vccd1
+ _25669_/D sky130_fd_sc_hd__o221a_1
X_15027_ _25823_/Q _15014_/S _16386_/S _15026_/X vssd1 vssd1 vccd1 vccd1 _15027_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19835_ _25666_/Q _19834_/C _25667_/Q vssd1 vssd1 vccd1 vccd1 _19835_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19766_ _19766_/A vssd1 vssd1 vccd1 vccd1 _19766_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_256_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16978_ _16983_/A _16983_/B _16978_/C vssd1 vssd1 vccd1 vccd1 _16978_/X sky130_fd_sc_hd__and3_1
XFILLER_256_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput4 coreIndex[3] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_4
XFILLER_272_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18717_ _19003_/A _18716_/X _18010_/X _24986_/A vssd1 vssd1 vccd1 vccd1 _19287_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_283_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15929_ _15925_/X _15928_/X _14807_/A vssd1 vssd1 vccd1 vccd1 _15929_/Y sky130_fd_sc_hd__o21ai_1
X_19697_ _19914_/A _19911_/A vssd1 vssd1 vccd1 vccd1 _19771_/A sky130_fd_sc_hd__nand2_1
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18648_ _18638_/Y _18647_/X _18003_/X vssd1 vssd1 vccd1 vccd1 _18648_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18579_ _18554_/X _18576_/X _18580_/B vssd1 vssd1 vccd1 vccd1 _18579_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20610_ _20609_/X _25720_/Q _20614_/S vssd1 vssd1 vccd1 vccd1 _20611_/A sky130_fd_sc_hd__mux2_1
X_21590_ _21585_/X _21588_/X _21589_/X vssd1 vssd1 vccd1 vccd1 _21590_/X sky130_fd_sc_hd__a21o_1
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20541_ _23549_/A vssd1 vssd1 vccd1 vccd1 _23725_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23260_ _26573_/Q _23105_/X _23266_/S vssd1 vssd1 vccd1 vccd1 _23261_/A sky130_fd_sc_hd__mux2_1
X_20472_ _20471_/A _20471_/B _20471_/C vssd1 vssd1 vccd1 vccd1 _20472_/X sky130_fd_sc_hd__a21o_1
X_22211_ input4/X input270/X _22226_/S vssd1 vssd1 vccd1 vccd1 _22211_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23191_ _23191_/A vssd1 vssd1 vccd1 vccd1 _26542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22142_ _26166_/Q _22136_/X _22141_/X _22132_/X vssd1 vssd1 vccd1 vccd1 _26166_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput330 _16724_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[7] sky130_fd_sc_hd__buf_2
XFILLER_105_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput341 _16894_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[16] sky130_fd_sc_hd__buf_2
XFILLER_126_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput352 _16960_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[26] sky130_fd_sc_hd__buf_2
X_26950_ _26987_/CLK _26950_/D vssd1 vssd1 vccd1 vccd1 _26950_/Q sky130_fd_sc_hd__dfxtp_1
X_22073_ _26145_/Q _20926_/X _22077_/S vssd1 vssd1 vccd1 vccd1 _22074_/A sky130_fd_sc_hd__mux2_1
Xoutput363 _16835_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[7] sky130_fd_sc_hd__buf_2
Xoutput374 _16661_/X vssd1 vssd1 vccd1 vccd1 csb1[0] sky130_fd_sc_hd__buf_2
XFILLER_259_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput385 _17033_/X vssd1 vssd1 vccd1 vccd1 din0[18] sky130_fd_sc_hd__buf_2
XFILLER_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput396 _17046_/X vssd1 vssd1 vccd1 vccd1 din0[28] sky130_fd_sc_hd__buf_2
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21024_ _25882_/Q _20913_/X _21026_/S vssd1 vssd1 vccd1 vccd1 _21025_/A sky130_fd_sc_hd__mux2_1
X_25901_ _26282_/CLK _25901_/D vssd1 vssd1 vccd1 vccd1 _25901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26881_ _26881_/CLK _26881_/D vssd1 vssd1 vccd1 vccd1 _26881_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_87_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25832_ _27267_/CLK _25832_/D vssd1 vssd1 vccd1 vccd1 _25832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_263_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22975_ _23032_/S vssd1 vssd1 vccd1 vccd1 _22984_/S sky130_fd_sc_hd__clkbuf_2
X_25763_ _26593_/CLK _25763_/D vssd1 vssd1 vccd1 vccd1 _25763_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_256_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21926_ _21926_/A vssd1 vssd1 vccd1 vccd1 _26079_/D sky130_fd_sc_hd__clkbuf_1
X_24714_ hold3/A vssd1 vssd1 vccd1 vccd1 _24715_/B sky130_fd_sc_hd__inv_2
XFILLER_35_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25694_ _26240_/CLK _25694_/D vssd1 vssd1 vccd1 vccd1 _25694_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24645_ _24765_/A _24645_/B vssd1 vssd1 vccd1 vccd1 _24645_/Y sky130_fd_sc_hd__nand2_2
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21857_ _21857_/A vssd1 vssd1 vccd1 vccd1 _26056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20808_ _25800_/Q vssd1 vssd1 vccd1 vccd1 _20809_/A sky130_fd_sc_hd__clkbuf_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24576_ _24615_/A vssd1 vssd1 vccd1 vccd1 _24576_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21788_ _21788_/A vssd1 vssd1 vccd1 vccd1 _26026_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26315_ _26319_/CLK _26315_/D vssd1 vssd1 vccd1 vccd1 _26315_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_184_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23527_ _23610_/S vssd1 vssd1 vccd1 vccd1 _23540_/S sky130_fd_sc_hd__clkbuf_4
X_20739_ _20529_/X _25767_/Q _20739_/S vssd1 vssd1 vccd1 vccd1 _20740_/A sky130_fd_sc_hd__mux2_1
X_27295_ _27295_/CLK _27295_/D vssd1 vssd1 vccd1 vccd1 _27295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14260_ _15990_/S _14256_/X _14259_/X _13863_/A vssd1 vssd1 vccd1 vccd1 _14260_/X
+ sky130_fd_sc_hd__a211o_1
X_26246_ _26248_/CLK _26246_/D vssd1 vssd1 vccd1 vccd1 _26246_/Q sky130_fd_sc_hd__dfxtp_1
X_23458_ _26661_/Q _23066_/X _23458_/S vssd1 vssd1 vccd1 vccd1 _23459_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13211_ _18028_/A _12738_/X _13529_/A vssd1 vssd1 vccd1 vccd1 _13212_/A sky130_fd_sc_hd__o21ai_1
X_22409_ _22379_/X _22361_/B _22405_/X _22408_/Y _22402_/X vssd1 vssd1 vccd1 vccd1
+ _26239_/D sky130_fd_sc_hd__o221a_1
X_26177_ _26186_/CLK _26177_/D vssd1 vssd1 vccd1 vccd1 _26177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14191_ _18001_/A _17776_/A vssd1 vssd1 vccd1 vccd1 _14193_/B sky130_fd_sc_hd__nor2_2
X_23389_ _26630_/Q _23069_/X _23397_/S vssd1 vssd1 vccd1 vccd1 _23390_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13142_ _13142_/A vssd1 vssd1 vccd1 vccd1 _13159_/A sky130_fd_sc_hd__buf_2
X_25128_ _27189_/Q _25112_/X _25127_/X vssd1 vssd1 vccd1 vccd1 _27189_/D sky130_fd_sc_hd__o21ba_1
XFILLER_100_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13073_ _15561_/B vssd1 vssd1 vccd1 vccd1 _15255_/A sky130_fd_sc_hd__buf_4
X_17950_ _17819_/B _15342_/B _17950_/S vssd1 vssd1 vccd1 vccd1 _17950_/X sky130_fd_sc_hd__mux2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25059_ _25113_/A vssd1 vssd1 vccd1 vccd1 _25059_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16901_ _16901_/A _16952_/A vssd1 vssd1 vccd1 vccd1 _16957_/B sky130_fd_sc_hd__or2_1
XFILLER_239_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17881_ _17810_/B _17779_/Y _17909_/S vssd1 vssd1 vccd1 vccd1 _17881_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19620_ _27064_/Q _26061_/Q _19620_/C vssd1 vssd1 vccd1 vccd1 _19620_/X sky130_fd_sc_hd__and3_1
X_16832_ _16832_/A vssd1 vssd1 vccd1 vccd1 _16832_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19551_ _19551_/A vssd1 vssd1 vccd1 vccd1 _19551_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16763_ _22513_/A _16756_/X _16757_/X _19118_/B vssd1 vssd1 vccd1 vccd1 _16763_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_247_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13975_ _15516_/A _13969_/X _13974_/X _13311_/A vssd1 vssd1 vccd1 vccd1 _13975_/X
+ sky130_fd_sc_hd__o211a_1
X_18502_ _17259_/X _18439_/X _18441_/X _25540_/Q vssd1 vssd1 vccd1 vccd1 _18502_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_280_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15714_ _15714_/A vssd1 vssd1 vccd1 vccd1 _15988_/S sky130_fd_sc_hd__buf_4
XFILLER_46_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12926_ _15345_/A _14237_/D vssd1 vssd1 vccd1 vccd1 _12926_/X sky130_fd_sc_hd__or2_1
XFILLER_34_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19482_ _20487_/A _19482_/B vssd1 vssd1 vccd1 vccd1 _19551_/A sky130_fd_sc_hd__or2_4
XFILLER_234_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16694_ _16586_/B _17998_/A _14564_/X vssd1 vssd1 vccd1 vccd1 _16696_/A sky130_fd_sc_hd__a21o_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18433_ _19772_/A _18432_/C _25730_/Q vssd1 vssd1 vccd1 vccd1 _18434_/B sky130_fd_sc_hd__a21oi_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15645_ _15643_/X _15644_/X _15645_/S vssd1 vssd1 vccd1 vccd1 _15645_/X sky130_fd_sc_hd__mux2_1
X_12857_ _12850_/Y _15708_/A _13916_/A _15706_/A vssd1 vssd1 vccd1 vccd1 _12857_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18364_ _18364_/A vssd1 vssd1 vccd1 vccd1 _18364_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_199_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15576_ _15576_/A _15576_/B vssd1 vssd1 vccd1 vccd1 _15576_/X sky130_fd_sc_hd__or2_1
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _12808_/A vssd1 vssd1 vccd1 vccd1 _13269_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _17334_/A _17322_/C vssd1 vssd1 vccd1 vccd1 _17315_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14527_ _12674_/A _14362_/B _14525_/X _14526_/X vssd1 vssd1 vccd1 vccd1 _16581_/B
+ sky130_fd_sc_hd__a22o_1
X_18295_ _27105_/Q _19056_/A _18291_/X _18294_/X vssd1 vssd1 vccd1 vccd1 _18295_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_159_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17246_ _25501_/Q _25502_/Q _25503_/Q _25504_/Q vssd1 vssd1 vccd1 vccd1 _17253_/C
+ sky130_fd_sc_hd__and4_1
X_14458_ _14456_/X _14457_/X _14458_/S vssd1 vssd1 vccd1 vccd1 _14458_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13409_ _13409_/A vssd1 vssd1 vccd1 vccd1 _15826_/S sky130_fd_sc_hd__clkbuf_8
X_14389_ _26098_/Q _25999_/Q _14389_/S vssd1 vssd1 vccd1 vccd1 _14389_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17177_ _25485_/Q _17185_/B vssd1 vssd1 vccd1 vccd1 _17177_/X sky130_fd_sc_hd__or2_1
XFILLER_190_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16128_ _19034_/A _16621_/B _16614_/B _19048_/A _16127_/X vssd1 vssd1 vccd1 vccd1
+ _16612_/B sky130_fd_sc_hd__o41a_2
XFILLER_227_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16059_ _16057_/X _16058_/X _16059_/S vssd1 vssd1 vccd1 vccd1 _16059_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19818_ _19790_/A _27072_/Q _19817_/X vssd1 vssd1 vccd1 vccd1 _19819_/B sky130_fd_sc_hd__o21ai_1
XFILLER_69_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19749_ _27136_/Q _27070_/Q _19687_/B vssd1 vssd1 vccd1 vccd1 _19753_/A sky130_fd_sc_hd__a21oi_1
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22760_ _22760_/A vssd1 vssd1 vccd1 vccd1 _26365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_266_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21711_ _21654_/C _21654_/D _21715_/A _21349_/B vssd1 vssd1 vccd1 vccd1 _21713_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_253_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22691_ _23734_/A vssd1 vssd1 vccd1 vccd1 _22691_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24430_ _27016_/Q _24421_/X _24429_/Y _24415_/X vssd1 vssd1 vccd1 vccd1 _27016_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_240_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21642_ _21284_/A _19471_/X _21286_/A _25828_/Q _21346_/X vssd1 vssd1 vccd1 vccd1
+ _21642_/X sky130_fd_sc_hd__a221o_1
XFILLER_178_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24361_ _14237_/B _21884_/X _24361_/S vssd1 vssd1 vccd1 vccd1 _24781_/B sky130_fd_sc_hd__mux2_4
XFILLER_166_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21573_ _21573_/A vssd1 vssd1 vccd1 vccd1 _21573_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_178_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26100_ _27267_/CLK _26100_/D vssd1 vssd1 vccd1 vccd1 _26100_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23312_ _23312_/A vssd1 vssd1 vccd1 vccd1 _26596_/D sky130_fd_sc_hd__clkbuf_1
X_20524_ _23536_/A vssd1 vssd1 vccd1 vccd1 _23712_/A sky130_fd_sc_hd__buf_4
X_27080_ _27198_/CLK _27080_/D vssd1 vssd1 vccd1 vccd1 _27080_/Q sky130_fd_sc_hd__dfxtp_1
X_24292_ _26987_/Q _24293_/C _26988_/Q vssd1 vssd1 vccd1 vccd1 _24294_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26031_ _26240_/CLK _26031_/D vssd1 vssd1 vccd1 vccd1 _26031_/Q sky130_fd_sc_hd__dfxtp_1
X_23243_ _23243_/A vssd1 vssd1 vccd1 vccd1 _26565_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20455_ _27163_/Q _27097_/Q vssd1 vssd1 vccd1 vccd1 _20457_/A sky130_fd_sc_hd__nand2_1
XFILLER_193_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23174_ _23196_/A vssd1 vssd1 vccd1 vccd1 _23183_/S sky130_fd_sc_hd__buf_4
XFILLER_137_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20386_ _27128_/Q _20248_/X _20276_/X _20385_/Y vssd1 vssd1 vccd1 vccd1 _20386_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_284_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22125_ _26160_/Q _22122_/X _22124_/X input253/X _22118_/X vssd1 vssd1 vccd1 vccd1
+ _22125_/X sky130_fd_sc_hd__a221o_1
XFILLER_279_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22056_ _22056_/A vssd1 vssd1 vccd1 vccd1 _26137_/D sky130_fd_sc_hd__clkbuf_1
X_26933_ _27258_/CLK _26933_/D vssd1 vssd1 vccd1 vccd1 _26933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21007_ _25874_/Q _20887_/X _21015_/S vssd1 vssd1 vccd1 vccd1 _21008_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26864_ _27315_/CLK _26864_/D vssd1 vssd1 vccd1 vccd1 _26864_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25815_ _26881_/CLK _25815_/D vssd1 vssd1 vccd1 vccd1 _25815_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26795_ _27249_/CLK _26795_/D vssd1 vssd1 vccd1 vccd1 _26795_/Q sky130_fd_sc_hd__dfxtp_1
X_13760_ _26072_/Q _15484_/S _13759_/X _13762_/A vssd1 vssd1 vccd1 vccd1 _13760_/X
+ sky130_fd_sc_hd__o211a_1
X_22958_ _26454_/Q _22739_/X _22960_/S vssd1 vssd1 vccd1 vccd1 _22959_/A sky130_fd_sc_hd__mux2_1
X_25746_ _26282_/CLK _25746_/D vssd1 vssd1 vccd1 vccd1 _25746_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21909_ _20525_/X _26072_/Q _21911_/S vssd1 vssd1 vccd1 vccd1 _21910_/A sky130_fd_sc_hd__mux2_1
X_12711_ _14268_/S vssd1 vssd1 vccd1 vccd1 _15983_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_204_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13691_ _13691_/A vssd1 vssd1 vccd1 vccd1 _18593_/A sky130_fd_sc_hd__buf_4
XFILLER_231_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22889_ _22889_/A vssd1 vssd1 vccd1 vccd1 _26423_/D sky130_fd_sc_hd__clkbuf_1
X_25677_ _26278_/CLK _25677_/D vssd1 vssd1 vccd1 vccd1 _25677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15430_ _15430_/A _15430_/B vssd1 vssd1 vccd1 vccd1 _15430_/Y sky130_fd_sc_hd__nor2_1
X_24628_ _27067_/Q _24553_/B _24627_/Y _24619_/X vssd1 vssd1 vccd1 vccd1 _27067_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15361_ _16060_/S vssd1 vssd1 vccd1 vccd1 _15374_/S sky130_fd_sc_hd__buf_2
XFILLER_212_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24559_ _24559_/A _24569_/B vssd1 vssd1 vccd1 vccd1 _24559_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17100_ _20487_/B vssd1 vssd1 vccd1 vccd1 _25208_/B sky130_fd_sc_hd__inv_2
X_14312_ _13239_/A _14310_/X _14311_/X _13540_/A vssd1 vssd1 vccd1 vccd1 _14312_/X
+ sky130_fd_sc_hd__a211o_1
X_15292_ _15292_/A vssd1 vssd1 vccd1 vccd1 _15596_/S sky130_fd_sc_hd__clkbuf_4
X_18080_ _18861_/A _18080_/B vssd1 vssd1 vccd1 vccd1 _18080_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27278_ _27278_/CLK _27278_/D vssd1 vssd1 vccd1 vccd1 _27278_/Q sky130_fd_sc_hd__dfxtp_1
X_14243_ _25633_/Q _15532_/B _13578_/X _25601_/Q _14242_/X vssd1 vssd1 vccd1 vccd1
+ _23520_/A sky130_fd_sc_hd__a221o_4
XFILLER_8_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17031_ _17028_/X _16899_/B _17025_/X input223/X vssd1 vssd1 vccd1 vccd1 _17031_/X
+ sky130_fd_sc_hd__a22o_4
X_26229_ _26520_/CLK _26229_/D vssd1 vssd1 vccd1 vccd1 _26229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14174_ _25801_/Q _14103_/X _14107_/A _14173_/X vssd1 vssd1 vccd1 vccd1 _14174_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13125_ _13857_/A vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__buf_2
XFILLER_113_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18982_ _17967_/X _18056_/X _18191_/X _18321_/A vssd1 vssd1 vccd1 vccd1 _18982_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _14114_/S vssd1 vssd1 vccd1 vccd1 _15895_/S sky130_fd_sc_hd__clkbuf_8
X_17933_ _14022_/A _17784_/B _17933_/S vssd1 vssd1 vccd1 vccd1 _17933_/X sky130_fd_sc_hd__mux2_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17864_ _18362_/A vssd1 vssd1 vccd1 vccd1 _18859_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_159_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27132_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19603_ _19603_/A vssd1 vssd1 vccd1 vccd1 _19943_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16815_ _16815_/A vssd1 vssd1 vccd1 vccd1 _16815_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17795_ _17795_/A _16287_/B vssd1 vssd1 vccd1 vccd1 _17795_/X sky130_fd_sc_hd__or2b_1
XFILLER_54_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19534_ _25648_/Q _19536_/B vssd1 vssd1 vccd1 vccd1 _19534_/X sky130_fd_sc_hd__or2_1
X_16746_ _22500_/A _16742_/X _16743_/X _16636_/C vssd1 vssd1 vccd1 vccd1 _16746_/X
+ sky130_fd_sc_hd__a22o_1
X_13958_ _27301_/Q _26558_/Q _16005_/S vssd1 vssd1 vccd1 vccd1 _13958_/X sky130_fd_sc_hd__mux2_1
XFILLER_253_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12909_ _12946_/A _13916_/C _13916_/D vssd1 vssd1 vccd1 vccd1 _13397_/B sky130_fd_sc_hd__nand3_2
X_19465_ _27164_/Q _19465_/B vssd1 vssd1 vccd1 vccd1 _19465_/X sky130_fd_sc_hd__or2_1
XFILLER_35_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16677_ _17020_/A vssd1 vssd1 vccd1 vccd1 _17042_/A sky130_fd_sc_hd__clkbuf_2
X_13889_ _13889_/A vssd1 vssd1 vccd1 vccd1 _15982_/S sky130_fd_sc_hd__buf_2
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18416_ _18197_/X _18208_/X _18416_/S vssd1 vssd1 vccd1 vccd1 _18416_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15628_ _25813_/Q _16151_/S _15633_/S _15627_/X vssd1 vssd1 vccd1 vccd1 _15628_/X
+ sky130_fd_sc_hd__o211a_1
X_19396_ _19388_/X _19391_/X _19394_/X _19395_/X vssd1 vssd1 vccd1 vccd1 _19396_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18347_ _18064_/X _18050_/X _18347_/S vssd1 vssd1 vccd1 vccd1 _18347_/X sky130_fd_sc_hd__mux2_1
X_15559_ _15557_/X _15558_/X _15559_/S vssd1 vssd1 vccd1 vccd1 _15559_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18278_ _18792_/A _18253_/X _18269_/Y _18277_/X vssd1 vssd1 vccd1 vccd1 _18278_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17229_ _25027_/A vssd1 vssd1 vccd1 vccd1 _25466_/A sky130_fd_sc_hd__clkbuf_16
Xinput40 core_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput51 dout0[17] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_2
Xinput62 dout0[27] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_2
Xinput73 dout0[37] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_1
Xinput84 dout0[47] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__clkbuf_1
X_20240_ _27154_/Q _27088_/Q vssd1 vssd1 vccd1 vccd1 _20240_/Y sky130_fd_sc_hd__nand2_1
Xinput95 dout0[57] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20171_ _20119_/B _20169_/X _19698_/X _20675_/A vssd1 vssd1 vccd1 vccd1 _20173_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23930_ _23785_/X _26843_/Q _23930_/S vssd1 vssd1 vccd1 vccd1 _23931_/A sky130_fd_sc_hd__mux2_1
XFILLER_258_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23861_ _23917_/A vssd1 vssd1 vccd1 vccd1 _23930_/S sky130_fd_sc_hd__buf_6
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22812_ _22812_/A vssd1 vssd1 vccd1 vccd1 _26389_/D sky130_fd_sc_hd__clkbuf_1
X_25600_ _25607_/CLK _25600_/D vssd1 vssd1 vccd1 vccd1 _25600_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23792_ _23792_/A vssd1 vssd1 vccd1 vccd1 _26780_/D sky130_fd_sc_hd__clkbuf_1
X_26580_ _26580_/CLK _26580_/D vssd1 vssd1 vccd1 vccd1 _26580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25531_ _25553_/CLK _25531_/D vssd1 vssd1 vccd1 vccd1 _25531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22743_ _26359_/Q _22742_/X _22743_/S vssd1 vssd1 vccd1 vccd1 _22744_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25462_ _25462_/A vssd1 vssd1 vccd1 vccd1 _27325_/D sky130_fd_sc_hd__clkbuf_1
X_22674_ _22674_/A vssd1 vssd1 vccd1 vccd1 _26337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24413_ _24674_/B vssd1 vssd1 vccd1 vccd1 _24572_/A sky130_fd_sc_hd__clkinv_2
X_27201_ _27203_/CLK _27201_/D vssd1 vssd1 vccd1 vccd1 _27201_/Q sky130_fd_sc_hd__dfxtp_1
X_21625_ input64/X input100/X _21646_/S vssd1 vssd1 vccd1 vccd1 _21626_/A sky130_fd_sc_hd__mux2_8
XFILLER_178_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25393_ _25393_/A _25393_/B vssd1 vssd1 vccd1 vccd1 _25450_/A sky130_fd_sc_hd__or2_4
XFILLER_240_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24344_ _24350_/S _25493_/Q _25492_/Q _17691_/X vssd1 vssd1 vccd1 vccd1 _24347_/B
+ sky130_fd_sc_hd__o31a_1
X_27132_ _27132_/CLK _27132_/D vssd1 vssd1 vccd1 vccd1 _27132_/Q sky130_fd_sc_hd__dfxtp_4
X_21556_ _21556_/A vssd1 vssd1 vccd1 vccd1 _21556_/X sky130_fd_sc_hd__buf_4
XFILLER_32_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20507_ _23523_/A vssd1 vssd1 vccd1 vccd1 _23699_/A sky130_fd_sc_hd__clkbuf_4
X_27063_ _27160_/CLK _27063_/D vssd1 vssd1 vccd1 vccd1 _27063_/Q sky130_fd_sc_hd__dfxtp_1
X_24275_ _26982_/Q _26981_/Q _24275_/C vssd1 vssd1 vccd1 vccd1 _24278_/B sky130_fd_sc_hd__and3_1
XFILLER_181_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21487_ _21480_/X _21486_/X _21473_/X vssd1 vssd1 vccd1 vccd1 _21487_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_154_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26014_ _27280_/CLK _26014_/D vssd1 vssd1 vccd1 vccd1 _26014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23226_ _23226_/A vssd1 vssd1 vccd1 vccd1 _26557_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20438_ _20436_/Y _20437_/X _20434_/A _19820_/S vssd1 vssd1 vccd1 vccd1 _20438_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_181_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23157_ _26527_/Q _23060_/X _23161_/S vssd1 vssd1 vccd1 vccd1 _23158_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20369_ _20367_/Y _20369_/B vssd1 vssd1 vccd1 vccd1 _20370_/B sky130_fd_sc_hd__and2b_1
XFILLER_107_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22108_ _22121_/A _22239_/B vssd1 vssd1 vccd1 vccd1 _22200_/A sky130_fd_sc_hd__nor2_1
XFILLER_267_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23088_ _23088_/A vssd1 vssd1 vccd1 vccd1 _26503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22039_ _22039_/A vssd1 vssd1 vccd1 vccd1 _26129_/D sky130_fd_sc_hd__clkbuf_1
X_26916_ _26916_/CLK _26916_/D vssd1 vssd1 vccd1 vccd1 _26916_/Q sky130_fd_sc_hd__dfxtp_1
X_14930_ _14724_/X _14839_/Y _14929_/X _14827_/X vssd1 vssd1 vccd1 vccd1 _19408_/A
+ sky130_fd_sc_hd__a211o_4
XTAP_5644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26847_ _27269_/CLK _26847_/D vssd1 vssd1 vccd1 vccd1 _26847_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14861_ _26093_/Q _14846_/B _14859_/X _14860_/X vssd1 vssd1 vccd1 vccd1 _14861_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ _16833_/A _19639_/B vssd1 vssd1 vccd1 vccd1 _16639_/B sky130_fd_sc_hd__and2_2
X_13812_ _13806_/X _13807_/X _13811_/X _13339_/A vssd1 vssd1 vccd1 vccd1 _13818_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17580_ _17595_/A _17580_/B vssd1 vssd1 vccd1 vccd1 _25576_/D sky130_fd_sc_hd__nor2_1
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14792_ _14792_/A vssd1 vssd1 vccd1 vccd1 _14793_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_90_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26778_ _27326_/CLK _26778_/D vssd1 vssd1 vccd1 vccd1 _26778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16531_ _26939_/Q _26423_/Q _16533_/A vssd1 vssd1 vccd1 vccd1 _16531_/X sky130_fd_sc_hd__mux2_1
X_13743_ _25918_/Q _13737_/A _13742_/Y _13748_/A vssd1 vssd1 vccd1 vccd1 _13744_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_25729_ _26271_/CLK _25729_/D vssd1 vssd1 vccd1 vccd1 _25729_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_250_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19250_ _19087_/X _19244_/X _19249_/X _18891_/X vssd1 vssd1 vccd1 vccd1 _19251_/B
+ sky130_fd_sc_hd__a22o_1
X_16462_ _16462_/A _16462_/B vssd1 vssd1 vccd1 vccd1 _25161_/A sky130_fd_sc_hd__xor2_4
X_13674_ _13791_/A _13672_/X _13673_/X _12754_/A vssd1 vssd1 vccd1 vccd1 _13674_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18201_ _17951_/X _17935_/X _18265_/S vssd1 vssd1 vccd1 vccd1 _18201_/X sky130_fd_sc_hd__mux2_1
X_15413_ _15405_/X _15412_/X _14818_/A vssd1 vssd1 vccd1 vccd1 _15413_/Y sky130_fd_sc_hd__o21ai_1
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19181_ _19087_/X _19177_/X _20251_/A _18884_/X vssd1 vssd1 vccd1 vccd1 _19182_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16393_ _15167_/X _26903_/Q _26775_/Q _15030_/S _15169_/X vssd1 vssd1 vccd1 vccd1
+ _16393_/X sky130_fd_sc_hd__a221o_1
XPHY_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18132_ _25502_/Q _18559_/A _18123_/X _18130_/X _18574_/A vssd1 vssd1 vccd1 vccd1
+ _18132_/X sky130_fd_sc_hd__o221a_1
XFILLER_157_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15344_ _15344_/A vssd1 vssd1 vccd1 vccd1 _19156_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18063_ _17957_/X _17953_/X _18063_/S vssd1 vssd1 vccd1 vccd1 _18063_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15275_ _26542_/Q _26150_/Q _15276_/S vssd1 vssd1 vccd1 vccd1 _15275_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17014_ _16810_/A _17008_/X _16883_/B _17013_/X input244/X vssd1 vssd1 vccd1 vccd1
+ _17014_/X sky130_fd_sc_hd__a32o_4
X_14226_ _13475_/A _14224_/X _14225_/X _15939_/A vssd1 vssd1 vccd1 vccd1 _14226_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_256_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14157_ _13614_/A _14150_/X _14156_/Y _12700_/A vssd1 vssd1 vccd1 vccd1 _14157_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13108_ _14713_/C vssd1 vssd1 vccd1 vccd1 _13717_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_258_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14088_ _14086_/X _14087_/X _14115_/S vssd1 vssd1 vccd1 vccd1 _14088_/X sky130_fd_sc_hd__mux2_1
X_18965_ _19037_/C _18965_/B vssd1 vssd1 vccd1 vccd1 _18965_/X sky130_fd_sc_hd__or2_2
XFILLER_26_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13039_ _14351_/S vssd1 vssd1 vccd1 vccd1 _14513_/S sky130_fd_sc_hd__clkbuf_2
X_17916_ _17983_/A vssd1 vssd1 vccd1 vccd1 _18349_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18896_ _18896_/A _18896_/B vssd1 vssd1 vccd1 vccd1 _18896_/X sky130_fd_sc_hd__or2_1
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17847_ _19237_/B _19237_/C _17846_/X vssd1 vssd1 vccd1 vccd1 _19355_/C sky130_fd_sc_hd__a21o_1
XFILLER_226_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17778_ _17671_/X _17768_/X _17775_/Y _16853_/A _19219_/A vssd1 vssd1 vccd1 vccd1
+ _18005_/C sky130_fd_sc_hd__a32o_1
XFILLER_214_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19517_ _25641_/Q _19523_/B vssd1 vssd1 vccd1 vccd1 _19517_/X sky130_fd_sc_hd__or2_1
XFILLER_240_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16729_ _18539_/A _16729_/B vssd1 vssd1 vccd1 vccd1 _18541_/A sky130_fd_sc_hd__xnor2_4
XFILLER_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_530 _17048_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_541 _25743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19448_ _19448_/A _19448_/B vssd1 vssd1 vccd1 vccd1 _19448_/Y sky130_fd_sc_hd__nand2_1
XINSDIODE2_552 _16992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19379_ _25752_/Q vssd1 vssd1 vccd1 vccd1 _19381_/A sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_56_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26599_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_188_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21410_ _21410_/A vssd1 vssd1 vccd1 vccd1 _21410_/Y sky130_fd_sc_hd__inv_2
X_22390_ _22390_/A _22390_/B vssd1 vssd1 vccd1 vccd1 _22390_/Y sky130_fd_sc_hd__nor2_1
XFILLER_163_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21341_ _25943_/Q _21310_/X _21340_/Y _21330_/X vssd1 vssd1 vccd1 vccd1 _25943_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_135_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24060_ _24060_/A vssd1 vssd1 vccd1 vccd1 _26900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_265_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21272_ _21407_/A _21269_/X _21271_/Y _21259_/X vssd1 vssd1 vccd1 vccd1 _21273_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_144_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23011_ _26477_/Q _22711_/X _23017_/S vssd1 vssd1 vccd1 vccd1 _23012_/A sky130_fd_sc_hd__mux2_1
X_20223_ _22638_/B vssd1 vssd1 vccd1 vccd1 _20223_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_265_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20154_ _20154_/A _20154_/B vssd1 vssd1 vccd1 vccd1 _20154_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24962_ _24605_/A _24941_/X _24938_/X vssd1 vssd1 vccd1 vccd1 _24962_/Y sky130_fd_sc_hd__a21oi_1
X_20085_ _20061_/X _20083_/X _20084_/Y vssd1 vssd1 vccd1 vccd1 _20085_/X sky130_fd_sc_hd__a21bo_1
XFILLER_246_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26701_ _26925_/CLK _26701_/D vssd1 vssd1 vccd1 vccd1 _26701_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23913_ _23760_/X _26835_/Q _23915_/S vssd1 vssd1 vccd1 vccd1 _23914_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24893_ _27131_/Q _24896_/B vssd1 vssd1 vccd1 vccd1 _24893_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26632_ _26920_/CLK _26632_/D vssd1 vssd1 vccd1 vccd1 _26632_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_261_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23844_ _23844_/A vssd1 vssd1 vccd1 vccd1 _26804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26563_ _27330_/A _26563_/D vssd1 vssd1 vccd1 vccd1 _26563_/Q sky130_fd_sc_hd__dfxtp_1
X_23775_ _23775_/A vssd1 vssd1 vccd1 vccd1 _26775_/D sky130_fd_sc_hd__clkbuf_1
X_20987_ _20987_/A vssd1 vssd1 vccd1 vccd1 _25865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_26_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25514_ _25518_/CLK _25514_/D vssd1 vssd1 vccd1 vccd1 _25514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22726_ _22726_/A vssd1 vssd1 vccd1 vccd1 _26353_/D sky130_fd_sc_hd__clkbuf_1
X_26494_ _27272_/CLK _26494_/D vssd1 vssd1 vccd1 vccd1 _26494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22657_ _26332_/Q _22656_/X _22657_/S vssd1 vssd1 vccd1 vccd1 _22658_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25445_ _25445_/A vssd1 vssd1 vccd1 vccd1 _27317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21608_ _21604_/Y _21607_/X _21556_/X vssd1 vssd1 vccd1 vccd1 _21608_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13390_ _25920_/Q _13737_/A _13389_/Y _25795_/Q vssd1 vssd1 vccd1 vccd1 _13391_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_22588_ _22580_/X _22586_/Y _22587_/X vssd1 vssd1 vccd1 vccd1 _26310_/D sky130_fd_sc_hd__a21oi_1
XFILLER_223_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25376_ _27287_/Q _23763_/A _25376_/S vssd1 vssd1 vccd1 vccd1 _25377_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27115_ _27117_/CLK _27115_/D vssd1 vssd1 vccd1 vccd1 _27115_/Q sky130_fd_sc_hd__dfxtp_4
X_24327_ _24327_/A _24327_/B _24331_/C vssd1 vssd1 vccd1 vccd1 _27000_/D sky130_fd_sc_hd__nor3_1
X_21539_ input57/X input92/X _21553_/S vssd1 vssd1 vccd1 vccd1 _21540_/A sky130_fd_sc_hd__mux2_8
XFILLER_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15060_ _15057_/X _15059_/X _15060_/S vssd1 vssd1 vccd1 vccd1 _15060_/X sky130_fd_sc_hd__mux2_1
X_24258_ _26976_/Q _26975_/Q _24258_/C vssd1 vssd1 vccd1 vccd1 _24260_/B sky130_fd_sc_hd__and3_1
X_27046_ _27049_/CLK _27046_/D vssd1 vssd1 vccd1 vccd1 _27046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14011_ _27269_/Q _26462_/Q _14252_/S vssd1 vssd1 vccd1 vccd1 _14011_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23209_ _26551_/Q _23136_/X _23209_/S vssd1 vssd1 vccd1 vccd1 _23210_/A sky130_fd_sc_hd__mux2_1
X_24189_ _26953_/Q _24191_/C _24188_/Y vssd1 vssd1 vccd1 vccd1 _26953_/D sky130_fd_sc_hd__o21a_1
XFILLER_175_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18750_ _27211_/Q _19462_/B vssd1 vssd1 vccd1 vccd1 _18750_/X sky130_fd_sc_hd__and2_1
XTAP_5430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15962_ _13585_/X _26404_/Q _15826_/S _15961_/X vssd1 vssd1 vccd1 vccd1 _15962_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput230 localMemory_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 input230/X sky130_fd_sc_hd__buf_6
XTAP_5452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput241 localMemory_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input241/X sky130_fd_sc_hd__buf_6
X_17701_ _17706_/A _17701_/B vssd1 vssd1 vccd1 vccd1 _17701_/X sky130_fd_sc_hd__and2_1
XTAP_5463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput252 localMemory_wb_we_i vssd1 vssd1 vccd1 vccd1 _21715_/A sky130_fd_sc_hd__clkbuf_1
X_14913_ _27324_/Q _26581_/Q _14996_/S vssd1 vssd1 vccd1 vccd1 _14913_/X sky130_fd_sc_hd__mux2_1
Xinput263 manufacturerID[9] vssd1 vssd1 vccd1 vccd1 input263/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18681_ _18681_/A vssd1 vssd1 vccd1 vccd1 _18682_/A sky130_fd_sc_hd__clkbuf_2
Xinput274 partID[4] vssd1 vssd1 vccd1 vccd1 input274/X sky130_fd_sc_hd__clkbuf_1
XTAP_5485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15893_ _15720_/S _15887_/X _15889_/X _15892_/X _13630_/X vssd1 vssd1 vccd1 vccd1
+ _15893_/X sky130_fd_sc_hd__a311o_1
XTAP_5496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ _19774_/A _17584_/X _17604_/X _17631_/X vssd1 vssd1 vccd1 vccd1 _17633_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_63_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14844_ _14878_/S vssd1 vssd1 vccd1 vccd1 _14960_/B sky130_fd_sc_hd__buf_2
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17563_ _17575_/A _17563_/B vssd1 vssd1 vccd1 vccd1 _25572_/D sky130_fd_sc_hd__nor2_1
XFILLER_251_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14775_ _16517_/A _14767_/X _14774_/X _12758_/A vssd1 vssd1 vccd1 vccd1 _14776_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19302_ _27159_/Q _19302_/B vssd1 vssd1 vccd1 vccd1 _19302_/X sky130_fd_sc_hd__or2_1
XFILLER_232_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16514_ _16533_/A vssd1 vssd1 vccd1 vccd1 _16526_/S sky130_fd_sc_hd__buf_2
X_13726_ _15633_/S _13724_/X _13725_/X _14647_/A vssd1 vssd1 vccd1 vccd1 _13726_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17494_ _26063_/Q vssd1 vssd1 vccd1 vccd1 _17706_/A sky130_fd_sc_hd__inv_2
XFILLER_31_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19233_ _18383_/A _19231_/Y _18705_/A vssd1 vssd1 vccd1 vccd1 _19234_/C sky130_fd_sc_hd__o21ba_1
X_16445_ _16336_/X _16443_/X _16444_/X _12756_/A vssd1 vssd1 vccd1 vccd1 _16445_/X
+ sky130_fd_sc_hd__o211a_1
X_13657_ _13657_/A vssd1 vssd1 vccd1 vccd1 _16021_/S sky130_fd_sc_hd__buf_4
XFILLER_189_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19164_ _27091_/Q _18815_/X _18816_/X _27189_/Q _18817_/X vssd1 vssd1 vccd1 vccd1
+ _19164_/X sky130_fd_sc_hd__a221o_1
XFILLER_192_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _25824_/Q _27258_/Q _16377_/S vssd1 vssd1 vccd1 vccd1 _16376_/X sky130_fd_sc_hd__mux2_1
X_13588_ _13402_/A _13581_/X _13587_/X _13433_/X vssd1 vssd1 vccd1 vccd1 _13588_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_185_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18115_ _27200_/Q _19331_/B _18110_/X _18114_/X vssd1 vssd1 vccd1 vccd1 _18115_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_9_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15327_ _26086_/Q _25891_/Q _16256_/B vssd1 vssd1 vccd1 vccd1 _15327_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19095_ _27057_/Q _18503_/A _19092_/X _19094_/X _18519_/A vssd1 vssd1 vccd1 vccd1
+ _19095_/X sky130_fd_sc_hd__o221a_2
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18046_ _18043_/X _18045_/X _18210_/S vssd1 vssd1 vccd1 vccd1 _18046_/X sky130_fd_sc_hd__mux2_1
X_15258_ _27253_/Q _16388_/B vssd1 vssd1 vccd1 vccd1 _15258_/X sky130_fd_sc_hd__or2_1
XFILLER_172_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14209_ _15588_/A _26100_/Q _26001_/Q _13675_/S _12738_/C vssd1 vssd1 vccd1 vccd1
+ _14209_/X sky130_fd_sc_hd__a221o_1
XFILLER_160_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15189_ _12704_/A _15177_/X _15188_/X _14710_/A vssd1 vssd1 vccd1 vccd1 _15189_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_99_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_174_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25725_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_235_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19997_ _27144_/Q _19957_/B _19996_/X vssd1 vssd1 vccd1 vccd1 _19999_/C sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_103_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26319_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_259_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18948_ _17287_/X _18556_/A _18557_/A _25549_/Q vssd1 vssd1 vccd1 vccd1 _18948_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18879_ _18741_/X _18876_/X _18878_/Y vssd1 vssd1 vccd1 vccd1 _18879_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_239_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20910_ _23725_/A vssd1 vssd1 vccd1 vccd1 _20910_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21890_ _21946_/A vssd1 vssd1 vccd1 vccd1 _21959_/S sky130_fd_sc_hd__buf_6
XFILLER_66_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20841_ _20841_/A vssd1 vssd1 vccd1 vccd1 _25816_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_270_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23560_ _26699_/Q _23558_/X _23572_/S vssd1 vssd1 vccd1 vccd1 _23561_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20772_ _20592_/X _25782_/Q _20772_/S vssd1 vssd1 vccd1 vccd1 _20773_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_360 input217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22511_ _22511_/A _22513_/B vssd1 vssd1 vccd1 vccd1 _22512_/A sky130_fd_sc_hd__and2_1
XINSDIODE2_371 _17064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_382 _16718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23491_ _26676_/Q _23114_/X _23491_/S vssd1 vssd1 vccd1 vccd1 _23492_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_393 _17034_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22442_ _24415_/A vssd1 vssd1 vccd1 vccd1 _22442_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_211_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25230_ _27221_/Q _25225_/X _25228_/X _24736_/B _25229_/X vssd1 vssd1 vccd1 vccd1
+ _27221_/D sky130_fd_sc_hd__o221a_1
XFILLER_136_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25161_ _25161_/A vssd1 vssd1 vccd1 vccd1 _25161_/Y sky130_fd_sc_hd__inv_2
X_22373_ _26235_/Q _26228_/Q _22376_/S vssd1 vssd1 vccd1 vccd1 _22374_/B sky130_fd_sc_hd__mux2_1
XFILLER_164_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24112_ _26923_/Q _23558_/X _24120_/S vssd1 vssd1 vccd1 vccd1 _24113_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21324_ _21320_/X _21323_/X _21290_/X vssd1 vssd1 vccd1 vccd1 _21324_/X sky130_fd_sc_hd__a21o_1
XFILLER_191_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25092_ _25119_/A vssd1 vssd1 vccd1 vccd1 _25092_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24043_ _24043_/A vssd1 vssd1 vccd1 vccd1 _26892_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21255_ _20626_/A _21545_/A _21279_/A _21254_/X vssd1 vssd1 vccd1 vccd1 _21255_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20206_ _20206_/A _20206_/B _20206_/C vssd1 vssd1 vccd1 vccd1 _20206_/X sky130_fd_sc_hd__or3_1
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21186_ _21186_/A vssd1 vssd1 vccd1 vccd1 _25932_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20137_ _27150_/Q _20135_/Y _20371_/S vssd1 vssd1 vccd1 vccd1 _20137_/X sky130_fd_sc_hd__mux2_2
X_25994_ _27156_/CLK _25994_/D vssd1 vssd1 vccd1 vccd1 _25994_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24945_ _27147_/Q _24930_/X _24944_/Y _24921_/X vssd1 vssd1 vccd1 vccd1 _27147_/D
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_20 _19043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20068_ _27116_/Q _19877_/X _19967_/X _20067_/X vssd1 vssd1 vccd1 vccd1 _20068_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_218_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_31 _19308_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_42 _20644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_53 _20643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_64 _20652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _15706_/C vssd1 vssd1 vccd1 vccd1 _14834_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24876_ _24873_/Y _24875_/X _24871_/X vssd1 vssd1 vccd1 vccd1 _27125_/D sky130_fd_sc_hd__a21oi_1
XINSDIODE2_75 _20694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_86 _21878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_97 _21441_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26615_ _27257_/CLK _26615_/D vssd1 vssd1 vccd1 vccd1 _26615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23827_ _23827_/A vssd1 vssd1 vccd1 vccd1 _26796_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26546_ _27292_/CLK _26546_/D vssd1 vssd1 vccd1 vccd1 _26546_/Q sky130_fd_sc_hd__dfxtp_1
X_14560_ _25724_/Q _14559_/X _14560_/S vssd1 vssd1 vccd1 vccd1 _17807_/A sky130_fd_sc_hd__mux2_2
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23758_ _23757_/X _26770_/Q _23764_/S vssd1 vssd1 vccd1 vccd1 _23759_/A sky130_fd_sc_hd__mux2_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _26918_/Q _26402_/Q _13535_/S vssd1 vssd1 vccd1 vccd1 _13511_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22709_ _26348_/Q _22707_/X _22721_/S vssd1 vssd1 vccd1 vccd1 _22710_/A sky130_fd_sc_hd__mux2_1
X_14491_ _13744_/X _14485_/Y _14237_/A vssd1 vssd1 vccd1 vccd1 _14491_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26477_ _26609_/CLK _26477_/D vssd1 vssd1 vccd1 vccd1 _26477_/Q sky130_fd_sc_hd__dfxtp_1
X_23689_ _23689_/A vssd1 vssd1 vccd1 vccd1 _26748_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _12705_/A _16221_/X _16229_/X _14710_/A vssd1 vssd1 vccd1 vccd1 _16230_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_70_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13442_ _12770_/A _26886_/Q _26758_/Q _15796_/S _13050_/A vssd1 vssd1 vccd1 vccd1
+ _13442_/X sky130_fd_sc_hd__a221o_1
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25428_ _25450_/A vssd1 vssd1 vccd1 vccd1 _25437_/S sky130_fd_sc_hd__buf_4
XFILLER_16_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16161_ _26117_/Q _26018_/Q _16161_/S vssd1 vssd1 vccd1 vccd1 _16161_/X sky130_fd_sc_hd__mux2_1
X_13373_ _17971_/B _18006_/C vssd1 vssd1 vccd1 vccd1 _14481_/B sky130_fd_sc_hd__or2_2
XFILLER_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25359_ _27279_/Q _23738_/A _25365_/S vssd1 vssd1 vccd1 vccd1 _25360_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15112_ _15111_/X _26710_/Q _26838_/Q _15121_/S _14771_/A vssd1 vssd1 vccd1 vccd1
+ _15112_/X sky130_fd_sc_hd__a221o_1
XFILLER_10_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27317_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16092_ _16348_/S _16090_/X _16091_/X _13274_/X vssd1 vssd1 vccd1 vccd1 _16093_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27029_ _27058_/CLK _27029_/D vssd1 vssd1 vccd1 vccd1 _27029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19920_ _19920_/A vssd1 vssd1 vccd1 vccd1 _20119_/B sky130_fd_sc_hd__buf_2
X_15043_ _14623_/A _15021_/X _15028_/X _15042_/X _14683_/A vssd1 vssd1 vccd1 vccd1
+ _15043_/X sky130_fd_sc_hd__a311o_1
XFILLER_253_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19851_ _20643_/A _19708_/A _19850_/X _19604_/X vssd1 vssd1 vccd1 vccd1 _19976_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_122_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18802_ _18548_/A _18801_/X _17829_/A _16038_/B vssd1 vssd1 vccd1 vccd1 _18803_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19782_ _19834_/C _19764_/Y _19765_/X _19781_/X vssd1 vssd1 vccd1 vccd1 _19782_/Y
+ sky130_fd_sc_hd__o211ai_1
X_16994_ _22480_/A _16988_/X _16990_/X _18357_/A vssd1 vssd1 vccd1 vccd1 _16994_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18733_ _18861_/A vssd1 vssd1 vccd1 vccd1 _18733_/X sky130_fd_sc_hd__buf_2
XFILLER_283_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15945_ _15933_/X _15936_/X _15944_/X vssd1 vssd1 vccd1 vccd1 _15945_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_37_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18664_ _19912_/A _19268_/B vssd1 vssd1 vccd1 vccd1 _18666_/B sky130_fd_sc_hd__nor2_1
XFILLER_236_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15876_ _25643_/Q _13803_/B _14611_/A vssd1 vssd1 vccd1 vccd1 _15876_/X sky130_fd_sc_hd__a21o_1
XFILLER_252_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ _17615_/A _17615_/B vssd1 vssd1 vccd1 vccd1 _25585_/D sky130_fd_sc_hd__nor2_1
XFILLER_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14827_ _14827_/A vssd1 vssd1 vccd1 vccd1 _14827_/X sky130_fd_sc_hd__buf_2
X_18595_ _18942_/B _19573_/B _18636_/A vssd1 vssd1 vccd1 vccd1 _18595_/X sky130_fd_sc_hd__o21a_1
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17546_ _25907_/Q _17544_/X _17545_/X vssd1 vssd1 vccd1 vccd1 _17546_/Y sky130_fd_sc_hd__o21ai_2
X_14758_ _14758_/A vssd1 vssd1 vccd1 vccd1 _14759_/A sky130_fd_sc_hd__buf_2
XFILLER_44_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13709_ _26628_/Q _26724_/Q _15548_/S vssd1 vssd1 vccd1 vccd1 _13709_/X sky130_fd_sc_hd__mux2_1
X_17477_ _16679_/B _17476_/Y _21868_/A vssd1 vssd1 vccd1 vccd1 _17482_/A sky130_fd_sc_hd__a21oi_1
X_14689_ _12777_/A _26906_/Q _26778_/Q _16467_/A _16484_/A vssd1 vssd1 vccd1 vccd1
+ _14689_/X sky130_fd_sc_hd__a221o_1
XFILLER_149_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19216_ _17738_/B _18972_/X _18973_/X _19215_/Y vssd1 vssd1 vccd1 vccd1 _19216_/X
+ sky130_fd_sc_hd__a211o_1
X_16428_ _25824_/Q _27258_/Q _16428_/S vssd1 vssd1 vccd1 vccd1 _16428_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19147_ _25744_/Q _19146_/C _25745_/Q vssd1 vssd1 vccd1 vccd1 _19148_/B sky130_fd_sc_hd__a21oi_1
X_16359_ _27288_/Q _26481_/Q _16359_/S vssd1 vssd1 vccd1 vccd1 _16359_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19078_ _19078_/A vssd1 vssd1 vccd1 vccd1 _19078_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18029_ _25725_/Q _19879_/A vssd1 vssd1 vccd1 vccd1 _18227_/C sky130_fd_sc_hd__or2_2
XFILLER_278_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21040_ _25889_/Q _20935_/X _21048_/S vssd1 vssd1 vccd1 vccd1 _21041_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22991_ _26468_/Q _22682_/X _22995_/S vssd1 vssd1 vccd1 vccd1 _22992_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24730_ _27089_/Q _24724_/X _24729_/Y _24720_/X vssd1 vssd1 vccd1 vccd1 _24731_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_21942_ _20588_/X _26087_/Q _21944_/S vssd1 vssd1 vccd1 vccd1 _21943_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21873_ _21873_/A vssd1 vssd1 vccd1 vccd1 _21874_/A sky130_fd_sc_hd__buf_2
X_24661_ _27073_/Q _24657_/X _24659_/Y _24660_/X vssd1 vssd1 vccd1 vccd1 _24662_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_leaf_71_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26462_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26400_ _26433_/CLK _26400_/D vssd1 vssd1 vccd1 vccd1 _26400_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_231_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20824_ _25808_/Q vssd1 vssd1 vccd1 vccd1 _20825_/A sky130_fd_sc_hd__clkbuf_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23612_ _25249_/C _23860_/B vssd1 vssd1 vccd1 vccd1 _23669_/A sky130_fd_sc_hd__nor2_2
X_24592_ _24948_/A _24595_/B vssd1 vssd1 vccd1 vccd1 _24592_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26331_ _26462_/CLK _26331_/D vssd1 vssd1 vccd1 vccd1 _26331_/Q sky130_fd_sc_hd__dfxtp_2
X_23543_ _23610_/S vssd1 vssd1 vccd1 vccd1 _23556_/S sky130_fd_sc_hd__buf_6
X_20755_ _20559_/X _25774_/Q _20761_/S vssd1 vssd1 vccd1 vccd1 _20756_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_190 _16827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26262_ _27110_/CLK _26262_/D vssd1 vssd1 vccd1 vccd1 _26262_/Q sky130_fd_sc_hd__dfxtp_1
X_23474_ _26668_/Q _23089_/X _23480_/S vssd1 vssd1 vccd1 vccd1 _23475_/A sky130_fd_sc_hd__mux2_1
X_20686_ _20686_/A vssd1 vssd1 vccd1 vccd1 _20686_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22425_ _26243_/Q _22430_/B vssd1 vssd1 vccd1 vccd1 _22425_/X sky130_fd_sc_hd__or2_1
XFILLER_195_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25213_ _27216_/Q _25204_/X _25207_/X _24715_/B _25212_/X vssd1 vssd1 vccd1 vccd1
+ _27216_/D sky130_fd_sc_hd__o221a_1
XFILLER_210_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26193_ _26297_/CLK _26193_/D vssd1 vssd1 vccd1 vccd1 _26193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22356_ _22356_/A _22533_/B vssd1 vssd1 vccd1 vccd1 _22357_/A sky130_fd_sc_hd__and2_1
XFILLER_136_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25144_ _27192_/Q _25137_/X _25141_/X _25143_/Y _22402_/X vssd1 vssd1 vccd1 vccd1
+ _27192_/D sky130_fd_sc_hd__o221a_1
XFILLER_237_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21307_ _21304_/Y _21306_/Y _21297_/X vssd1 vssd1 vccd1 vccd1 _21307_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_152_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25075_ _22498_/A _25065_/X _25060_/X _16635_/C _25052_/X vssd1 vssd1 vccd1 vccd1
+ _25075_/X sky130_fd_sc_hd__a221o_1
X_22287_ _26207_/Q _22279_/X _22285_/X _26308_/Q _22286_/X vssd1 vssd1 vccd1 vccd1
+ _22287_/X sky130_fd_sc_hd__a221o_1
XFILLER_105_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24026_ _26885_/Q _23539_/X _24026_/S vssd1 vssd1 vccd1 vccd1 _24027_/A sky130_fd_sc_hd__mux2_1
X_21238_ _21231_/X _21234_/X _21237_/X vssd1 vssd1 vccd1 vccd1 _21238_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_105_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21169_ _21172_/A _21169_/B vssd1 vssd1 vccd1 vccd1 _21170_/A sky130_fd_sc_hd__or2_1
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25977_ _27022_/CLK _25977_/D vssd1 vssd1 vccd1 vccd1 _25977_/Q sky130_fd_sc_hd__dfxtp_4
X_13991_ _13084_/A _26690_/Q _26818_/Q _15890_/S _13611_/A vssd1 vssd1 vccd1 vccd1
+ _13991_/X sky130_fd_sc_hd__a221o_1
XFILLER_19_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15730_ _27310_/Q _26567_/Q _15734_/S vssd1 vssd1 vccd1 vccd1 _15730_/X sky130_fd_sc_hd__mux2_1
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _12942_/A vssd1 vssd1 vccd1 vccd1 _14325_/S sky130_fd_sc_hd__clkbuf_2
X_24928_ _24572_/A _24917_/X _24909_/X vssd1 vssd1 vccd1 vccd1 _24928_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _26668_/Q _25708_/Q _16086_/S vssd1 vssd1 vccd1 vccd1 _15661_/X sky130_fd_sc_hd__mux2_1
XFILLER_234_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12873_ _12873_/A vssd1 vssd1 vccd1 vccd1 _14486_/A sky130_fd_sc_hd__clkbuf_2
X_24859_ _24877_/A vssd1 vssd1 vccd1 vccd1 _24873_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17400_ _17428_/A _17400_/B _17401_/B vssd1 vssd1 vccd1 vccd1 _25551_/D sky130_fd_sc_hd__nor3_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14612_ _14612_/A vssd1 vssd1 vccd1 vccd1 _15135_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ _19772_/A _18432_/C vssd1 vssd1 vccd1 vccd1 _19768_/B sky130_fd_sc_hd__or2_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _15676_/A _27280_/Q _26473_/Q _16178_/S _15576_/A vssd1 vssd1 vccd1 vccd1
+ _15592_/X sky130_fd_sc_hd__a221o_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _25529_/Q _25530_/Q _17331_/C vssd1 vssd1 vccd1 vccd1 _17333_/B sky130_fd_sc_hd__and3_1
XFILLER_202_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _27295_/Q _26552_/Q _14544_/S vssd1 vssd1 vccd1 vccd1 _14543_/X sky130_fd_sc_hd__mux2_1
X_26529_ _27304_/CLK _26529_/D vssd1 vssd1 vccd1 vccd1 _26529_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17262_ _17259_/X _17263_/C _25509_/Q vssd1 vssd1 vccd1 vccd1 _17264_/B sky130_fd_sc_hd__a21oi_1
X_14474_ _26653_/Q _25693_/Q _14474_/S vssd1 vssd1 vccd1 vccd1 _14474_/X sky130_fd_sc_hd__mux2_1
X_19001_ _18003_/X _18984_/X _19000_/X _18927_/X vssd1 vssd1 vccd1 vccd1 _19001_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_16213_ _14601_/A _16211_/Y _16212_/X _15135_/X vssd1 vssd1 vccd1 vccd1 _16213_/X
+ sky130_fd_sc_hd__o22a_1
X_13425_ _15727_/S vssd1 vssd1 vccd1 vccd1 _13698_/A sky130_fd_sc_hd__buf_2
XFILLER_139_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17193_ _25490_/Q _20630_/B vssd1 vssd1 vccd1 vccd1 _17193_/X sky130_fd_sc_hd__or2_1
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16144_ _16142_/X _16143_/X _16144_/S vssd1 vssd1 vccd1 vccd1 _16144_/X sky130_fd_sc_hd__mux2_1
X_13356_ _13535_/S vssd1 vssd1 vccd1 vccd1 _15484_/S sky130_fd_sc_hd__buf_6
XFILLER_127_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16075_ _12772_/A _26895_/Q _26767_/Q _15623_/B vssd1 vssd1 vccd1 vccd1 _16075_/X
+ sky130_fd_sc_hd__a22o_1
X_13287_ _13675_/S vssd1 vssd1 vccd1 vccd1 _15582_/A sky130_fd_sc_hd__buf_4
XFILLER_143_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19903_ _19894_/X _19901_/X _19902_/X vssd1 vssd1 vccd1 vccd1 _19903_/X sky130_fd_sc_hd__a21o_1
X_15026_ _27257_/Q _15026_/B vssd1 vssd1 vccd1 vccd1 _15026_/X sky130_fd_sc_hd__or2_1
X_19834_ _25667_/Q _25666_/Q _19834_/C vssd1 vssd1 vccd1 vccd1 _19845_/B sky130_fd_sc_hd__and3_1
XFILLER_268_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19765_ _19941_/A vssd1 vssd1 vccd1 vccd1 _19765_/X sky130_fd_sc_hd__buf_2
X_16977_ _14716_/X _16952_/X _16887_/X vssd1 vssd1 vccd1 vccd1 _16980_/B sky130_fd_sc_hd__o21ai_2
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 coreIndex[4] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15928_ _15300_/A _15926_/X _15927_/X _13367_/A vssd1 vssd1 vccd1 vccd1 _15928_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18716_ _18895_/A vssd1 vssd1 vccd1 vccd1 _18716_/X sky130_fd_sc_hd__buf_2
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19696_ _25727_/Q vssd1 vssd1 vccd1 vccd1 _20630_/A sky130_fd_sc_hd__buf_4
XFILLER_271_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18647_ _19358_/A _18641_/Y _18642_/Y _19454_/A _18646_/X vssd1 vssd1 vccd1 vccd1
+ _18647_/X sky130_fd_sc_hd__o221a_1
XFILLER_65_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15859_ _15859_/A _15859_/B vssd1 vssd1 vccd1 vccd1 _15859_/X sky130_fd_sc_hd__or2_1
XFILLER_91_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18578_ _19231_/B _19849_/A vssd1 vssd1 vccd1 vccd1 _18580_/B sky130_fd_sc_hd__and2b_1
XFILLER_212_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17529_ _17529_/A vssd1 vssd1 vccd1 vccd1 _17529_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_205_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20540_ _20540_/A vssd1 vssd1 vccd1 vccd1 _25703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20471_ _20471_/A _20471_/B _20471_/C vssd1 vssd1 vccd1 vccd1 _20471_/Y sky130_fd_sc_hd__nand3_1
XFILLER_146_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22210_ _22210_/A vssd1 vssd1 vccd1 vccd1 _22226_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23190_ _26542_/Q _23108_/X _23194_/S vssd1 vssd1 vccd1 vccd1 _23191_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22141_ _26165_/Q _22113_/X _22140_/X input259/X _22137_/X vssd1 vssd1 vccd1 vccd1
+ _22141_/X sky130_fd_sc_hd__a221o_1
Xoutput320 _16771_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[23] sky130_fd_sc_hd__buf_2
Xoutput331 _16730_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[8] sky130_fd_sc_hd__buf_2
Xoutput342 _16900_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[17] sky130_fd_sc_hd__buf_2
Xoutput353 _16966_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[27] sky130_fd_sc_hd__buf_2
X_22072_ _22072_/A vssd1 vssd1 vccd1 vccd1 _26144_/D sky130_fd_sc_hd__clkbuf_1
Xoutput364 _16845_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[8] sky130_fd_sc_hd__buf_2
XFILLER_126_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput375 _20990_/B vssd1 vssd1 vccd1 vccd1 csb1[1] sky130_fd_sc_hd__buf_2
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21023_ _21023_/A vssd1 vssd1 vccd1 vccd1 _25881_/D sky130_fd_sc_hd__clkbuf_1
X_25900_ _27326_/CLK _25900_/D vssd1 vssd1 vccd1 vccd1 _25900_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput386 _17034_/X vssd1 vssd1 vccd1 vccd1 din0[19] sky130_fd_sc_hd__buf_2
XFILLER_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput397 _17047_/X vssd1 vssd1 vccd1 vccd1 din0[29] sky130_fd_sc_hd__buf_2
XFILLER_102_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26880_ _26880_/CLK _26880_/D vssd1 vssd1 vccd1 vccd1 _26880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25831_ _26240_/CLK _25831_/D vssd1 vssd1 vccd1 vccd1 _25831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25762_ _26592_/CLK _25762_/D vssd1 vssd1 vccd1 vccd1 _25762_/Q sky130_fd_sc_hd__dfxtp_1
X_22974_ _22974_/A vssd1 vssd1 vccd1 vccd1 _26460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_262_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24713_ _24722_/A _24713_/B vssd1 vssd1 vccd1 vccd1 _27085_/D sky130_fd_sc_hd__nor2_1
XFILLER_271_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21925_ _20554_/X _26079_/Q _21933_/S vssd1 vssd1 vccd1 vccd1 _21926_/A sky130_fd_sc_hd__mux2_1
XFILLER_262_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25693_ _26240_/CLK _25693_/D vssd1 vssd1 vccd1 vccd1 _25693_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_28_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24644_ _27069_/Q _24636_/X _24643_/X _24631_/X vssd1 vssd1 vccd1 vccd1 _27069_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21856_ _26056_/Q _20958_/X _21860_/S vssd1 vssd1 vccd1 vccd1 _21857_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20807_ _20807_/A vssd1 vssd1 vccd1 vccd1 _25799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24575_ _27046_/Q _24562_/X _24574_/Y _24567_/X vssd1 vssd1 vccd1 vccd1 _27046_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21787_ _20613_/X _26026_/Q _21787_/S vssd1 vssd1 vccd1 vccd1 _21788_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26314_ _26322_/CLK _26314_/D vssd1 vssd1 vccd1 vccd1 _26314_/Q sky130_fd_sc_hd__dfxtp_2
X_23526_ _23526_/A vssd1 vssd1 vccd1 vccd1 _23526_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20738_ _20738_/A vssd1 vssd1 vccd1 vccd1 _25766_/D sky130_fd_sc_hd__clkbuf_1
X_27294_ _27326_/CLK _27294_/D vssd1 vssd1 vccd1 vccd1 _27294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26245_ _26248_/CLK _26245_/D vssd1 vssd1 vccd1 vccd1 _26245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23457_ _23457_/A vssd1 vssd1 vccd1 vccd1 _26660_/D sky130_fd_sc_hd__clkbuf_1
X_20669_ _26278_/Q _20660_/X _20668_/X _20658_/X vssd1 vssd1 vccd1 vccd1 _25741_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13210_ _13210_/A vssd1 vssd1 vccd1 vccd1 _13529_/A sky130_fd_sc_hd__buf_4
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22408_ _22405_/A _22406_/X _22407_/X vssd1 vssd1 vccd1 vccd1 _22408_/Y sky130_fd_sc_hd__o21ai_1
X_26176_ _26238_/CLK _26176_/D vssd1 vssd1 vccd1 vccd1 _26176_/Q sky130_fd_sc_hd__dfxtp_1
X_14190_ _19455_/B _17856_/A _12803_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _17776_/A
+ sky130_fd_sc_hd__a211oi_4
X_23388_ _23434_/S vssd1 vssd1 vccd1 vccd1 _23397_/S sky130_fd_sc_hd__buf_6
XFILLER_109_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13141_ _13141_/A vssd1 vssd1 vccd1 vccd1 _13142_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_192_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25127_ _24736_/Y _25124_/X _25126_/Y _25109_/X vssd1 vssd1 vccd1 vccd1 _25127_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_124_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22339_ _22335_/Y _22336_/X _22338_/X _22330_/X vssd1 vssd1 vccd1 vccd1 _26225_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13072_ _13052_/X _13067_/X _13703_/A vssd1 vssd1 vccd1 vccd1 _13072_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25058_ _25159_/B vssd1 vssd1 vccd1 vccd1 _25058_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16900_ _16900_/A vssd1 vssd1 vccd1 vccd1 _16900_/X sky130_fd_sc_hd__clkbuf_1
X_24009_ _26877_/Q _23514_/X _24015_/S vssd1 vssd1 vccd1 vccd1 _24010_/A sky130_fd_sc_hd__mux2_1
XFILLER_279_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17880_ _17873_/X _17878_/X _18050_/S vssd1 vssd1 vccd1 vccd1 _17880_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16831_ _16834_/A _16895_/A _16878_/B vssd1 vssd1 vccd1 vccd1 _16832_/A sky130_fd_sc_hd__and3_2
XFILLER_238_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19550_ _19538_/X _19230_/X _19549_/X _19541_/X vssd1 vssd1 vccd1 vccd1 _25654_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16762_ _16762_/A vssd1 vssd1 vccd1 vccd1 _19118_/B sky130_fd_sc_hd__buf_4
X_13974_ _13239_/A _13972_/X _13973_/X _13540_/A vssd1 vssd1 vccd1 vccd1 _13974_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_58_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18501_ _18484_/X _18495_/Y _18500_/Y _18375_/X vssd1 vssd1 vccd1 vccd1 _18501_/X
+ sky130_fd_sc_hd__o31a_1
X_15713_ _13585_/A _26699_/Q _26827_/Q _15805_/S vssd1 vssd1 vccd1 vccd1 _15713_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_262_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12925_ _25921_/Q _12916_/X _12922_/Y _13928_/A vssd1 vssd1 vccd1 vccd1 _14237_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_74_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19481_ _25629_/Q _18719_/A _19480_/X _19352_/X vssd1 vssd1 vccd1 vccd1 _25629_/D
+ sky130_fd_sc_hd__o211a_1
X_16693_ _16769_/A vssd1 vssd1 vccd1 vccd1 _16693_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18432_ _25730_/Q _19772_/A _18432_/C vssd1 vssd1 vccd1 vccd1 _18530_/B sky130_fd_sc_hd__and3_1
XFILLER_262_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15644_ _15063_/A _26700_/Q _26828_/Q _16050_/B vssd1 vssd1 vccd1 vccd1 _15644_/X
+ sky130_fd_sc_hd__a22o_1
X_12856_ _12891_/A _12893_/A _17653_/C _12899_/A _25933_/Q vssd1 vssd1 vccd1 vccd1
+ _15706_/A sky130_fd_sc_hd__o32a_2
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _18858_/S _18207_/X _18271_/X vssd1 vssd1 vccd1 vccd1 _18363_/X sky130_fd_sc_hd__o21a_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _26637_/Q _26733_/Q _15582_/A vssd1 vssd1 vccd1 vccd1 _15576_/B sky130_fd_sc_hd__mux2_1
XFILLER_15_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _16635_/A vssd1 vssd1 vccd1 vccd1 _16996_/A sky130_fd_sc_hd__clkbuf_2
X_17314_ _25525_/Q _17314_/B vssd1 vssd1 vccd1 vccd1 _17322_/C sky130_fd_sc_hd__and2_1
XFILLER_159_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _25572_/Q _14187_/A _14193_/B vssd1 vssd1 vccd1 vccd1 _14526_/X sky130_fd_sc_hd__o21a_1
X_18294_ _27073_/Q _18815_/A _18816_/A _27171_/Q _18817_/A vssd1 vssd1 vccd1 vccd1
+ _18294_/X sky130_fd_sc_hd__a221o_1
XFILLER_230_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17245_ _24966_/A vssd1 vssd1 vccd1 vccd1 _17285_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14457_ _26909_/Q _26393_/Q _14472_/S vssd1 vssd1 vccd1 vccd1 _14457_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13408_ _14178_/S vssd1 vssd1 vccd1 vccd1 _13409_/A sky130_fd_sc_hd__clkbuf_2
X_17176_ _16540_/S _17170_/X _17174_/X _17175_/X vssd1 vssd1 vccd1 vccd1 _25484_/D
+ sky130_fd_sc_hd__o211a_1
X_14388_ _26522_/Q _26130_/Q _14389_/S vssd1 vssd1 vccd1 vccd1 _14388_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16127_ _16124_/Y _19016_/S _16125_/A vssd1 vssd1 vccd1 vccd1 _16127_/X sky130_fd_sc_hd__a21o_1
X_13339_ _13339_/A vssd1 vssd1 vccd1 vccd1 _13340_/A sky130_fd_sc_hd__buf_2
XFILLER_116_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16058_ _26507_/Q _26379_/Q _16069_/S vssd1 vssd1 vccd1 vccd1 _16058_/X sky130_fd_sc_hd__mux2_1
X_15009_ _15001_/X _15008_/X _17179_/A vssd1 vssd1 vccd1 vccd1 _15009_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_257_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19817_ _27138_/Q _27072_/Q _19785_/Y vssd1 vssd1 vccd1 vccd1 _19817_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19748_ _20712_/A vssd1 vssd1 vccd1 vccd1 _19748_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19679_ _27103_/Q _20079_/A _19905_/A _19678_/X vssd1 vssd1 vccd1 vccd1 _19679_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21710_ _25994_/Q _20973_/A _20986_/B _16669_/B _21662_/S vssd1 vssd1 vccd1 vccd1
+ _25994_/D sky130_fd_sc_hd__a41o_1
XFILLER_53_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22690_ _22690_/A vssd1 vssd1 vccd1 vccd1 _26342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21641_ _21641_/A _21641_/B vssd1 vssd1 vccd1 vccd1 _21641_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21572_ _25960_/Q _21506_/X _21571_/Y _21531_/X vssd1 vssd1 vccd1 vccd1 _25960_/D
+ sky130_fd_sc_hd__a211o_1
X_24360_ _24472_/A vssd1 vssd1 vccd1 vccd1 _24361_/S sky130_fd_sc_hd__buf_2
XFILLER_162_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20523_ _20523_/A vssd1 vssd1 vccd1 vccd1 _25699_/D sky130_fd_sc_hd__clkbuf_1
X_23311_ _20525_/X _26596_/Q _23313_/S vssd1 vssd1 vccd1 vccd1 _23312_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24291_ _24291_/A vssd1 vssd1 vccd1 vccd1 _24327_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_192_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26030_ _27265_/CLK _26030_/D vssd1 vssd1 vccd1 vccd1 _26030_/Q sky130_fd_sc_hd__dfxtp_2
X_23242_ _26565_/Q _23079_/X _23244_/S vssd1 vssd1 vccd1 vccd1 _23243_/A sky130_fd_sc_hd__mux2_1
X_20454_ _27131_/Q _19765_/X _24768_/A _20453_/Y vssd1 vssd1 vccd1 vccd1 _20454_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23173_ _23173_/A vssd1 vssd1 vccd1 vccd1 _26534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20385_ _20385_/A _20385_/B vssd1 vssd1 vccd1 vccd1 _20385_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22124_ _22179_/A vssd1 vssd1 vccd1 vccd1 _22124_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22055_ _26137_/Q _20900_/X _22055_/S vssd1 vssd1 vccd1 vccd1 _22056_/A sky130_fd_sc_hd__mux2_1
X_26932_ _26932_/CLK _26932_/D vssd1 vssd1 vccd1 vccd1 _26932_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21006_ _21063_/S vssd1 vssd1 vccd1 vccd1 _21015_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26863_ _27311_/CLK _26863_/D vssd1 vssd1 vccd1 vccd1 _26863_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25814_ _26843_/CLK _25814_/D vssd1 vssd1 vccd1 vccd1 _25814_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26794_ _27309_/CLK _26794_/D vssd1 vssd1 vccd1 vccd1 _26794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25745_ _26282_/CLK _25745_/D vssd1 vssd1 vccd1 vccd1 _25745_/Q sky130_fd_sc_hd__dfxtp_4
X_22957_ _22957_/A vssd1 vssd1 vccd1 vccd1 _26453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12710_ _25589_/Q vssd1 vssd1 vccd1 vccd1 _14268_/S sky130_fd_sc_hd__clkbuf_2
X_21908_ _21908_/A vssd1 vssd1 vccd1 vccd1 _26071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25676_ _26278_/CLK _25676_/D vssd1 vssd1 vccd1 vccd1 _25676_/Q sky130_fd_sc_hd__dfxtp_1
X_13690_ _18604_/S _13690_/B vssd1 vssd1 vccd1 vccd1 _13691_/A sky130_fd_sc_hd__or2_1
X_22888_ _26423_/Q _22742_/X _22888_/S vssd1 vssd1 vccd1 vccd1 _22889_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24627_ _24627_/A _24629_/B vssd1 vssd1 vccd1 vccd1 _24627_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21839_ _21839_/A vssd1 vssd1 vccd1 vccd1 _26048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15360_ _15142_/X _15354_/X _15359_/X _14660_/A vssd1 vssd1 vccd1 vccd1 _15360_/X
+ sky130_fd_sc_hd__a211o_1
X_24558_ _27040_/Q _24546_/X _24557_/Y _24551_/X vssd1 vssd1 vccd1 vccd1 _27040_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14311_ _13521_/A _26591_/Q _14365_/S _26331_/Q _14390_/S vssd1 vssd1 vccd1 vccd1
+ _14311_/X sky130_fd_sc_hd__o221a_1
XFILLER_196_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23509_ _24004_/B _23860_/B vssd1 vssd1 vccd1 vccd1 _23591_/A sky130_fd_sc_hd__nor2_2
X_27277_ _27277_/CLK _27277_/D vssd1 vssd1 vccd1 vccd1 _27277_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_184_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15291_ _12706_/A _16284_/S _15244_/X _15290_/Y vssd1 vssd1 vccd1 vccd1 _17793_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24489_ _27026_/Q _24480_/X _24488_/Y _24470_/X vssd1 vssd1 vccd1 vccd1 _27026_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17030_ _17028_/X _16893_/B _17025_/X input222/X vssd1 vssd1 vccd1 vccd1 _17030_/X
+ sky130_fd_sc_hd__a22o_4
X_26228_ _26520_/CLK _26228_/D vssd1 vssd1 vccd1 vccd1 _26228_/Q sky130_fd_sc_hd__dfxtp_1
X_14242_ _14237_/Y _14239_/Y _14241_/X _14602_/A _13558_/A vssd1 vssd1 vccd1 vccd1
+ _14242_/X sky130_fd_sc_hd__o221a_1
XFILLER_172_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14173_ _27235_/Q _14173_/B vssd1 vssd1 vccd1 vccd1 _14173_/X sky130_fd_sc_hd__or2_1
X_26159_ _26939_/CLK _26159_/D vssd1 vssd1 vccd1 vccd1 _26159_/Q sky130_fd_sc_hd__dfxtp_1
X_13124_ _13124_/A vssd1 vssd1 vccd1 vccd1 _13857_/A sky130_fd_sc_hd__buf_2
XFILLER_139_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18981_ _16043_/Y _18371_/X _18366_/A _16621_/B _17503_/X vssd1 vssd1 vccd1 vccd1
+ _18981_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_140_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13055_ _14344_/S vssd1 vssd1 vccd1 vccd1 _14114_/S sky130_fd_sc_hd__clkbuf_2
X_17932_ _17926_/X _17930_/X _18265_/S vssd1 vssd1 vccd1 vccd1 _17932_/X sky130_fd_sc_hd__mux2_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17863_ _17966_/A vssd1 vssd1 vccd1 vccd1 _18362_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19602_ _19658_/A _19659_/B vssd1 vssd1 vccd1 vccd1 _19607_/A sky130_fd_sc_hd__xnor2_2
XFILLER_282_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16814_ _16828_/A _16824_/B _16848_/B vssd1 vssd1 vccd1 vccd1 _16815_/A sky130_fd_sc_hd__and3_4
X_17794_ _15344_/A _17792_/X _17793_/X vssd1 vssd1 vccd1 vccd1 _17794_/X sky130_fd_sc_hd__o21a_1
XFILLER_4_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19533_ _19525_/X _18995_/X _19532_/X _19528_/X vssd1 vssd1 vccd1 vccd1 _25647_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_35_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16745_ _25674_/Q vssd1 vssd1 vccd1 vccd1 _22500_/A sky130_fd_sc_hd__clkbuf_4
X_13957_ _14389_/S vssd1 vssd1 vccd1 vccd1 _16005_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_35_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_199_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26739_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_222_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12908_ _12933_/B _12907_/Y _12872_/A vssd1 vssd1 vccd1 vccd1 _13923_/B sky130_fd_sc_hd__a21oi_2
X_19464_ _27132_/Q _18748_/X _19462_/X _19463_/X vssd1 vssd1 vccd1 vccd1 _19464_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_35_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16676_ _16676_/A _16676_/B vssd1 vssd1 vccd1 vccd1 _17020_/A sky130_fd_sc_hd__nor2_4
XFILLER_234_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13888_ _14431_/A vssd1 vssd1 vccd1 vccd1 _13889_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_128_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27058_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_261_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18415_ _18413_/Y _18414_/X _18896_/A vssd1 vssd1 vccd1 vccd1 _18415_/X sky130_fd_sc_hd__mux2_1
X_15627_ _27247_/Q _16073_/B vssd1 vssd1 vccd1 vccd1 _15627_/X sky130_fd_sc_hd__or2_1
XFILLER_22_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19395_ _18682_/X _18212_/X _18193_/B _18342_/A vssd1 vssd1 vccd1 vccd1 _19395_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12839_ _16657_/A _25792_/Q vssd1 vssd1 vccd1 vccd1 _13389_/A sky130_fd_sc_hd__nand2_2
XFILLER_61_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18346_ _18344_/Y _18345_/X _18487_/A vssd1 vssd1 vccd1 vccd1 _18346_/X sky130_fd_sc_hd__mux2_1
X_15558_ _12771_/A _26701_/Q _26829_/Q _15548_/S vssd1 vssd1 vccd1 vccd1 _15558_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14509_ _14502_/X _14508_/X _14421_/A vssd1 vssd1 vccd1 vccd1 _14509_/X sky130_fd_sc_hd__o21a_1
XFILLER_147_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18277_ _18602_/A _19358_/B _18276_/X _17503_/X vssd1 vssd1 vccd1 vccd1 _18277_/X
+ sky130_fd_sc_hd__o211a_1
X_15489_ _15488_/X _26702_/Q _26830_/Q _15834_/S _15486_/A vssd1 vssd1 vccd1 vccd1
+ _15489_/X sky130_fd_sc_hd__a221o_1
XFILLER_238_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17228_ _25176_/A vssd1 vssd1 vccd1 vccd1 _25027_/A sky130_fd_sc_hd__buf_4
Xinput30 core_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_1
Xinput41 core_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_1
XFILLER_238_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput52 dout0[18] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_2
Xinput63 dout0[28] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_2
X_17159_ _17224_/B vssd1 vssd1 vccd1 vccd1 _17159_/X sky130_fd_sc_hd__clkbuf_2
Xinput74 dout0[38] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__clkbuf_1
Xinput85 dout0[48] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__clkbuf_1
Xinput96 dout0[58] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_5_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_192_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20170_ _25743_/Q vssd1 vssd1 vccd1 vccd1 _20675_/A sky130_fd_sc_hd__buf_8
XFILLER_170_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23860_ _23860_/A _23860_/B vssd1 vssd1 vccd1 vccd1 _23917_/A sky130_fd_sc_hd__or2_4
XFILLER_272_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22811_ _26389_/Q _22736_/X _22811_/S vssd1 vssd1 vccd1 vccd1 _22812_/A sky130_fd_sc_hd__mux2_1
XFILLER_272_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23791_ _23684_/X _26780_/Q _23799_/S vssd1 vssd1 vccd1 vccd1 _23792_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25530_ _25553_/CLK _25530_/D vssd1 vssd1 vccd1 vccd1 _25530_/Q sky130_fd_sc_hd__dfxtp_1
X_22742_ _23785_/A vssd1 vssd1 vccd1 vccd1 _22742_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_213_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25461_ _23782_/X _27325_/Q _25463_/S vssd1 vssd1 vccd1 vccd1 _25462_/A sky130_fd_sc_hd__mux2_1
X_22673_ _26337_/Q _22672_/X _22673_/S vssd1 vssd1 vccd1 vccd1 _22674_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27200_ _27203_/CLK _27200_/D vssd1 vssd1 vccd1 vccd1 _27200_/Q sky130_fd_sc_hd__dfxtp_1
X_24412_ _24381_/X _25606_/Q _24411_/X vssd1 vssd1 vccd1 vccd1 _24674_/B sky130_fd_sc_hd__o21a_4
X_21624_ _21276_/A _21623_/X _21603_/X vssd1 vssd1 vccd1 vccd1 _21624_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_179_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25392_ _25392_/A vssd1 vssd1 vccd1 vccd1 _27294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27131_ _27132_/CLK _27131_/D vssd1 vssd1 vccd1 vccd1 _27131_/Q sky130_fd_sc_hd__dfxtp_4
X_24343_ _21203_/A _25496_/Q _17471_/A _24342_/Y vssd1 vssd1 vccd1 vccd1 _24347_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_138_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21555_ _21552_/X _25864_/Q _21554_/Y _21518_/X vssd1 vssd1 vccd1 vccd1 _21555_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20506_ _20506_/A vssd1 vssd1 vccd1 vccd1 _25695_/D sky130_fd_sc_hd__clkbuf_1
X_27062_ _27062_/CLK _27062_/D vssd1 vssd1 vccd1 vccd1 _27062_/Q sky130_fd_sc_hd__dfxtp_2
X_24274_ _26981_/Q _24275_/C _26982_/Q vssd1 vssd1 vccd1 vccd1 _24276_/B sky130_fd_sc_hd__a21oi_1
X_21486_ _20670_/A _21481_/X _21459_/X _21485_/X vssd1 vssd1 vccd1 vccd1 _21486_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26013_ _26796_/CLK _26013_/D vssd1 vssd1 vccd1 vccd1 _26013_/Q sky130_fd_sc_hd__dfxtp_1
X_23225_ _26557_/Q _23053_/X _23233_/S vssd1 vssd1 vccd1 vccd1 _23226_/A sky130_fd_sc_hd__mux2_1
X_20437_ _20433_/X _20434_/Y _20435_/Y _19787_/A vssd1 vssd1 vccd1 vccd1 _20437_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_162_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23156_ _23156_/A vssd1 vssd1 vccd1 vccd1 _26526_/D sky130_fd_sc_hd__clkbuf_1
X_20368_ _27159_/Q _27093_/Q vssd1 vssd1 vccd1 vccd1 _20369_/B sky130_fd_sc_hd__nand2_1
X_22107_ _22230_/C _22236_/C _26230_/Q vssd1 vssd1 vccd1 vccd1 _22239_/B sky130_fd_sc_hd__o21ai_2
X_23087_ _26503_/Q _23085_/X _23099_/S vssd1 vssd1 vccd1 vccd1 _23088_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20299_ _20299_/A _20299_/B vssd1 vssd1 vccd1 vccd1 _20300_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22038_ _26129_/Q _20875_/X _22044_/S vssd1 vssd1 vccd1 vccd1 _22039_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26915_ _26916_/CLK _26915_/D vssd1 vssd1 vccd1 vccd1 _26915_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26846_ _27297_/CLK _26846_/D vssd1 vssd1 vccd1 vccd1 _26846_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14860_ _25898_/Q _15026_/B vssd1 vssd1 vccd1 vccd1 _14860_/X sky130_fd_sc_hd__or2_1
XFILLER_102_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13811_ _16015_/A _13811_/B vssd1 vssd1 vccd1 vccd1 _13811_/X sky130_fd_sc_hd__or2_1
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26777_ _26905_/CLK _26777_/D vssd1 vssd1 vccd1 vccd1 _26777_/Q sky130_fd_sc_hd__dfxtp_1
X_14791_ _14791_/A vssd1 vssd1 vccd1 vccd1 _14792_/A sky130_fd_sc_hd__buf_2
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23989_ _23989_/A vssd1 vssd1 vccd1 vccd1 _23998_/S sky130_fd_sc_hd__buf_4
XFILLER_244_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16530_ _27326_/Q _26583_/Q _16533_/A vssd1 vssd1 vccd1 vccd1 _16530_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13742_ _14133_/A _13742_/B vssd1 vssd1 vccd1 vccd1 _13742_/Y sky130_fd_sc_hd__nor2_1
X_25728_ _26271_/CLK _25728_/D vssd1 vssd1 vccd1 vccd1 _25728_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16461_ _16461_/A _16461_/B vssd1 vssd1 vccd1 vccd1 _16462_/B sky130_fd_sc_hd__nand2_1
X_25659_ _26248_/CLK _25659_/D vssd1 vssd1 vccd1 vccd1 _25659_/Q sky130_fd_sc_hd__dfxtp_1
X_13673_ _12738_/D _26885_/Q _26757_/Q _15931_/S _14768_/A vssd1 vssd1 vccd1 vccd1
+ _13673_/X sky130_fd_sc_hd__a221o_1
XFILLER_189_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18200_ _17939_/X _17926_/X _18265_/S vssd1 vssd1 vccd1 vccd1 _18200_/X sky130_fd_sc_hd__mux2_1
X_15412_ _15227_/S _15407_/X _15411_/X _14786_/A vssd1 vssd1 vccd1 vccd1 _15412_/X
+ sky130_fd_sc_hd__a31o_1
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19180_ _19246_/C _19180_/B vssd1 vssd1 vccd1 vccd1 _20251_/A sky130_fd_sc_hd__or2_2
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16392_ _26679_/Q _25719_/Q _16402_/S vssd1 vssd1 vccd1 vccd1 _16392_/X sky130_fd_sc_hd__mux2_1
XPHY_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18131_ _18468_/A vssd1 vssd1 vccd1 vccd1 _18574_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15343_ _19158_/S _15343_/B vssd1 vssd1 vccd1 vccd1 _15344_/A sky130_fd_sc_hd__nor2_1
X_27329_ _27329_/A vssd1 vssd1 vccd1 vccd1 _27329_/X sky130_fd_sc_hd__buf_2
XPHY_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18062_ _17954_/X _17902_/X _18062_/S vssd1 vssd1 vccd1 vccd1 _18062_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15274_ _15165_/X _15271_/X _15273_/X vssd1 vssd1 vccd1 vccd1 _15274_/X sky130_fd_sc_hd__o21a_1
XFILLER_145_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17013_ _17016_/A vssd1 vssd1 vccd1 vccd1 _17013_/X sky130_fd_sc_hd__clkbuf_2
X_14225_ _13937_/X _26592_/Q _16004_/S _26332_/Q _13653_/S vssd1 vssd1 vccd1 vccd1
+ _14225_/X sky130_fd_sc_hd__o221a_1
XFILLER_256_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14156_ _14165_/A _14156_/B vssd1 vssd1 vccd1 vccd1 _14156_/Y sky130_fd_sc_hd__nand2_1
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13107_ _13107_/A vssd1 vssd1 vccd1 vccd1 _14713_/C sky130_fd_sc_hd__buf_2
X_14087_ _26101_/Q _26002_/Q _14095_/A vssd1 vssd1 vccd1 vccd1 _14087_/X sky130_fd_sc_hd__mux2_1
X_18964_ _25740_/Q _18964_/B vssd1 vssd1 vccd1 vccd1 _18965_/B sky130_fd_sc_hd__nor2_1
XFILLER_113_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13038_ _12771_/A _26695_/Q _26823_/Q _15561_/B vssd1 vssd1 vccd1 vccd1 _13038_/X
+ sky130_fd_sc_hd__a22o_1
X_17915_ _17905_/X _17913_/X _18318_/S vssd1 vssd1 vccd1 vccd1 _17915_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18895_ _18895_/A vssd1 vssd1 vccd1 vccd1 _18895_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_267_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17846_ _17846_/A _17846_/B _17846_/C _17846_/D vssd1 vssd1 vccd1 vccd1 _17846_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_208_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17777_ _18339_/A vssd1 vssd1 vccd1 vccd1 _19219_/A sky130_fd_sc_hd__buf_2
X_14989_ _14890_/X _26904_/Q _26776_/Q _14981_/S _14772_/A vssd1 vssd1 vccd1 vccd1
+ _14989_/X sky130_fd_sc_hd__a221o_1
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19516_ _19512_/X _18663_/X _19514_/X _19515_/X vssd1 vssd1 vccd1 vccd1 _25640_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16728_ _18549_/S _16728_/B vssd1 vssd1 vccd1 vccd1 _18539_/A sky130_fd_sc_hd__or2_2
XINSDIODE2_520 _17023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_531 _17048_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_542 _25753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19447_ _18891_/X _19422_/X _19446_/X _18929_/X vssd1 vssd1 vccd1 vccd1 _19448_/B
+ sky130_fd_sc_hd__a22o_1
X_16659_ _20796_/B vssd1 vssd1 vccd1 vccd1 _20973_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_263_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_553 _20990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19378_ _18003_/X _19362_/X _19377_/X _18841_/X vssd1 vssd1 vccd1 vccd1 _19378_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_210_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18329_ _18329_/A _18904_/A vssd1 vssd1 vccd1 vccd1 _18329_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21340_ _21337_/Y _21339_/Y _21297_/X vssd1 vssd1 vccd1 vccd1 _21340_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_108_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_96_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27295_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_135_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21271_ _21271_/A _21271_/B vssd1 vssd1 vccd1 vccd1 _21271_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_25_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27293_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_265_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20222_ _22130_/A vssd1 vssd1 vccd1 vccd1 _22638_/B sky130_fd_sc_hd__buf_12
XFILLER_144_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23010_ _23010_/A vssd1 vssd1 vccd1 vccd1 _26476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20153_ _19833_/X _20164_/B _20152_/Y _20100_/X vssd1 vssd1 vccd1 vccd1 _20154_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_134_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24961_ _27153_/Q _24953_/X _24960_/Y _24949_/X vssd1 vssd1 vccd1 vccd1 _27153_/D
+ sky130_fd_sc_hd__o211a_1
X_20084_ _20084_/A _20084_/B vssd1 vssd1 vccd1 vccd1 _20084_/Y sky130_fd_sc_hd__nand2_1
XFILLER_258_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26700_ _27314_/CLK _26700_/D vssd1 vssd1 vccd1 vccd1 _26700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_258_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23912_ _23912_/A vssd1 vssd1 vccd1 vccd1 _26834_/D sky130_fd_sc_hd__clkbuf_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24892_ _24890_/Y _24891_/X _21242_/X vssd1 vssd1 vccd1 vccd1 _27130_/D sky130_fd_sc_hd__a21oi_1
XFILLER_273_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26631_ _27330_/A _26631_/D vssd1 vssd1 vccd1 vccd1 _26631_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23843_ _23763_/X _26804_/Q _23843_/S vssd1 vssd1 vccd1 vccd1 _23844_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26562_ _26599_/CLK _26562_/D vssd1 vssd1 vccd1 vccd1 _26562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23774_ _23773_/X _26775_/Q _23780_/S vssd1 vssd1 vccd1 vccd1 _23775_/A sky130_fd_sc_hd__mux2_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20986_ _26587_/Q _20986_/B _20986_/C vssd1 vssd1 vccd1 vccd1 _20987_/A sky130_fd_sc_hd__and3_1
XFILLER_26_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25513_ _27049_/CLK _25513_/D vssd1 vssd1 vccd1 vccd1 _25513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22725_ _26353_/Q _22723_/X _22737_/S vssd1 vssd1 vccd1 vccd1 _22726_/A sky130_fd_sc_hd__mux2_1
X_26493_ _26751_/CLK _26493_/D vssd1 vssd1 vccd1 vccd1 _26493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25444_ _23757_/X _27317_/Q _25448_/S vssd1 vssd1 vccd1 vccd1 _25445_/A sky130_fd_sc_hd__mux2_1
X_22656_ _23699_/A vssd1 vssd1 vccd1 vccd1 _22656_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_179_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21607_ _21552_/X _21566_/X _21606_/Y _21581_/X vssd1 vssd1 vccd1 vccd1 _21607_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_178_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25375_ _25375_/A vssd1 vssd1 vccd1 vccd1 _27286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_279_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22587_ _22600_/A vssd1 vssd1 vccd1 vccd1 _22587_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27114_ _27117_/CLK _27114_/D vssd1 vssd1 vccd1 vccd1 _27114_/Q sky130_fd_sc_hd__dfxtp_4
X_24326_ _27000_/Q _26999_/Q _24326_/C vssd1 vssd1 vccd1 vccd1 _24331_/C sky130_fd_sc_hd__and3_1
X_21538_ _21480_/X _21536_/X _21537_/X vssd1 vssd1 vccd1 vccd1 _21538_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_139_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27045_ _27049_/CLK _27045_/D vssd1 vssd1 vccd1 vccd1 _27045_/Q sky130_fd_sc_hd__dfxtp_1
X_24257_ _26975_/Q _24258_/C _26976_/Q vssd1 vssd1 vccd1 vccd1 _24259_/B sky130_fd_sc_hd__a21oi_1
XFILLER_107_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21469_ _25485_/Q _21495_/B vssd1 vssd1 vccd1 vccd1 _21469_/X sky130_fd_sc_hd__or2_1
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _14008_/X _14009_/X _14010_/S vssd1 vssd1 vccd1 vccd1 _14010_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23208_ _23208_/A vssd1 vssd1 vccd1 vccd1 _26550_/D sky130_fd_sc_hd__clkbuf_1
X_24188_ _24188_/A _24188_/B vssd1 vssd1 vccd1 vccd1 _24188_/Y sky130_fd_sc_hd__nor2_1
XFILLER_150_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23139_ _23139_/A _25393_/A vssd1 vssd1 vccd1 vccd1 _23196_/A sky130_fd_sc_hd__nor2_4
XFILLER_150_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15961_ _26920_/Q _15961_/B vssd1 vssd1 vccd1 vccd1 _15961_/X sky130_fd_sc_hd__or2_1
XFILLER_122_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput220 localMemory_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input220/X sky130_fd_sc_hd__buf_6
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput231 localMemory_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 input231/X sky130_fd_sc_hd__buf_8
XTAP_5442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput242 localMemory_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input242/X sky130_fd_sc_hd__buf_6
X_17700_ _20189_/A _17465_/A _17706_/A vssd1 vssd1 vccd1 vccd1 _17736_/B sky130_fd_sc_hd__mux2_1
X_14912_ _15088_/S vssd1 vssd1 vccd1 vccd1 _14996_/S sky130_fd_sc_hd__buf_2
XFILLER_76_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput253 manufacturerID[0] vssd1 vssd1 vccd1 vccd1 input253/X sky130_fd_sc_hd__buf_2
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15892_ _15982_/S _15890_/X _15891_/X _13614_/A vssd1 vssd1 vccd1 vccd1 _15892_/X
+ sky130_fd_sc_hd__o211a_1
X_18680_ _17824_/A _13380_/Y _18366_/X vssd1 vssd1 vccd1 vccd1 _18680_/Y sky130_fd_sc_hd__a21oi_1
Xinput264 partID[0] vssd1 vssd1 vccd1 vccd1 input264/X sky130_fd_sc_hd__clkbuf_1
XFILLER_276_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput275 partID[5] vssd1 vssd1 vccd1 vccd1 input275/X sky130_fd_sc_hd__clkbuf_1
XTAP_5486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_264_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17631_ _25927_/Q _17554_/A _13561_/Y _17577_/X vssd1 vssd1 vccd1 vccd1 _17631_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_14843_ _16384_/S vssd1 vssd1 vccd1 vccd1 _14878_/S sky130_fd_sc_hd__buf_2
XFILLER_236_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26829_ _27312_/CLK _26829_/D vssd1 vssd1 vccd1 vccd1 _26829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_252_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17562_ _25572_/Q _17529_/X _17540_/X _17561_/Y vssd1 vssd1 vccd1 vccd1 _17563_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14774_ _16513_/A _26714_/Q _26842_/Q _14767_/S _14773_/X vssd1 vssd1 vccd1 vccd1
+ _14774_/X sky130_fd_sc_hd__a221o_1
XFILLER_263_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16513_ _16513_/A vssd1 vssd1 vccd1 vccd1 _16513_/X sky130_fd_sc_hd__clkbuf_4
X_19301_ _27127_/Q _18812_/X _19299_/X _19300_/X vssd1 vssd1 vccd1 vccd1 _19301_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_216_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13725_ _13086_/X _26596_/Q _15634_/S _26336_/Q _15547_/A vssd1 vssd1 vccd1 vccd1
+ _13725_/X sky130_fd_sc_hd__o221a_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17493_ _21219_/A _21208_/D _21219_/B vssd1 vssd1 vccd1 vccd1 _21221_/A sky130_fd_sc_hd__or3_1
XFILLER_205_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16444_ _15321_/X _26903_/Q _26775_/Q _15228_/S _15210_/X vssd1 vssd1 vccd1 vccd1
+ _16444_/X sky130_fd_sc_hd__a221o_1
X_19232_ _18608_/X _19230_/X _19231_/Y vssd1 vssd1 vccd1 vccd1 _19234_/B sky130_fd_sc_hd__a21oi_1
X_13656_ _14060_/A vssd1 vssd1 vccd1 vccd1 _13657_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19163_ _27221_/Q _19299_/B vssd1 vssd1 vccd1 vccd1 _19163_/X sky130_fd_sc_hd__and2_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16375_ _19237_/A _16572_/B _19277_/A _16374_/X vssd1 vssd1 vccd1 vccd1 _16567_/B
+ sky130_fd_sc_hd__a31o_2
X_13587_ _13585_/X _26597_/Q _13065_/A _13586_/X vssd1 vssd1 vccd1 vccd1 _13587_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18114_ _27006_/Q _18238_/A _19060_/A _27102_/Q _18113_/X vssd1 vssd1 vccd1 vccd1
+ _18114_/X sky130_fd_sc_hd__a221o_1
XFILLER_158_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15326_ _15834_/S vssd1 vssd1 vccd1 vccd1 _16256_/B sky130_fd_sc_hd__clkbuf_4
X_19094_ _27025_/Q _18514_/A _19093_/X _18455_/A vssd1 vssd1 vccd1 vccd1 _19094_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18045_ _17974_/Y _18044_/X _18197_/S vssd1 vssd1 vccd1 vccd1 _18045_/X sky130_fd_sc_hd__mux2_1
X_15257_ _26866_/Q _25780_/Q _16301_/S vssd1 vssd1 vccd1 vccd1 _15257_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14208_ _26524_/Q _26132_/Q _15292_/A vssd1 vssd1 vccd1 vccd1 _14208_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15188_ _16405_/A _15182_/X _15186_/Y _15187_/X vssd1 vssd1 vccd1 vccd1 _15188_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14139_ input127/X input163/X _14402_/S vssd1 vssd1 vccd1 vccd1 _14139_/X sky130_fd_sc_hd__mux2_8
XFILLER_99_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19996_ _27144_/Q _27078_/Q _19959_/Y vssd1 vssd1 vccd1 vccd1 _19996_/X sky130_fd_sc_hd__a21o_1
XFILLER_113_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18947_ _18947_/A _18947_/B vssd1 vssd1 vccd1 vccd1 _18947_/Y sky130_fd_sc_hd__nor2_1
XFILLER_274_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18878_ _20034_/A _19442_/B vssd1 vssd1 vccd1 vccd1 _18878_/Y sky130_fd_sc_hd__nor2_1
XFILLER_251_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_143_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26940_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_251_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17829_ _17829_/A _16038_/B vssd1 vssd1 vccd1 vccd1 _18855_/B sky130_fd_sc_hd__or2b_1
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20840_ _25816_/Q vssd1 vssd1 vccd1 vccd1 _20841_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_54_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20771_ _20771_/A vssd1 vssd1 vccd1 vccd1 _25781_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_350 _19612_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_361 input228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22510_ _22510_/A vssd1 vssd1 vccd1 vccd1 _26279_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_372 _17064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_383 _16661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23490_ _23490_/A vssd1 vssd1 vccd1 vccd1 _26675_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_394 _17034_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22441_ _24441_/A vssd1 vssd1 vccd1 vccd1 _24415_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_195_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25160_ _27196_/Q _25151_/B _25158_/X _25159_/Y _22380_/X vssd1 vssd1 vccd1 vccd1
+ _27196_/D sky130_fd_sc_hd__o221a_1
X_22372_ _22372_/A vssd1 vssd1 vccd1 vccd1 _26234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24111_ _24133_/A vssd1 vssd1 vccd1 vccd1 _24120_/S sky130_fd_sc_hd__buf_2
XFILLER_163_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21323_ _21284_/X _18471_/X _21286_/X _25803_/Q _21322_/X vssd1 vssd1 vccd1 vccd1
+ _21323_/X sky130_fd_sc_hd__a221o_1
X_25091_ _27182_/Q _25085_/X _25090_/X vssd1 vssd1 vccd1 vccd1 _27182_/D sky130_fd_sc_hd__o21ba_1
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21254_ _21248_/X _21252_/X _21589_/A vssd1 vssd1 vccd1 vccd1 _21254_/X sky130_fd_sc_hd__a21o_1
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24042_ _26892_/Q _23562_/X _24048_/S vssd1 vssd1 vccd1 vccd1 _24043_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20205_ _20301_/A _20205_/B vssd1 vssd1 vccd1 vccd1 _20206_/C sky130_fd_sc_hd__and2b_1
X_21185_ _21188_/A _21185_/B vssd1 vssd1 vccd1 vccd1 _21186_/A sky130_fd_sc_hd__or2_1
XFILLER_132_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20136_ _20461_/S vssd1 vssd1 vccd1 vccd1 _20371_/S sky130_fd_sc_hd__buf_2
X_25993_ _27327_/CLK _25993_/D vssd1 vssd1 vccd1 vccd1 _25993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24944_ _24944_/A _24951_/B vssd1 vssd1 vccd1 vccd1 _24944_/Y sky130_fd_sc_hd__nand2_1
XINSDIODE2_10 _18693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20067_ _20067_/A _20067_/B _20067_/C vssd1 vssd1 vccd1 vccd1 _20067_/X sky130_fd_sc_hd__or3_1
XFILLER_219_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_21 _19099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_32 _19308_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_43 _19574_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_54 _20643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24875_ _20687_/A _19905_/X _24746_/Y _24896_/B vssd1 vssd1 vccd1 vccd1 _24875_/X
+ sky130_fd_sc_hd__o22a_1
XINSDIODE2_65 _20654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_76 _20694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_87 _21878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26614_ _27321_/CLK _26614_/D vssd1 vssd1 vccd1 vccd1 _26614_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_98 _21453_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23826_ _23738_/X _26796_/Q _23832_/S vssd1 vssd1 vccd1 vccd1 _23827_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26545_ _27259_/CLK _26545_/D vssd1 vssd1 vccd1 vccd1 _26545_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23757_ _23757_/A vssd1 vssd1 vccd1 vccd1 _23757_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20969_ _20969_/A vssd1 vssd1 vccd1 vccd1 _25859_/D sky130_fd_sc_hd__clkbuf_1
X_13510_ _27305_/Q _26562_/Q _13535_/S vssd1 vssd1 vccd1 vccd1 _13510_/X sky130_fd_sc_hd__mux2_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22708_ _22724_/A vssd1 vssd1 vccd1 vccd1 _22721_/S sky130_fd_sc_hd__clkbuf_4
X_14490_ _25902_/Q _13922_/B _14489_/Y _13928_/A vssd1 vssd1 vccd1 vccd1 _14490_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_26476_ _26609_/CLK _26476_/D vssd1 vssd1 vccd1 vccd1 _26476_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23688_ _23684_/X _26748_/Q _23700_/S vssd1 vssd1 vccd1 vccd1 _23689_/A sky130_fd_sc_hd__mux2_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25427_ _25427_/A vssd1 vssd1 vccd1 vccd1 _27309_/D sky130_fd_sc_hd__clkbuf_1
X_13441_ _26662_/Q _25702_/Q _13441_/S vssd1 vssd1 vccd1 vccd1 _13441_/X sky130_fd_sc_hd__mux2_1
X_22639_ _22639_/A vssd1 vssd1 vccd1 vccd1 _26327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16160_ _16320_/S _16160_/B vssd1 vssd1 vccd1 vccd1 _16160_/X sky130_fd_sc_hd__or2_1
X_25358_ _25358_/A vssd1 vssd1 vccd1 vccd1 _27278_/D sky130_fd_sc_hd__clkbuf_1
X_13372_ _23546_/A _14789_/A _15127_/A _13371_/Y vssd1 vssd1 vccd1 vccd1 _19947_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_103_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15111_ _15111_/A vssd1 vssd1 vccd1 vccd1 _15111_/X sky130_fd_sc_hd__buf_2
XFILLER_127_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24309_ _26994_/Q _26993_/Q _24309_/C vssd1 vssd1 vccd1 vccd1 _24311_/B sky130_fd_sc_hd__and3_1
XFILLER_127_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16091_ _13267_/X _26895_/Q _26767_/Q _16189_/S _13221_/A vssd1 vssd1 vccd1 vccd1
+ _16091_/X sky130_fd_sc_hd__a221o_1
XFILLER_127_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25289_ _23741_/X _27248_/Q _25293_/S vssd1 vssd1 vccd1 vccd1 _25290_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27028_ _27154_/CLK _27028_/D vssd1 vssd1 vccd1 vccd1 _27028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15042_ _15020_/X _15033_/X _15041_/X _14679_/A vssd1 vssd1 vccd1 vccd1 _15042_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19850_ _20252_/B _18582_/X _19671_/A _19849_/X vssd1 vssd1 vccd1 vccd1 _19850_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_150_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18801_ _18734_/A _18643_/A _18801_/S vssd1 vssd1 vccd1 vccd1 _18801_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19781_ _19766_/X _19778_/Y _19780_/X vssd1 vssd1 vccd1 vccd1 _19781_/X sky130_fd_sc_hd__a21o_1
X_16993_ _22478_/A _16988_/X _16990_/X _18329_/A vssd1 vssd1 vccd1 vccd1 _16993_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_283_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18732_ _18362_/X _18260_/X _18364_/X vssd1 vssd1 vccd1 vccd1 _18732_/Y sky130_fd_sc_hd__o21ai_1
XTAP_5250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15944_ _15940_/X _15943_/X _13313_/A vssd1 vssd1 vccd1 vccd1 _15944_/X sky130_fd_sc_hd__o21a_2
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18663_ _18437_/X _18652_/X _18662_/X vssd1 vssd1 vccd1 vccd1 _18663_/X sky130_fd_sc_hd__a21o_4
X_15875_ _12871_/A _15872_/Y _15873_/Y _13575_/X _15874_/X vssd1 vssd1 vccd1 vccd1
+ _15875_/X sky130_fd_sc_hd__o32a_1
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826_ _14826_/A vssd1 vssd1 vccd1 vccd1 _14827_/A sky130_fd_sc_hd__buf_8
X_17614_ _17712_/B _17612_/X _17608_/X _17613_/X vssd1 vssd1 vccd1 vccd1 _17615_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18594_ _18634_/B _18594_/B vssd1 vssd1 vccd1 vccd1 _19573_/B sky130_fd_sc_hd__nor2_1
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ _17653_/A _17556_/B _17545_/C vssd1 vssd1 vccd1 vccd1 _17545_/X sky130_fd_sc_hd__or3_1
X_14757_ _14757_/A vssd1 vssd1 vccd1 vccd1 _14758_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_17_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13708_ _15464_/B vssd1 vssd1 vccd1 vccd1 _15548_/S sky130_fd_sc_hd__clkbuf_4
X_17476_ _21244_/A _22536_/A vssd1 vssd1 vccd1 vccd1 _17476_/Y sky130_fd_sc_hd__nor2_1
X_14688_ _14688_/A vssd1 vssd1 vccd1 vccd1 _16484_/A sky130_fd_sc_hd__buf_2
XFILLER_189_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19215_ _18144_/A _19187_/X _19214_/X vssd1 vssd1 vccd1 vccd1 _19215_/Y sky130_fd_sc_hd__o21ai_4
X_13639_ _27272_/Q _26465_/Q _15923_/S vssd1 vssd1 vccd1 vccd1 _13639_/X sky130_fd_sc_hd__mux2_1
X_16427_ _16425_/X _16426_/X _16442_/S vssd1 vssd1 vccd1 vccd1 _16427_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19146_ _25745_/Q _25744_/Q _19146_/C vssd1 vssd1 vccd1 vccd1 _19179_/B sky130_fd_sc_hd__and3_1
X_16358_ _26089_/Q _25894_/Q _16359_/S vssd1 vssd1 vccd1 vccd1 _16358_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15309_ _15297_/X _15301_/X _15305_/X _15308_/X _14758_/A _14778_/A vssd1 vssd1 vccd1
+ vccd1 _15310_/B sky130_fd_sc_hd__mux4_1
X_16289_ _16289_/A vssd1 vssd1 vccd1 vccd1 _19191_/B sky130_fd_sc_hd__buf_4
X_19077_ _19482_/B _19074_/Y _19075_/X _19045_/Y _19076_/X vssd1 vssd1 vccd1 vccd1
+ _19077_/X sky130_fd_sc_hd__o32a_2
XFILLER_246_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18028_ _18028_/A _18028_/B vssd1 vssd1 vccd1 vccd1 _19879_/A sky130_fd_sc_hd__or2_4
XFILLER_246_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_259_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19979_ _19919_/B _19951_/A _19976_/Y _19977_/X _19978_/X vssd1 vssd1 vccd1 vccd1
+ _19982_/B sky130_fd_sc_hd__a311o_1
XFILLER_99_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22990_ _22990_/A vssd1 vssd1 vccd1 vccd1 _26467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21941_ _21941_/A vssd1 vssd1 vccd1 vccd1 _26086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24660_ _24740_/A vssd1 vssd1 vccd1 vccd1 _24660_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_282_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21872_ _26295_/Q _21869_/X _21871_/X input237/X vssd1 vssd1 vccd1 vccd1 _21872_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23611_ _23611_/A vssd1 vssd1 vccd1 vccd1 _26715_/D sky130_fd_sc_hd__clkbuf_1
X_20823_ _20823_/A vssd1 vssd1 vccd1 vccd1 _25807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24591_ _27052_/Q _24589_/X _24590_/Y _24580_/X vssd1 vssd1 vccd1 vccd1 _27052_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_270_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26330_ _27266_/CLK _26330_/D vssd1 vssd1 vccd1 vccd1 _26330_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23542_ _23542_/A vssd1 vssd1 vccd1 vccd1 _23542_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_196_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20754_ _20754_/A vssd1 vssd1 vccd1 vccd1 _25773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_180 _13747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_191 _15902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26261_ _26264_/CLK _26261_/D vssd1 vssd1 vccd1 vccd1 _26261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23473_ _23473_/A vssd1 vssd1 vccd1 vccd1 _26667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20685_ _26284_/Q _20673_/X _20683_/X _20684_/X vssd1 vssd1 vccd1 vccd1 _25747_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_40_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26925_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_25212_ _27054_/Q _21874_/A input178/X _25209_/X _25199_/A vssd1 vssd1 vccd1 vccd1
+ _25212_/X sky130_fd_sc_hd__a41o_1
X_22424_ _26194_/Q _22418_/X _22423_/X _22348_/X vssd1 vssd1 vccd1 vccd1 _26242_/D
+ sky130_fd_sc_hd__o211a_1
X_26192_ _26222_/CLK _26192_/D vssd1 vssd1 vccd1 vccd1 _26192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25143_ _25143_/A _25151_/B vssd1 vssd1 vccd1 vccd1 _25143_/Y sky130_fd_sc_hd__nand2_1
X_22355_ _22515_/A vssd1 vssd1 vccd1 vccd1 _22533_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_156_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21306_ _21231_/X _21305_/X _21237_/X vssd1 vssd1 vccd1 vccd1 _21306_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_124_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25074_ _27179_/Q _25058_/X _25073_/X vssd1 vssd1 vccd1 vccd1 _27179_/D sky130_fd_sc_hd__o21ba_1
X_22286_ _22317_/A vssd1 vssd1 vccd1 vccd1 _22286_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24025_ _24025_/A vssd1 vssd1 vccd1 vccd1 _26884_/D sky130_fd_sc_hd__clkbuf_1
X_21237_ _21259_/A vssd1 vssd1 vccd1 vccd1 _21237_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21168_ _25927_/Q _21166_/X _21167_/X input27/X vssd1 vssd1 vccd1 vccd1 _21169_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_277_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20119_ _20119_/A _20119_/B vssd1 vssd1 vccd1 vccd1 _20125_/D sky130_fd_sc_hd__nand2_1
X_25976_ _27022_/CLK _25976_/D vssd1 vssd1 vccd1 vccd1 _25976_/Q sky130_fd_sc_hd__dfxtp_4
X_13990_ _26626_/Q _26722_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _13990_/X sky130_fd_sc_hd__mux2_1
X_21099_ _25908_/Q _21094_/X _21095_/X input38/X vssd1 vssd1 vccd1 vccd1 _21100_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_218_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12941_ _12941_/A _13569_/C vssd1 vssd1 vccd1 vccd1 _12941_/Y sky130_fd_sc_hd__nand2_1
X_24927_ _24957_/A vssd1 vssd1 vccd1 vccd1 _24927_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ _14765_/A _16122_/S _15244_/A _15659_/Y vssd1 vssd1 vccd1 vccd1 _17837_/A
+ sky130_fd_sc_hd__o22a_2
X_12872_ _12872_/A vssd1 vssd1 vccd1 vccd1 _14407_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24858_ _24856_/Y _24857_/X _24854_/X vssd1 vssd1 vccd1 vccd1 _27120_/D sky130_fd_sc_hd__a21oi_1
XFILLER_74_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _14611_/A vssd1 vssd1 vccd1 vccd1 _14612_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23809_ _23809_/A vssd1 vssd1 vccd1 vccd1 _26788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _15914_/S vssd1 vssd1 vccd1 vccd1 _16178_/S sky130_fd_sc_hd__clkbuf_4
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24789_ _24810_/A vssd1 vssd1 vccd1 vccd1 _24789_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17330_ _17327_/X _17331_/C _25530_/Q vssd1 vssd1 vccd1 vccd1 _17332_/B sky130_fd_sc_hd__a21oi_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _14542_/A _14542_/B _14542_/C vssd1 vssd1 vccd1 vccd1 _14542_/X sky130_fd_sc_hd__or3_1
X_26528_ _27303_/CLK _26528_/D vssd1 vssd1 vccd1 vccd1 _26528_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _17259_/X _17263_/C _17260_/Y vssd1 vssd1 vccd1 vccd1 _25508_/D sky130_fd_sc_hd__o21a_1
XFILLER_202_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26459_ _27267_/CLK _26459_/D vssd1 vssd1 vccd1 vccd1 _26459_/Q sky130_fd_sc_hd__dfxtp_1
X_14473_ _14471_/X _14472_/X _14473_/S vssd1 vssd1 vccd1 vccd1 _14473_/X sky130_fd_sc_hd__mux2_2
XFILLER_198_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16212_ _25653_/Q _16212_/B vssd1 vssd1 vccd1 vccd1 _16212_/X sky130_fd_sc_hd__and2_1
XFILLER_174_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19000_ _18740_/X _18997_/Y _18999_/X _18975_/Y _18777_/X vssd1 vssd1 vccd1 vccd1
+ _19000_/X sky130_fd_sc_hd__o32a_2
X_13424_ _15903_/S vssd1 vssd1 vccd1 vccd1 _15727_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17192_ _20674_/A vssd1 vssd1 vccd1 vccd1 _20630_/B sky130_fd_sc_hd__buf_2
XFILLER_155_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16143_ _26509_/Q _26381_/Q _16143_/S vssd1 vssd1 vccd1 vccd1 _16143_/X sky130_fd_sc_hd__mux2_1
X_13355_ _16004_/S vssd1 vssd1 vccd1 vccd1 _13535_/S sky130_fd_sc_hd__buf_2
XFILLER_139_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16074_ _26671_/Q _16151_/S _16073_/X _15169_/A vssd1 vssd1 vccd1 vccd1 _16074_/X
+ sky130_fd_sc_hd__o211a_1
X_13286_ _13652_/S vssd1 vssd1 vccd1 vccd1 _13675_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_182_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19902_ _20186_/A vssd1 vssd1 vccd1 vccd1 _19902_/X sky130_fd_sc_hd__clkbuf_2
X_15025_ _26870_/Q _25784_/Q _16235_/S vssd1 vssd1 vccd1 vccd1 _15025_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19833_ _19833_/A vssd1 vssd1 vccd1 vccd1 _19833_/X sky130_fd_sc_hd__buf_2
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19764_ _22480_/A _19762_/B _19763_/X vssd1 vssd1 vccd1 vccd1 _19764_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_256_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16976_ _16976_/A vssd1 vssd1 vccd1 vccd1 _16976_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_272_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18715_ _18715_/A vssd1 vssd1 vccd1 vccd1 _25609_/D sky130_fd_sc_hd__clkbuf_1
Xinput6 coreIndex[5] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15927_ _13266_/A _26857_/Q _25771_/Q _13262_/A _15924_/A vssd1 vssd1 vccd1 vccd1
+ _15927_/X sky130_fd_sc_hd__a221o_1
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19695_ _17738_/B _18377_/A _20092_/B _25575_/Q vssd1 vssd1 vccd1 vccd1 _19704_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_77_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18646_ _18548_/X _18645_/X _13553_/B vssd1 vssd1 vccd1 vccd1 _18646_/X sky130_fd_sc_hd__a21o_1
XFILLER_37_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15858_ _25811_/Q _27245_/Q _15858_/S vssd1 vssd1 vccd1 vccd1 _15859_/B sky130_fd_sc_hd__mux2_1
XFILLER_209_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14809_ _14794_/X _14797_/X _14805_/X _17181_/A vssd1 vssd1 vccd1 vccd1 _14809_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_206_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18577_ _18577_/A vssd1 vssd1 vccd1 vccd1 _19231_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_212_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15789_ _18901_/S _15789_/B vssd1 vssd1 vccd1 vccd1 _18906_/A sky130_fd_sc_hd__nor2_4
XFILLER_205_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17528_ _17548_/A _17528_/B vssd1 vssd1 vccd1 vccd1 _25566_/D sky130_fd_sc_hd__nor2_1
XFILLER_33_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17459_ _17459_/A vssd1 vssd1 vccd1 vccd1 _17460_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_220_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20470_ _20470_/A _20470_/B vssd1 vssd1 vccd1 vccd1 _20471_/C sky130_fd_sc_hd__xnor2_1
X_19129_ _25522_/Q _18556_/X _18557_/X _25554_/Q vssd1 vssd1 vccd1 vccd1 _19129_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22140_ _22179_/A vssd1 vssd1 vccd1 vccd1 _22140_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput310 _16746_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[14] sky130_fd_sc_hd__buf_2
Xoutput321 _16774_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[24] sky130_fd_sc_hd__buf_2
Xoutput332 _16733_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[9] sky130_fd_sc_hd__buf_2
Xoutput343 _16905_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[18] sky130_fd_sc_hd__buf_2
X_22071_ _26144_/Q _20923_/X _22077_/S vssd1 vssd1 vccd1 vccd1 _22072_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput354 _16971_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[28] sky130_fd_sc_hd__buf_2
XFILLER_99_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput365 _16851_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[9] sky130_fd_sc_hd__buf_2
Xoutput376 _17004_/X vssd1 vssd1 vccd1 vccd1 din0[0] sky130_fd_sc_hd__buf_2
X_21022_ _25881_/Q _20910_/X _21026_/S vssd1 vssd1 vccd1 vccd1 _21023_/A sky130_fd_sc_hd__mux2_1
Xoutput387 _17005_/X vssd1 vssd1 vccd1 vccd1 din0[1] sky130_fd_sc_hd__buf_2
XFILLER_248_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput398 _17007_/X vssd1 vssd1 vccd1 vccd1 din0[2] sky130_fd_sc_hd__buf_2
XFILLER_259_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25830_ _27265_/CLK _25830_/D vssd1 vssd1 vccd1 vccd1 _25830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25761_ _26592_/CLK _25761_/D vssd1 vssd1 vccd1 vccd1 _25761_/Q sky130_fd_sc_hd__dfxtp_1
X_22973_ _26460_/Q _22656_/X _22973_/S vssd1 vssd1 vccd1 vccd1 _22974_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24712_ _27085_/Q _24701_/X _24711_/Y _24697_/X vssd1 vssd1 vccd1 vccd1 _24713_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_21924_ _21946_/A vssd1 vssd1 vccd1 vccd1 _21933_/S sky130_fd_sc_hd__buf_4
X_25692_ _26240_/CLK _25692_/D vssd1 vssd1 vccd1 vccd1 _25692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_270_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24643_ _24768_/A _24781_/B _24639_/X _24771_/A _24701_/A vssd1 vssd1 vccd1 vccd1
+ _24643_/X sky130_fd_sc_hd__a221o_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21855_ _21855_/A vssd1 vssd1 vccd1 vccd1 _26055_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20806_ _25799_/Q vssd1 vssd1 vccd1 vccd1 _20807_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_212_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24574_ _24932_/A _24582_/B vssd1 vssd1 vccd1 vccd1 _24574_/Y sky130_fd_sc_hd__nand2_1
XFILLER_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21786_ _21786_/A vssd1 vssd1 vccd1 vccd1 _26025_/D sky130_fd_sc_hd__clkbuf_1
X_26313_ _26322_/CLK _26313_/D vssd1 vssd1 vccd1 vccd1 _26313_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_223_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23525_ _23525_/A vssd1 vssd1 vccd1 vccd1 _26688_/D sky130_fd_sc_hd__clkbuf_1
X_20737_ _20525_/X _25766_/Q _20739_/S vssd1 vssd1 vccd1 vccd1 _20738_/A sky130_fd_sc_hd__mux2_1
X_27293_ _27293_/CLK _27293_/D vssd1 vssd1 vccd1 vccd1 _27293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26244_ _26248_/CLK _26244_/D vssd1 vssd1 vccd1 vccd1 _26244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23456_ _26660_/Q _23063_/X _23458_/S vssd1 vssd1 vccd1 vccd1 _23457_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20668_ _20668_/A _20670_/B vssd1 vssd1 vccd1 vccd1 _20668_/X sky130_fd_sc_hd__or2_1
XFILLER_177_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22407_ _22394_/A _22381_/X _22383_/X _22337_/A vssd1 vssd1 vccd1 vccd1 _22407_/X
+ sky130_fd_sc_hd__o211a_1
X_26175_ _26238_/CLK _26175_/D vssd1 vssd1 vccd1 vccd1 _26175_/Q sky130_fd_sc_hd__dfxtp_1
X_23387_ _23387_/A vssd1 vssd1 vccd1 vccd1 _26629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20599_ _20599_/A vssd1 vssd1 vccd1 vccd1 _25717_/D sky130_fd_sc_hd__clkbuf_1
X_13140_ _13140_/A vssd1 vssd1 vccd1 vccd1 _13141_/A sky130_fd_sc_hd__buf_2
X_25126_ _20681_/A _25113_/X _25125_/X vssd1 vssd1 vccd1 vccd1 _25126_/Y sky130_fd_sc_hd__o21ai_1
X_22338_ _22337_/X _17078_/X _26225_/Q vssd1 vssd1 vccd1 vccd1 _22338_/X sky130_fd_sc_hd__a21o_1
XFILLER_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13071_ _13071_/A vssd1 vssd1 vccd1 vccd1 _13703_/A sky130_fd_sc_hd__buf_4
X_25057_ _27176_/Q _25030_/X _25056_/X vssd1 vssd1 vccd1 vccd1 _27176_/D sky130_fd_sc_hd__o21ba_1
X_22269_ _22269_/A vssd1 vssd1 vccd1 vccd1 _22269_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24008_ _24008_/A vssd1 vssd1 vccd1 vccd1 _26876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16830_ _16982_/B _16830_/B vssd1 vssd1 vccd1 vccd1 _16878_/B sky130_fd_sc_hd__and2_2
XFILLER_265_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13973_ _13521_/A _26594_/Q _13652_/S _26334_/Q _13244_/A vssd1 vssd1 vccd1 vccd1
+ _13973_/X sky130_fd_sc_hd__o221a_1
X_16761_ _25680_/Q vssd1 vssd1 vccd1 vccd1 _22513_/A sky130_fd_sc_hd__buf_2
XFILLER_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25959_ _26995_/CLK _25959_/D vssd1 vssd1 vccd1 vccd1 _25959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18500_ _18544_/A _18497_/X _18499_/X vssd1 vssd1 vccd1 vccd1 _18500_/Y sky130_fd_sc_hd__o21ai_1
X_15712_ _25613_/Q _14595_/A _15711_/Y _12977_/A vssd1 vssd1 vccd1 vccd1 _15750_/A
+ sky130_fd_sc_hd__o22a_2
X_12924_ _13748_/A vssd1 vssd1 vccd1 vccd1 _13928_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16692_ _25662_/Q vssd1 vssd1 vccd1 vccd1 _22474_/A sky130_fd_sc_hd__clkbuf_4
X_19480_ _20249_/A _18720_/X _18788_/X _19479_/Y vssd1 vssd1 vccd1 vccd1 _19480_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_262_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18431_ _18421_/Y _18425_/X _18430_/Y _18375_/X vssd1 vssd1 vccd1 vccd1 _18431_/X
+ sky130_fd_sc_hd__o31a_1
X_12855_ input131/X input166/X _25868_/Q vssd1 vssd1 vccd1 vccd1 _17653_/C sky130_fd_sc_hd__mux2_8
XFILLER_34_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15643_ _26636_/Q _26732_/Q _15643_/S vssd1 vssd1 vccd1 vccd1 _15643_/X sky130_fd_sc_hd__mux2_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15574_ _26669_/Q _25709_/Q _16087_/S vssd1 vssd1 vccd1 vccd1 _15574_/X sky130_fd_sc_hd__mux2_1
X_18362_ _18362_/A vssd1 vssd1 vccd1 vccd1 _18362_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12786_ _25688_/Q _16685_/B _14580_/C vssd1 vssd1 vccd1 vccd1 _16635_/A sky130_fd_sc_hd__nor3_4
XFILLER_15_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _17332_/A _17313_/B _17314_/B vssd1 vssd1 vccd1 vccd1 _25524_/D sky130_fd_sc_hd__nor3_1
XFILLER_202_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _16809_/B _16809_/C _16578_/B vssd1 vssd1 vccd1 vccd1 _14525_/X sky130_fd_sc_hd__a21o_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18293_ _18293_/A vssd1 vssd1 vccd1 vccd1 _18817_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14456_ _27296_/Q _26553_/Q _14472_/S vssd1 vssd1 vccd1 vccd1 _14456_/X sky130_fd_sc_hd__mux2_1
X_17244_ _24208_/A vssd1 vssd1 vccd1 vccd1 _24966_/A sky130_fd_sc_hd__buf_2
XFILLER_179_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13407_ _14349_/S vssd1 vssd1 vccd1 vccd1 _14178_/S sky130_fd_sc_hd__clkbuf_2
X_17175_ _22377_/A vssd1 vssd1 vccd1 vccd1 _17175_/X sky130_fd_sc_hd__clkbuf_2
X_14387_ _14535_/A _14387_/B _14387_/C vssd1 vssd1 vccd1 vccd1 _14387_/X sky130_fd_sc_hd__or3_1
XFILLER_190_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16126_ _19045_/B vssd1 vssd1 vccd1 vccd1 _19048_/A sky130_fd_sc_hd__inv_2
X_13338_ _13475_/A vssd1 vssd1 vccd1 vccd1 _13339_/A sky130_fd_sc_hd__buf_2
XFILLER_143_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16057_ _26347_/Q _26607_/Q _16078_/S vssd1 vssd1 vccd1 vccd1 _16057_/X sky130_fd_sc_hd__mux2_1
X_13269_ _13269_/A vssd1 vssd1 vccd1 vccd1 _17658_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_29_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15008_ _14804_/A _15004_/X _15007_/X _14818_/X vssd1 vssd1 vccd1 vccd1 _15008_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19816_ _19814_/Y _19816_/B vssd1 vssd1 vccd1 vccd1 _19819_/A sky130_fd_sc_hd__and2b_1
XFILLER_284_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_257_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19747_ _24848_/A vssd1 vssd1 vccd1 vccd1 _20712_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_284_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16959_ _16980_/A _16959_/B _16959_/C vssd1 vssd1 vccd1 vccd1 _16960_/A sky130_fd_sc_hd__and3_2
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19678_ _19657_/X _19674_/Y _19675_/X _19677_/Y vssd1 vssd1 vccd1 vccd1 _19678_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_237_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18629_ _13685_/X _18285_/A _18628_/X _18409_/X _25607_/Q vssd1 vssd1 vccd1 vccd1
+ _18630_/B sky130_fd_sc_hd__a32o_1
XFILLER_213_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21640_ _25499_/Q vssd1 vssd1 vccd1 vccd1 _21641_/A sky130_fd_sc_hd__inv_2
XFILLER_75_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21571_ _21565_/Y _21570_/X _21556_/X vssd1 vssd1 vccd1 vccd1 _21571_/Y sky130_fd_sc_hd__a21oi_4
X_23310_ _23310_/A vssd1 vssd1 vccd1 vccd1 _26595_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20522_ _20521_/X _25699_/Q _20530_/S vssd1 vssd1 vccd1 vccd1 _20523_/A sky130_fd_sc_hd__mux2_1
X_24290_ _26987_/Q _24293_/C _24289_/Y vssd1 vssd1 vccd1 vccd1 _26987_/D sky130_fd_sc_hd__o21a_1
XFILLER_192_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23241_ _23241_/A vssd1 vssd1 vccd1 vccd1 _26564_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20453_ _19740_/X _20442_/Y _20452_/X _19765_/X vssd1 vssd1 vccd1 vccd1 _20453_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_119_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23172_ _26534_/Q _23082_/X _23172_/S vssd1 vssd1 vccd1 vccd1 _23173_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20384_ _19657_/X _20420_/C _20383_/Y _20100_/X vssd1 vssd1 vccd1 vccd1 _20385_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_284_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22123_ _22210_/A _22206_/A vssd1 vssd1 vccd1 vccd1 _22179_/A sky130_fd_sc_hd__and2_2
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22054_ _22054_/A vssd1 vssd1 vccd1 vccd1 _26136_/D sky130_fd_sc_hd__clkbuf_1
X_26931_ _26931_/CLK _26931_/D vssd1 vssd1 vccd1 vccd1 _26931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21005_ _21005_/A vssd1 vssd1 vccd1 vccd1 _25873_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26862_ _27311_/CLK _26862_/D vssd1 vssd1 vccd1 vccd1 _26862_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25813_ _26917_/CLK _25813_/D vssd1 vssd1 vccd1 vccd1 _25813_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26793_ _26827_/CLK _26793_/D vssd1 vssd1 vccd1 vccd1 _26793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25744_ _26282_/CLK _25744_/D vssd1 vssd1 vccd1 vccd1 _25744_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22956_ _26453_/Q _22736_/X _22956_/S vssd1 vssd1 vccd1 vccd1 _22957_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21907_ _20521_/X _26071_/Q _21911_/S vssd1 vssd1 vccd1 vccd1 _21908_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25675_ _27122_/CLK _25675_/D vssd1 vssd1 vccd1 vccd1 _25675_/Q sky130_fd_sc_hd__dfxtp_1
X_22887_ _22887_/A vssd1 vssd1 vccd1 vccd1 _26422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24626_ _27066_/Q _24615_/X _24625_/Y _24619_/X vssd1 vssd1 vccd1 vccd1 _27066_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_243_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21838_ _26048_/Q _20932_/X _21838_/S vssd1 vssd1 vccd1 vccd1 _21839_/A sky130_fd_sc_hd__mux2_1
XFILLER_270_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24557_ _24915_/A _24569_/B vssd1 vssd1 vccd1 vccd1 _24557_/Y sky130_fd_sc_hd__nand2_1
XFILLER_157_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21769_ _21769_/A vssd1 vssd1 vccd1 vccd1 _26017_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14310_ _26491_/Q _26363_/Q _14310_/S vssd1 vssd1 vccd1 vccd1 _14310_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23508_ _23508_/A vssd1 vssd1 vccd1 vccd1 _23508_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_169_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27276_ _27276_/CLK _27276_/D vssd1 vssd1 vccd1 vccd1 _27276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15290_ _15290_/A _16927_/A vssd1 vssd1 vccd1 vccd1 _15290_/Y sky130_fd_sc_hd__nor2_1
XFILLER_183_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24488_ _24492_/A _24605_/A vssd1 vssd1 vccd1 vccd1 _24488_/Y sky130_fd_sc_hd__nand2_1
XFILLER_157_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26227_ _27297_/CLK _26227_/D vssd1 vssd1 vccd1 vccd1 _26227_/Q sky130_fd_sc_hd__dfxtp_1
X_14241_ _13911_/X _14489_/A _14240_/X _12916_/X _25905_/Q vssd1 vssd1 vccd1 vccd1
+ _14241_/X sky130_fd_sc_hd__o32a_1
X_23439_ _26652_/Q _23034_/X _23447_/S vssd1 vssd1 vccd1 vccd1 _23440_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14172_ _26848_/Q _25762_/Q _15714_/A vssd1 vssd1 vccd1 vccd1 _14172_/X sky130_fd_sc_hd__mux2_1
X_26158_ _26938_/CLK _26158_/D vssd1 vssd1 vccd1 vccd1 _26158_/Q sky130_fd_sc_hd__dfxtp_1
X_13123_ _14111_/A vssd1 vssd1 vccd1 vccd1 _13124_/A sky130_fd_sc_hd__clkbuf_2
X_25109_ _25109_/A vssd1 vssd1 vccd1 vccd1 _25109_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18980_ _18683_/A _18858_/X _18859_/Y _18682_/X vssd1 vssd1 vccd1 vccd1 _18980_/X
+ sky130_fd_sc_hd__o211a_1
X_26089_ _26677_/CLK _26089_/D vssd1 vssd1 vccd1 vccd1 _26089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _14348_/S vssd1 vssd1 vccd1 vccd1 _14344_/S sky130_fd_sc_hd__clkbuf_2
X_17931_ _18050_/S vssd1 vssd1 vccd1 vccd1 _18265_/S sky130_fd_sc_hd__clkbuf_2
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17862_ _18899_/A vssd1 vssd1 vccd1 vccd1 _19358_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19601_ _25573_/Q _19600_/X _18027_/A _17697_/B vssd1 vssd1 vccd1 vccd1 _19659_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_78_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16813_ _16833_/A _16813_/B _16813_/C vssd1 vssd1 vccd1 vccd1 _16848_/B sky130_fd_sc_hd__and3_4
XFILLER_213_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17793_ _17793_/A _15342_/B vssd1 vssd1 vccd1 vccd1 _17793_/X sky130_fd_sc_hd__or2b_1
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19532_ _25647_/Q _19536_/B vssd1 vssd1 vccd1 vccd1 _19532_/X sky130_fd_sc_hd__or2_1
XFILLER_4_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16744_ _22498_/A _16742_/X _16743_/X _16635_/C vssd1 vssd1 vccd1 vccd1 _16744_/X
+ sky130_fd_sc_hd__a22o_1
X_13956_ _16006_/A vssd1 vssd1 vccd1 vccd1 _15760_/A sky130_fd_sc_hd__buf_4
XFILLER_219_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12907_ _21429_/A _12878_/B _12873_/A vssd1 vssd1 vccd1 vccd1 _12907_/Y sky130_fd_sc_hd__o21ai_1
X_19463_ _27100_/Q _18751_/X _18752_/X _27198_/Q _18753_/X vssd1 vssd1 vccd1 vccd1
+ _19463_/X sky130_fd_sc_hd__a221o_1
X_13887_ _26659_/Q _15734_/S _13886_/X _15716_/S vssd1 vssd1 vccd1 vccd1 _13887_/X
+ sky130_fd_sc_hd__o211a_1
X_16675_ _20977_/A _16668_/B vssd1 vssd1 vccd1 vccd1 _16679_/B sky130_fd_sc_hd__nor2b_4
XFILLER_235_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18414_ _18209_/X _18206_/X _18416_/S vssd1 vssd1 vccd1 vccd1 _18414_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12838_ _25861_/Q vssd1 vssd1 vccd1 vccd1 _16657_/A sky130_fd_sc_hd__clkbuf_4
X_15626_ _26860_/Q _25774_/Q _16143_/S vssd1 vssd1 vccd1 vccd1 _15626_/X sky130_fd_sc_hd__mux2_1
XFILLER_261_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19394_ _16556_/A _18548_/X _19392_/Y _16794_/B _19393_/Y vssd1 vssd1 vccd1 vccd1
+ _19394_/X sky130_fd_sc_hd__o221a_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18345_ _18053_/X _18043_/X _18345_/S vssd1 vssd1 vccd1 vccd1 _18345_/X sky130_fd_sc_hd__mux2_1
X_12769_ _12769_/A vssd1 vssd1 vccd1 vccd1 _12770_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15557_ _26637_/Q _26733_/Q _15557_/S vssd1 vssd1 vccd1 vccd1 _15557_/X sky130_fd_sc_hd__mux2_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_168_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26292_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14508_ _15979_/S _14503_/X _14504_/X _14507_/X _13162_/A vssd1 vssd1 vccd1 vccd1
+ _14508_/X sky130_fd_sc_hd__o311a_1
X_15488_ _15488_/A vssd1 vssd1 vccd1 vccd1 _15488_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18276_ _16707_/B _17997_/A _18275_/X _16713_/A vssd1 vssd1 vccd1 vccd1 _18276_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_175_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17227_ _20487_/B vssd1 vssd1 vccd1 vccd1 _25176_/A sky130_fd_sc_hd__buf_4
Xinput20 core_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_1
X_14439_ _13029_/A _14435_/Y _14438_/X _14331_/X vssd1 vssd1 vccd1 vccd1 _14439_/X
+ sky130_fd_sc_hd__o2bb2a_1
Xinput31 core_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
XFILLER_175_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput42 core_wb_error_i vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_1
Xinput53 dout0[19] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput64 dout0[29] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput75 dout0[39] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__clkbuf_1
X_17158_ _17158_/A vssd1 vssd1 vccd1 vccd1 _25479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput86 dout0[49] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput97 dout0[59] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16109_ _27314_/Q _26571_/Q _16178_/S vssd1 vssd1 vccd1 vccd1 _16109_/X sky130_fd_sc_hd__mux2_1
X_17089_ _26236_/Q _26233_/Q _26232_/Q _17085_/A vssd1 vssd1 vccd1 vccd1 _17089_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_89_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22810_ _22810_/A vssd1 vssd1 vccd1 vccd1 _26388_/D sky130_fd_sc_hd__clkbuf_1
X_23790_ _23858_/S vssd1 vssd1 vccd1 vccd1 _23799_/S sky130_fd_sc_hd__buf_4
XFILLER_272_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22741_ _22741_/A vssd1 vssd1 vccd1 vccd1 _26358_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25460_ _25460_/A vssd1 vssd1 vccd1 vccd1 _27324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_279_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22672_ _23715_/A vssd1 vssd1 vccd1 vccd1 _22672_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_241_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24411_ _26301_/Q _24382_/X _24383_/X input245/X _24384_/X vssd1 vssd1 vccd1 vccd1
+ _24411_/X sky130_fd_sc_hd__a221o_1
X_21623_ _20699_/A _21278_/A _21563_/A _21622_/X vssd1 vssd1 vccd1 vccd1 _21623_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_178_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25391_ _27294_/Q _23785_/A _25391_/S vssd1 vssd1 vccd1 vccd1 _25392_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27130_ _27130_/CLK _27130_/D vssd1 vssd1 vccd1 vccd1 _27130_/Q sky130_fd_sc_hd__dfxtp_2
X_24342_ _24342_/A vssd1 vssd1 vccd1 vccd1 _24342_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21554_ _21554_/A vssd1 vssd1 vccd1 vccd1 _21554_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20505_ _20504_/X _25695_/Q _20509_/S vssd1 vssd1 vccd1 vccd1 _20506_/A sky130_fd_sc_hd__mux2_1
X_27061_ _27062_/CLK _27061_/D vssd1 vssd1 vccd1 vccd1 _27061_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_154_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24273_ _26981_/Q _24275_/C _24272_/Y vssd1 vssd1 vccd1 vccd1 _26981_/D sky130_fd_sc_hd__o21a_1
XFILLER_165_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21485_ _21482_/X _21484_/X _21433_/X vssd1 vssd1 vccd1 vccd1 _21485_/X sky130_fd_sc_hd__a21o_1
X_26012_ _26531_/CLK _26012_/D vssd1 vssd1 vccd1 vccd1 _26012_/Q sky130_fd_sc_hd__dfxtp_1
X_23224_ _23281_/S vssd1 vssd1 vccd1 vccd1 _23233_/S sky130_fd_sc_hd__buf_4
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20436_ _20433_/X _20434_/Y _20435_/Y vssd1 vssd1 vccd1 vccd1 _20436_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_181_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23155_ _26526_/Q _23057_/X _23161_/S vssd1 vssd1 vccd1 vccd1 _23156_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20367_ _27159_/Q _27093_/Q vssd1 vssd1 vccd1 vccd1 _20367_/Y sky130_fd_sc_hd__nor2_1
X_22106_ _22393_/A _26237_/Q _22395_/A vssd1 vssd1 vccd1 vccd1 _22236_/C sky130_fd_sc_hd__and3_1
XFILLER_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23086_ _23118_/A vssd1 vssd1 vccd1 vccd1 _23099_/S sky130_fd_sc_hd__buf_4
X_20298_ _22520_/A _20225_/X _20290_/X _20297_/X _20223_/X vssd1 vssd1 vccd1 vccd1
+ _25683_/D sky130_fd_sc_hd__o221a_1
XTAP_5602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22037_ _22037_/A vssd1 vssd1 vccd1 vccd1 _26128_/D sky130_fd_sc_hd__clkbuf_1
X_26914_ _26917_/CLK _26914_/D vssd1 vssd1 vccd1 vccd1 _26914_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26845_ _26845_/CLK _26845_/D vssd1 vssd1 vccd1 vccd1 _26845_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ _26495_/Q _26367_/Q _16014_/S vssd1 vssd1 vccd1 vccd1 _13811_/B sky130_fd_sc_hd__mux2_1
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14790_ _16281_/S vssd1 vssd1 vccd1 vccd1 _14790_/X sky130_fd_sc_hd__clkbuf_4
X_23988_ _23988_/A vssd1 vssd1 vccd1 vccd1 _26868_/D sky130_fd_sc_hd__clkbuf_1
X_26776_ _27259_/CLK _26776_/D vssd1 vssd1 vccd1 vccd1 _26776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_263_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13741_ input114/X input149/X _13741_/S vssd1 vssd1 vccd1 vccd1 _13742_/B sky130_fd_sc_hd__mux2_8
XFILLER_272_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25727_ _26264_/CLK _25727_/D vssd1 vssd1 vccd1 vccd1 _25727_/Q sky130_fd_sc_hd__dfxtp_4
X_22939_ _26445_/Q _22711_/X _22945_/S vssd1 vssd1 vccd1 vccd1 _22940_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13672_ _26661_/Q _25701_/Q _15842_/S vssd1 vssd1 vccd1 vccd1 _13672_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16460_ _16560_/A _16562_/A _19393_/A _16561_/B vssd1 vssd1 vccd1 vccd1 _16461_/B
+ sky130_fd_sc_hd__a211o_1
X_25658_ _26248_/CLK _25658_/D vssd1 vssd1 vccd1 vccd1 _25658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15411_ _15406_/X _27283_/Q _26476_/Q _16440_/S _15318_/A vssd1 vssd1 vccd1 vccd1
+ _15411_/X sky130_fd_sc_hd__a221o_1
X_24609_ _27059_/Q _24602_/X _24608_/Y _24606_/X vssd1 vssd1 vccd1 vccd1 _27059_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16391_ _14650_/A _16386_/X _16390_/X _14679_/X vssd1 vssd1 vccd1 vccd1 _16391_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25589_ _26684_/CLK _25589_/D vssd1 vssd1 vccd1 vccd1 _25589_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18130_ _25534_/Q _18568_/A _18127_/X _19069_/A _18572_/A vssd1 vssd1 vccd1 vccd1
+ _18130_/X sky130_fd_sc_hd__a221o_1
XFILLER_197_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15342_ _17793_/A _15342_/B vssd1 vssd1 vccd1 vccd1 _15343_/B sky130_fd_sc_hd__nor2_1
XPHY_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18061_ _18061_/A vssd1 vssd1 vccd1 vccd1 _18061_/Y sky130_fd_sc_hd__inv_2
X_15273_ _15065_/A _26898_/Q _26770_/Q _16399_/S _15169_/X vssd1 vssd1 vccd1 vccd1
+ _15273_/X sky130_fd_sc_hd__a221o_1
XFILLER_185_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27259_ _27259_/CLK _27259_/D vssd1 vssd1 vccd1 vccd1 _27259_/Q sky130_fd_sc_hd__dfxtp_1
X_14224_ _26492_/Q _26364_/Q _16014_/S vssd1 vssd1 vccd1 vccd1 _14224_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17012_ _16810_/A _17008_/X _16878_/B _17006_/X input243/X vssd1 vssd1 vccd1 vccd1
+ _17012_/X sky130_fd_sc_hd__a32o_4
XFILLER_172_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14155_ _13889_/A _14152_/X _14154_/X vssd1 vssd1 vccd1 vccd1 _14156_/B sky130_fd_sc_hd__o21ai_1
XFILLER_256_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13106_ _14100_/A vssd1 vssd1 vccd1 vccd1 _13107_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14086_ _26525_/Q _26133_/Q _14095_/A vssd1 vssd1 vccd1 vccd1 _14086_/X sky130_fd_sc_hd__mux2_1
X_18963_ _25740_/Q _18964_/B vssd1 vssd1 vccd1 vccd1 _19037_/C sky130_fd_sc_hd__and2_1
X_13037_ _15453_/A vssd1 vssd1 vccd1 vccd1 _15561_/B sky130_fd_sc_hd__buf_2
X_17914_ _17941_/A vssd1 vssd1 vccd1 vccd1 _18318_/S sky130_fd_sc_hd__clkbuf_2
X_18894_ _18964_/B _18894_/B vssd1 vssd1 vccd1 vccd1 _18894_/X sky130_fd_sc_hd__or2_2
XFILLER_121_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17845_ _19109_/B _19109_/C _17844_/X _16289_/A _19156_/A vssd1 vssd1 vccd1 vccd1
+ _19237_/C sky130_fd_sc_hd__a2111o_1
XFILLER_78_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17776_ _17776_/A vssd1 vssd1 vccd1 vccd1 _18339_/A sky130_fd_sc_hd__buf_2
XFILLER_35_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14988_ _26680_/Q _25720_/Q _14991_/S vssd1 vssd1 vccd1 vccd1 _14988_/X sky130_fd_sc_hd__mux2_1
XFILLER_242_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19515_ _19541_/A vssd1 vssd1 vccd1 vccd1 _19515_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_235_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16727_ _16770_/A vssd1 vssd1 vccd1 vccd1 _16727_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13939_ _13939_/A vssd1 vssd1 vccd1 vccd1 _13939_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_208_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_510 _17066_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_521 _17023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19446_ _18895_/X _19430_/X _19445_/X _18927_/X vssd1 vssd1 vccd1 vccd1 _19446_/X
+ sky130_fd_sc_hd__a22o_1
XINSDIODE2_532 _17049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_543 _25727_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16658_ _16660_/A _20796_/B vssd1 vssd1 vccd1 vccd1 _20990_/B sky130_fd_sc_hd__nand2_8
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_554 _25728_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15609_ _15606_/X _15607_/X _15608_/X _13367_/A vssd1 vssd1 vccd1 vccd1 _15610_/B
+ sky130_fd_sc_hd__a31o_1
X_19377_ _19234_/A _19375_/Y _19376_/X _19385_/B _18839_/X vssd1 vssd1 vccd1 vccd1
+ _19377_/X sky130_fd_sc_hd__o32a_1
XFILLER_250_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16589_ _16853_/A _16589_/B vssd1 vssd1 vccd1 vccd1 _16782_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18328_ _18328_/A _18328_/B vssd1 vssd1 vccd1 vccd1 _18328_/X sky130_fd_sc_hd__or2_1
XFILLER_249_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18259_ _18257_/X _18258_/X _18348_/S vssd1 vssd1 vccd1 vccd1 _18259_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21270_ input65/X input70/X _21356_/S vssd1 vssd1 vccd1 vccd1 _21271_/B sky130_fd_sc_hd__mux2_8
XFILLER_144_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20221_ _19991_/X _20220_/X _20052_/X vssd1 vssd1 vccd1 vccd1 _20221_/Y sky130_fd_sc_hd__o21ai_1
X_20152_ _25677_/Q _20151_/C _22509_/A vssd1 vssd1 vccd1 vccd1 _20152_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_277_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_65_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27272_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_24960_ _24960_/A _24972_/B vssd1 vssd1 vccd1 vccd1 _24960_/Y sky130_fd_sc_hd__nand2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20083_ _20084_/A _20084_/B vssd1 vssd1 vccd1 vccd1 _20083_/X sky130_fd_sc_hd__or2_1
XFILLER_281_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23911_ _23757_/X _26834_/Q _23915_/S vssd1 vssd1 vccd1 vccd1 _23912_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24891_ _20699_/A _19963_/X _25159_/A _24779_/A vssd1 vssd1 vccd1 vccd1 _24891_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_258_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26630_ _27309_/CLK _26630_/D vssd1 vssd1 vccd1 vccd1 _26630_/Q sky130_fd_sc_hd__dfxtp_1
X_23842_ _23842_/A vssd1 vssd1 vccd1 vccd1 _26803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26561_ _27303_/CLK _26561_/D vssd1 vssd1 vccd1 vccd1 _26561_/Q sky130_fd_sc_hd__dfxtp_1
X_23773_ _23773_/A vssd1 vssd1 vccd1 vccd1 _23773_/X sky130_fd_sc_hd__buf_2
X_20985_ _20985_/A vssd1 vssd1 vccd1 vccd1 _25864_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25512_ _27014_/CLK _25512_/D vssd1 vssd1 vccd1 vccd1 _25512_/Q sky130_fd_sc_hd__dfxtp_1
X_22724_ _22724_/A vssd1 vssd1 vccd1 vccd1 _22737_/S sky130_fd_sc_hd__buf_4
X_26492_ _26657_/CLK _26492_/D vssd1 vssd1 vccd1 vccd1 _26492_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_225_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25443_ _25443_/A vssd1 vssd1 vccd1 vccd1 _27316_/D sky130_fd_sc_hd__clkbuf_1
X_22655_ _22655_/A vssd1 vssd1 vccd1 vccd1 _26331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21606_ _21606_/A vssd1 vssd1 vccd1 vccd1 _21606_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25374_ _27286_/Q _23760_/A _25376_/S vssd1 vssd1 vccd1 vccd1 _25375_/A sky130_fd_sc_hd__mux2_1
X_22586_ _26310_/Q _22591_/B vssd1 vssd1 vccd1 vccd1 _22586_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24325_ _26999_/Q _24326_/C _27000_/Q vssd1 vssd1 vccd1 vccd1 _24327_/B sky130_fd_sc_hd__a21oi_1
X_27113_ _27196_/CLK _27113_/D vssd1 vssd1 vccd1 vccd1 _27113_/Q sky130_fd_sc_hd__dfxtp_4
X_21537_ _21603_/A vssd1 vssd1 vccd1 vccd1 _21537_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27044_ _27044_/CLK _27044_/D vssd1 vssd1 vccd1 vccd1 _27044_/Q sky130_fd_sc_hd__dfxtp_1
X_24256_ _26975_/Q _24258_/C _24255_/Y vssd1 vssd1 vccd1 vccd1 _26975_/D sky130_fd_sc_hd__o21a_1
X_21468_ _25952_/Q _21443_/X _21466_/Y _21467_/X vssd1 vssd1 vccd1 vccd1 _25952_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_181_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23207_ _26550_/Q _23133_/X _23209_/S vssd1 vssd1 vccd1 vccd1 _23208_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20419_ _25689_/Q vssd1 vssd1 vccd1 vccd1 _22531_/A sky130_fd_sc_hd__buf_2
X_24187_ _26953_/Q _24191_/C vssd1 vssd1 vccd1 vccd1 _24188_/B sky130_fd_sc_hd__and2_1
XFILLER_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21399_ _24208_/A vssd1 vssd1 vccd1 vccd1 _21597_/A sky130_fd_sc_hd__buf_8
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23138_ _23138_/A vssd1 vssd1 vccd1 vccd1 _26519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_268_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23069_ _23542_/A vssd1 vssd1 vccd1 vccd1 _23069_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15960_ _27307_/Q _26564_/Q _15964_/S vssd1 vssd1 vccd1 vccd1 _15960_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput210 localMemory_wb_adr_i[6] vssd1 vssd1 vccd1 vccd1 input210/X sky130_fd_sc_hd__clkbuf_1
XTAP_5432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput221 localMemory_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input221/X sky130_fd_sc_hd__buf_6
XFILLER_68_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput232 localMemory_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 input232/X sky130_fd_sc_hd__buf_8
XFILLER_264_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14911_ _14779_/A _14907_/X _14910_/X _14787_/X vssd1 vssd1 vccd1 vccd1 _14911_/Y
+ sky130_fd_sc_hd__o31ai_2
XTAP_5454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput243 localMemory_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input243/X sky130_fd_sc_hd__buf_6
Xinput254 manufacturerID[10] vssd1 vssd1 vccd1 vccd1 input254/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15891_ _13585_/A _26697_/Q _26825_/Q _15726_/S _13049_/A vssd1 vssd1 vccd1 vccd1
+ _15891_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput265 partID[10] vssd1 vssd1 vccd1 vccd1 input265/X sky130_fd_sc_hd__clkbuf_1
XTAP_5476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput276 partID[6] vssd1 vssd1 vccd1 vccd1 input276/X sky130_fd_sc_hd__clkbuf_1
X_17630_ _17633_/A _17630_/B vssd1 vssd1 vccd1 vccd1 _25589_/D sky130_fd_sc_hd__nor2_1
XFILLER_84_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ _16396_/S vssd1 vssd1 vccd1 vccd1 _16384_/S sky130_fd_sc_hd__clkbuf_4
X_26828_ _27314_/CLK _26828_/D vssd1 vssd1 vccd1 vccd1 _26828_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17561_ _17560_/X _12846_/X _17544_/X _25909_/Q vssd1 vssd1 vccd1 vccd1 _17561_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_90_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26759_ _26889_/CLK _26759_/D vssd1 vssd1 vccd1 vccd1 _26759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14773_ _14773_/A vssd1 vssd1 vccd1 vccd1 _14773_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_216_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19300_ _27095_/Q _18815_/X _18816_/X _27193_/Q _18817_/X vssd1 vssd1 vccd1 vccd1
+ _19300_/X sky130_fd_sc_hd__a221o_1
XFILLER_216_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16512_ _26651_/Q _26747_/Q _16523_/S vssd1 vssd1 vccd1 vccd1 _16512_/X sky130_fd_sc_hd__mux2_1
X_13724_ _26496_/Q _26368_/Q _16067_/S vssd1 vssd1 vccd1 vccd1 _13724_/X sky130_fd_sc_hd__mux2_1
X_17492_ _17683_/A _21218_/C vssd1 vssd1 vccd1 vccd1 _21219_/B sky130_fd_sc_hd__nand2_1
XFILLER_182_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19231_ _19231_/A _19231_/B vssd1 vssd1 vccd1 vccd1 _19231_/Y sky130_fd_sc_hd__nor2_1
X_16443_ _26679_/Q _25719_/Q _16443_/S vssd1 vssd1 vccd1 vccd1 _16443_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13655_ _25806_/Q _27240_/Q _14221_/S vssd1 vssd1 vccd1 vccd1 _13655_/X sky130_fd_sc_hd__mux2_1
XFILLER_231_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19162_ _17308_/X _18807_/X _18808_/X _25555_/Q vssd1 vssd1 vccd1 vccd1 _19162_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13586_ _26337_/Q _15807_/S vssd1 vssd1 vccd1 vccd1 _13586_/X sky130_fd_sc_hd__or2_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16374_ _19273_/A _19240_/S _16370_/A vssd1 vssd1 vccd1 vccd1 _16374_/X sky130_fd_sc_hd__o21a_1
XFILLER_83_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18113_ _27134_/Q _18454_/A _18103_/A vssd1 vssd1 vccd1 vccd1 _18113_/X sky130_fd_sc_hd__a21bo_1
X_15325_ _15313_/X _15320_/X _15324_/X _14792_/A vssd1 vssd1 vccd1 vccd1 _15325_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_118_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19093_ _27153_/Q _19367_/B vssd1 vssd1 vccd1 vccd1 _19093_/X sky130_fd_sc_hd__or2_1
XFILLER_8_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18044_ _17891_/X _17881_/X _18044_/S vssd1 vssd1 vccd1 vccd1 _18044_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15256_ _16315_/S vssd1 vssd1 vccd1 vccd1 _16301_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_173_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14207_ _13941_/X _14205_/X _14206_/X _13945_/X vssd1 vssd1 vccd1 vccd1 _14211_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_160_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15187_ _15187_/A vssd1 vssd1 vccd1 vccd1 _15187_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_141_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14138_ _15874_/A _14138_/B vssd1 vssd1 vccd1 vccd1 _14138_/Y sky130_fd_sc_hd__nand2_1
XFILLER_259_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19995_ _27145_/Q _27079_/Q vssd1 vssd1 vccd1 vccd1 _19999_/B sky130_fd_sc_hd__nor2_1
X_14069_ _25582_/Q _14069_/B _14069_/C vssd1 vssd1 vccd1 vccd1 _14077_/B sky130_fd_sc_hd__or3_1
XFILLER_86_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18946_ _18946_/A _19231_/B vssd1 vssd1 vccd1 vccd1 _18947_/B sky130_fd_sc_hd__nor2_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18877_ _19140_/A vssd1 vssd1 vccd1 vccd1 _19442_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17828_ _17828_/A _16035_/B vssd1 vssd1 vccd1 vccd1 _18794_/A sky130_fd_sc_hd__or2b_1
XFILLER_95_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17759_ _18454_/A vssd1 vssd1 vccd1 vccd1 _18821_/A sky130_fd_sc_hd__buf_2
XFILLER_282_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_183_wb_clk_i _26681_/CLK vssd1 vssd1 vccd1 vccd1 _27324_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_251_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20770_ _20588_/X _25781_/Q _20772_/S vssd1 vssd1 vccd1 vccd1 _20771_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_340 _19609_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_112_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26980_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XINSDIODE2_351 _19612_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_362 input231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19429_ _18602_/X _18075_/Y _18084_/X _18342_/A _19428_/X vssd1 vssd1 vccd1 vccd1
+ _19429_/X sky130_fd_sc_hd__o221a_1
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_373 _16992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_384 _17004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_395 _17034_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22440_ _26249_/Q _22444_/B vssd1 vssd1 vccd1 vccd1 _22440_/X sky130_fd_sc_hd__or2_1
XFILLER_148_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22371_ _25466_/A _22371_/B vssd1 vssd1 vccd1 vccd1 _22372_/A sky130_fd_sc_hd__or2_1
XFILLER_109_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24110_ _24110_/A vssd1 vssd1 vccd1 vccd1 _26922_/D sky130_fd_sc_hd__clkbuf_1
X_21322_ _21547_/A vssd1 vssd1 vccd1 vccd1 _21322_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_276_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25090_ _24707_/Y _25070_/X _25089_/Y _25082_/X vssd1 vssd1 vccd1 vccd1 _25090_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_190_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24041_ _24041_/A vssd1 vssd1 vccd1 vccd1 _26891_/D sky130_fd_sc_hd__clkbuf_1
X_21253_ _21289_/A vssd1 vssd1 vccd1 vccd1 _21589_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20204_ _20204_/A _20204_/B _20200_/Y vssd1 vssd1 vccd1 vccd1 _20301_/A sky130_fd_sc_hd__or3b_1
XFILLER_278_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21184_ _25932_/Q _21112_/A _21113_/A input33/X vssd1 vssd1 vccd1 vccd1 _21185_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_131_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20135_ _20135_/A _20135_/B vssd1 vssd1 vccd1 vccd1 _20135_/Y sky130_fd_sc_hd__xnor2_1
X_25992_ _25992_/CLK _25992_/D vssd1 vssd1 vccd1 vccd1 _25992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24943_ _27146_/Q _24927_/X _24942_/Y vssd1 vssd1 vccd1 vccd1 _27146_/D sky130_fd_sc_hd__o21a_1
X_20066_ _22502_/A _20098_/C _20065_/Y vssd1 vssd1 vccd1 vccd1 _20067_/C sky130_fd_sc_hd__a21oi_1
XFILLER_100_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_11 _18694_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_22 _19103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_33 _19315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_44 _20630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_55 _20643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24874_ _24874_/A vssd1 vssd1 vccd1 vccd1 _24896_/B sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_66 _20654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_77 _20699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_88 _21878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26613_ _27324_/CLK _26613_/D vssd1 vssd1 vccd1 vccd1 _26613_/Q sky130_fd_sc_hd__dfxtp_1
X_23825_ _23825_/A vssd1 vssd1 vccd1 vccd1 _26795_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_99 _21464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26544_ _26739_/CLK _26544_/D vssd1 vssd1 vccd1 vccd1 _26544_/Q sky130_fd_sc_hd__dfxtp_1
X_23756_ _23756_/A vssd1 vssd1 vccd1 vccd1 _26769_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20968_ _25859_/Q _20967_/X _20971_/S vssd1 vssd1 vccd1 vccd1 _20969_/A sky130_fd_sc_hd__mux2_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22707_ _23750_/A vssd1 vssd1 vccd1 vccd1 _22707_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23687_ _23786_/S vssd1 vssd1 vccd1 vccd1 _23700_/S sky130_fd_sc_hd__buf_4
X_26475_ _26796_/CLK _26475_/D vssd1 vssd1 vccd1 vccd1 _26475_/Q sky130_fd_sc_hd__dfxtp_1
X_20899_ _20899_/A vssd1 vssd1 vccd1 vccd1 _25837_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13440_ _15825_/S vssd1 vssd1 vccd1 vccd1 _13441_/S sky130_fd_sc_hd__clkbuf_4
X_22638_ _22638_/A _22638_/B _22638_/C _22638_/D vssd1 vssd1 vccd1 vccd1 _22639_/A
+ sky130_fd_sc_hd__and4_1
X_25426_ _23731_/X _27309_/Q _25426_/S vssd1 vssd1 vccd1 vccd1 _25427_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25357_ _27278_/Q _23734_/A _25365_/S vssd1 vssd1 vccd1 vccd1 _25358_/A sky130_fd_sc_hd__mux2_1
X_13371_ _13276_/Y _13315_/Y _13370_/Y _13314_/X _14789_/A vssd1 vssd1 vccd1 vccd1
+ _13371_/Y sky130_fd_sc_hd__o221ai_4
X_22569_ _26303_/Q _22578_/B vssd1 vssd1 vccd1 vccd1 _22569_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15110_ _15110_/A vssd1 vssd1 vccd1 vccd1 _15111_/A sky130_fd_sc_hd__buf_2
X_24308_ _26993_/Q _24309_/C _26994_/Q vssd1 vssd1 vccd1 vccd1 _24310_/B sky130_fd_sc_hd__a21oi_1
XFILLER_194_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16090_ _13267_/X _26703_/Q _26831_/Q _16186_/S _16088_/A vssd1 vssd1 vccd1 vccd1
+ _16090_/X sky130_fd_sc_hd__a221o_1
X_25288_ _25288_/A vssd1 vssd1 vccd1 vccd1 _27247_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15041_ _15060_/S _15036_/X _15038_/X _15040_/X vssd1 vssd1 vccd1 vccd1 _15041_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_108_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24239_ _24239_/A vssd1 vssd1 vccd1 vccd1 _24269_/A sky130_fd_sc_hd__buf_2
X_27027_ _27058_/CLK _27027_/D vssd1 vssd1 vccd1 vccd1 _27027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18800_ _18859_/A _18798_/X _18799_/Y _18321_/A vssd1 vssd1 vccd1 vccd1 _18803_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_268_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19780_ _20015_/A vssd1 vssd1 vccd1 vccd1 _19780_/X sky130_fd_sc_hd__buf_2
X_16992_ _22476_/A _16988_/X _16990_/X _18230_/B vssd1 vssd1 vccd1 vccd1 _16992_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_95_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18731_ _18859_/A _18273_/Y _18730_/X vssd1 vssd1 vccd1 vccd1 _18731_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_62_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15943_ _15205_/A _15941_/X _15942_/X _13366_/A vssd1 vssd1 vccd1 vccd1 _15943_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_62_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18662_ _17268_/X _18444_/X _18659_/X _18661_/X _18469_/X vssd1 vssd1 vccd1 vccd1
+ _18662_/X sky130_fd_sc_hd__o221a_1
XTAP_5295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _15874_/A _15874_/B _15874_/C vssd1 vssd1 vccd1 vccd1 _15874_/X sky130_fd_sc_hd__and3_1
XFILLER_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17613_ _25922_/Q _17597_/X _14133_/Y _17518_/X vssd1 vssd1 vccd1 vccd1 _17613_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ _18028_/A _12738_/X _14806_/A vssd1 vssd1 vccd1 vccd1 _14826_/A sky130_fd_sc_hd__o21a_1
XFILLER_28_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18593_ _18593_/A _18593_/B _18593_/C vssd1 vssd1 vccd1 vccd1 _18594_/B sky130_fd_sc_hd__nor3_1
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17544_ _17554_/A vssd1 vssd1 vccd1 vccd1 _17544_/X sky130_fd_sc_hd__buf_2
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14756_ _16513_/A _25859_/Q _26059_/Q _14767_/S _14755_/X vssd1 vssd1 vccd1 vccd1
+ _14756_/X sky130_fd_sc_hd__a221o_1
XFILLER_205_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13707_ _15734_/S vssd1 vssd1 vccd1 vccd1 _15464_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17475_ _21208_/A _21214_/A _17475_/C _21208_/B vssd1 vssd1 vccd1 vccd1 _17475_/X
+ sky130_fd_sc_hd__or4b_1
X_14687_ _15048_/A vssd1 vssd1 vccd1 vccd1 _14688_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_220_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19214_ _18976_/X _19212_/X _20279_/A _19003_/X vssd1 vssd1 vccd1 vccd1 _19214_/X
+ sky130_fd_sc_hd__a22o_2
X_16426_ _26935_/Q _26419_/Q _16440_/S vssd1 vssd1 vccd1 vccd1 _16426_/X sky130_fd_sc_hd__mux2_1
X_13638_ _13638_/A vssd1 vssd1 vccd1 vccd1 _13638_/X sky130_fd_sc_hd__buf_6
XFILLER_146_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19145_ _18716_/X _19128_/X _19144_/X _19078_/X vssd1 vssd1 vccd1 vccd1 _19145_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16357_ _14753_/A _16354_/X _16356_/X _14792_/A vssd1 vssd1 vccd1 vccd1 _16357_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_173_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13569_ _13569_/A _13569_/B _13569_/C vssd1 vssd1 vccd1 vccd1 _13570_/A sky130_fd_sc_hd__and3_1
X_15308_ _15306_/X _15307_/X _15308_/S vssd1 vssd1 vccd1 vccd1 _15308_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19076_ _19076_/A vssd1 vssd1 vccd1 vccd1 _19076_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16288_ _16288_/A _16288_/B vssd1 vssd1 vccd1 vccd1 _16289_/A sky130_fd_sc_hd__nor2_1
XFILLER_173_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18027_ _18027_/A vssd1 vssd1 vccd1 vccd1 _18027_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15239_ _17782_/A _17781_/A vssd1 vssd1 vccd1 vccd1 _15240_/B sky130_fd_sc_hd__and2_1
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19978_ _19978_/A _19978_/B vssd1 vssd1 vccd1 vccd1 _19978_/X sky130_fd_sc_hd__and2_1
XFILLER_99_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18929_ _19087_/A vssd1 vssd1 vccd1 vccd1 _18929_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_268_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21940_ _20584_/X _26086_/Q _21944_/S vssd1 vssd1 vccd1 vccd1 _21941_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21871_ _24456_/A vssd1 vssd1 vccd1 vccd1 _21871_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_215_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23610_ _26715_/Q _23609_/X _23610_/S vssd1 vssd1 vccd1 vccd1 _23611_/A sky130_fd_sc_hd__mux2_1
XFILLER_270_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20822_ _25807_/Q vssd1 vssd1 vccd1 vccd1 _20823_/A sky130_fd_sc_hd__clkbuf_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24590_ _24590_/A _24595_/B vssd1 vssd1 vccd1 vccd1 _24590_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23541_ _23541_/A vssd1 vssd1 vccd1 vccd1 _26693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20753_ _20554_/X _25773_/Q _20761_/S vssd1 vssd1 vccd1 vccd1 _20754_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_170 _14449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_181 _19849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26260_ _26974_/CLK _26260_/D vssd1 vssd1 vccd1 vccd1 _26260_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_192 _15902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23472_ _26667_/Q _23085_/X _23480_/S vssd1 vssd1 vccd1 vccd1 _23473_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20684_ _21878_/A vssd1 vssd1 vccd1 vccd1 _20684_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25211_ _27215_/Q _25204_/X _25207_/X _24711_/B _25210_/X vssd1 vssd1 vccd1 vccd1
+ _27215_/D sky130_fd_sc_hd__o221a_1
XFILLER_10_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22423_ _26242_/Q _22430_/B vssd1 vssd1 vccd1 vccd1 _22423_/X sky130_fd_sc_hd__or2_1
X_26191_ _26238_/CLK _26191_/D vssd1 vssd1 vccd1 vccd1 _26191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25142_ _25142_/A vssd1 vssd1 vccd1 vccd1 _25151_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_22354_ _22356_/A _26231_/Q _17235_/X _22353_/Y vssd1 vssd1 vccd1 vccd1 _26230_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_136_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27238_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21305_ input87/X input72/X _21327_/S vssd1 vssd1 vccd1 vccd1 _21305_/X sky130_fd_sc_hd__mux2_8
XFILLER_237_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25073_ _24693_/Y _25070_/X _25072_/Y _25055_/X vssd1 vssd1 vccd1 vccd1 _25073_/X
+ sky130_fd_sc_hd__a31o_1
X_22285_ _22630_/B vssd1 vssd1 vccd1 vccd1 _22285_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24024_ _26884_/Q _23536_/X _24026_/S vssd1 vssd1 vccd1 vccd1 _24025_/A sky130_fd_sc_hd__mux2_1
X_21236_ _21581_/A vssd1 vssd1 vccd1 vccd1 _21259_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21167_ _21167_/A vssd1 vssd1 vccd1 vccd1 _21167_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20118_ _20118_/A _20118_/B vssd1 vssd1 vccd1 vccd1 _20127_/A sky130_fd_sc_hd__or2_1
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25975_ _27058_/CLK _25975_/D vssd1 vssd1 vccd1 vccd1 _25975_/Q sky130_fd_sc_hd__dfxtp_4
X_21098_ _21098_/A vssd1 vssd1 vccd1 vccd1 _25907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12940_ _14407_/A _14025_/B _13559_/B _12940_/D vssd1 vssd1 vccd1 vccd1 _14239_/A
+ sky130_fd_sc_hd__or4_2
X_24926_ _19839_/A _24902_/X _24925_/Y vssd1 vssd1 vccd1 vccd1 _27140_/D sky130_fd_sc_hd__o21a_1
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20049_ _20022_/Y _20024_/Y _20046_/X _20047_/Y vssd1 vssd1 vccd1 vccd1 _20049_/Y
+ sky130_fd_sc_hd__a211oi_2
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _12871_/A vssd1 vssd1 vccd1 vccd1 _12871_/Y sky130_fd_sc_hd__inv_2
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24857_ _20675_/A _24848_/X _24725_/Y _24849_/X vssd1 vssd1 vccd1 vccd1 _24857_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _14610_/A _14610_/B vssd1 vssd1 vccd1 vccd1 _14611_/A sky130_fd_sc_hd__nand2_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23808_ _23712_/X _26788_/Q _23810_/S vssd1 vssd1 vccd1 vccd1 _23809_/A sky130_fd_sc_hd__mux2_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _15676_/A _26345_/Q _26605_/Q _16194_/S _15670_/A vssd1 vssd1 vccd1 vccd1
+ _15590_/X sky130_fd_sc_hd__a221o_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24788_ _27103_/Q _24798_/B vssd1 vssd1 vccd1 vccd1 _24788_/Y sky130_fd_sc_hd__nand2_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26527_ _27272_/CLK _26527_/D vssd1 vssd1 vccd1 vccd1 _26527_/Q sky130_fd_sc_hd__dfxtp_1
X_14541_ _13941_/A _14539_/X _14540_/X _13939_/A vssd1 vssd1 vccd1 vccd1 _14542_/C
+ sky130_fd_sc_hd__o211a_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23739_ _23738_/X _26764_/Q _23748_/S vssd1 vssd1 vccd1 vccd1 _23740_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _17259_/X _17263_/C _17235_/X vssd1 vssd1 vccd1 vccd1 _17260_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_197_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26458_ _27266_/CLK _26458_/D vssd1 vssd1 vccd1 vccd1 _26458_/Q sky130_fd_sc_hd__dfxtp_2
X_14472_ _26097_/Q _25998_/Q _14472_/S vssd1 vssd1 vccd1 vccd1 _14472_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16211_ _15245_/X _15704_/Y _14604_/A vssd1 vssd1 vccd1 vccd1 _16211_/Y sky130_fd_sc_hd__a21oi_1
X_13423_ _14115_/S vssd1 vssd1 vccd1 vccd1 _15903_/S sky130_fd_sc_hd__buf_6
X_25409_ _23706_/X _27301_/Q _25415_/S vssd1 vssd1 vccd1 vccd1 _25410_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17191_ _25465_/S vssd1 vssd1 vccd1 vccd1 _20674_/A sky130_fd_sc_hd__buf_4
X_26389_ _27292_/CLK _26389_/D vssd1 vssd1 vccd1 vccd1 _26389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13354_ _14310_/S vssd1 vssd1 vccd1 vccd1 _16004_/S sky130_fd_sc_hd__clkbuf_2
X_16142_ _26349_/Q _26609_/Q _16143_/S vssd1 vssd1 vccd1 vccd1 _16142_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13285_ _14536_/S vssd1 vssd1 vccd1 vccd1 _13652_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_154_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16073_ _25711_/Q _16073_/B vssd1 vssd1 vccd1 vccd1 _16073_/X sky130_fd_sc_hd__or2_1
XFILLER_142_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15024_ _15030_/S vssd1 vssd1 vccd1 vccd1 _16235_/S sky130_fd_sc_hd__buf_2
X_19901_ _19899_/Y _19900_/X _19896_/A _20323_/B vssd1 vssd1 vccd1 vccd1 _19901_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19832_ _19766_/X _19830_/Y _19831_/X _19780_/X vssd1 vssd1 vccd1 vccd1 _19837_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_69_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19763_ _20452_/A vssd1 vssd1 vccd1 vccd1 _19763_/X sky130_fd_sc_hd__buf_2
X_16975_ _16980_/A _16975_/B _16975_/C vssd1 vssd1 vccd1 vccd1 _16976_/A sky130_fd_sc_hd__and3_2
XFILLER_7_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18714_ _22368_/A _18714_/B vssd1 vssd1 vccd1 vccd1 _18715_/A sky130_fd_sc_hd__and2_1
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15926_ _13266_/A _26921_/Q _26405_/Q _13262_/A _15916_/A vssd1 vssd1 vccd1 vccd1
+ _15926_/X sky130_fd_sc_hd__a221o_1
XFILLER_265_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19694_ _19879_/A vssd1 vssd1 vccd1 vccd1 _19766_/A sky130_fd_sc_hd__clkbuf_2
Xinput7 coreIndex[6] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_283_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18645_ _18686_/B _19192_/B _18645_/S vssd1 vssd1 vccd1 vccd1 _18645_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15857_ _27309_/Q _26566_/Q _15857_/S vssd1 vssd1 vccd1 vccd1 _15857_/X sky130_fd_sc_hd__mux2_1
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14808_ _14808_/A vssd1 vssd1 vccd1 vccd1 _17181_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18576_ _18555_/X _18558_/X _18575_/X vssd1 vssd1 vccd1 vccd1 _18576_/X sky130_fd_sc_hd__a21o_4
XFILLER_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15788_ _17826_/A _15788_/B vssd1 vssd1 vccd1 vccd1 _15789_/B sky130_fd_sc_hd__nor2_1
XFILLER_45_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17527_ _25566_/Q _20686_/A _17516_/X _17526_/X vssd1 vssd1 vccd1 vccd1 _17528_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14739_ _14811_/S vssd1 vssd1 vccd1 vccd1 _16510_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_205_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17458_ _21244_/A _17458_/B vssd1 vssd1 vccd1 vccd1 _17459_/A sky130_fd_sc_hd__nor2_1
XFILLER_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16409_ _16409_/A _16409_/B vssd1 vssd1 vccd1 vccd1 _16409_/Y sky130_fd_sc_hd__nor2_1
X_17389_ _25547_/Q _25548_/Q _17389_/C vssd1 vssd1 vccd1 vccd1 _17392_/B sky130_fd_sc_hd__and3_1
XFILLER_118_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19128_ _18636_/X _19124_/X _19127_/X vssd1 vssd1 vccd1 vccd1 _19128_/X sky130_fd_sc_hd__a21o_1
XFILLER_257_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19059_ _19059_/A vssd1 vssd1 vccd1 vccd1 _19059_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput300 _16998_/X vssd1 vssd1 vccd1 vccd1 addr1[6] sky130_fd_sc_hd__buf_2
XFILLER_146_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput311 _16749_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[15] sky130_fd_sc_hd__buf_2
Xoutput322 _16777_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[25] sky130_fd_sc_hd__buf_2
X_22070_ _22070_/A vssd1 vssd1 vccd1 vccd1 _26143_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput333 _21195_/A vssd1 vssd1 vccd1 vccd1 core_wb_cyc_o sky130_fd_sc_hd__buf_2
XFILLER_160_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput344 _16915_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[19] sky130_fd_sc_hd__buf_2
Xoutput355 _16976_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[29] sky130_fd_sc_hd__buf_2
X_21021_ _21021_/A vssd1 vssd1 vccd1 vccd1 _25880_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput366 _16786_/X vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[0] sky130_fd_sc_hd__buf_2
XFILLER_99_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput377 _17022_/X vssd1 vssd1 vccd1 vccd1 din0[10] sky130_fd_sc_hd__buf_2
Xoutput388 _17036_/X vssd1 vssd1 vccd1 vccd1 din0[20] sky130_fd_sc_hd__buf_2
Xoutput399 _17048_/X vssd1 vssd1 vccd1 vccd1 din0[30] sky130_fd_sc_hd__buf_2
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22972_ _22972_/A vssd1 vssd1 vccd1 vccd1 _26459_/D sky130_fd_sc_hd__clkbuf_1
X_25760_ _26909_/CLK _25760_/D vssd1 vssd1 vccd1 vccd1 _25760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24711_ _24725_/A _24711_/B vssd1 vssd1 vccd1 vccd1 _24711_/Y sky130_fd_sc_hd__nand2_2
XFILLER_283_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21923_ _21923_/A vssd1 vssd1 vccd1 vccd1 _26078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25691_ _27132_/CLK _25691_/D vssd1 vssd1 vccd1 vccd1 _25691_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_215_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21854_ _26055_/Q _20955_/X _21860_/S vssd1 vssd1 vccd1 vccd1 _21855_/A sky130_fd_sc_hd__mux2_1
X_24642_ _24744_/A vssd1 vssd1 vccd1 vccd1 _24701_/A sky130_fd_sc_hd__buf_2
XFILLER_222_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20805_ _20805_/A vssd1 vssd1 vccd1 vccd1 _25798_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_24573_ _27045_/Q _24562_/X _24572_/Y _24567_/X vssd1 vssd1 vccd1 vccd1 _27045_/D
+ sky130_fd_sc_hd__o211a_1
X_21785_ _20609_/X _26025_/Q _21787_/S vssd1 vssd1 vccd1 vccd1 _21786_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26312_ _26322_/CLK _26312_/D vssd1 vssd1 vccd1 vccd1 _26312_/Q sky130_fd_sc_hd__dfxtp_2
X_20736_ _20736_/A vssd1 vssd1 vccd1 vccd1 _25765_/D sky130_fd_sc_hd__clkbuf_1
X_23524_ _26688_/Q _23523_/X _23524_/S vssd1 vssd1 vccd1 vccd1 _23525_/A sky130_fd_sc_hd__mux2_1
X_27292_ _27292_/CLK _27292_/D vssd1 vssd1 vccd1 vccd1 _27292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26243_ _26248_/CLK _26243_/D vssd1 vssd1 vccd1 vccd1 _26243_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_195_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23455_ _23455_/A vssd1 vssd1 vccd1 vccd1 _26659_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20667_ _26277_/Q _20660_/X _20666_/X _20658_/X vssd1 vssd1 vccd1 vccd1 _25740_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_196_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22406_ _22406_/A _22406_/B vssd1 vssd1 vccd1 vccd1 _22406_/X sky130_fd_sc_hd__or2_1
XFILLER_13_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26174_ _26238_/CLK _26174_/D vssd1 vssd1 vccd1 vccd1 _26174_/Q sky130_fd_sc_hd__dfxtp_1
X_23386_ _26629_/Q _23066_/X _23386_/S vssd1 vssd1 vccd1 vccd1 _23387_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20598_ _20596_/X _25717_/Q _20614_/S vssd1 vssd1 vccd1 vccd1 _20599_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22337_ _22337_/A vssd1 vssd1 vccd1 vccd1 _22337_/X sky130_fd_sc_hd__buf_2
X_25125_ _22518_/A _25119_/X _25114_/X _16638_/A _25106_/X vssd1 vssd1 vccd1 vccd1
+ _25125_/X sky130_fd_sc_hd__a221o_1
XFILLER_137_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13070_ _13998_/S vssd1 vssd1 vccd1 vccd1 _13071_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25056_ _24682_/Y _25043_/X _25054_/Y _25055_/X vssd1 vssd1 vccd1 vccd1 _25056_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_279_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22268_ _26202_/Q _22254_/X _22267_/X _22258_/X vssd1 vssd1 vccd1 vccd1 _26202_/D
+ sky130_fd_sc_hd__o211a_1
X_24007_ _26876_/Q _23508_/X _24015_/S vssd1 vssd1 vccd1 vccd1 _24008_/A sky130_fd_sc_hd__mux2_1
X_21219_ _21219_/A _21219_/B _21221_/B _21208_/D vssd1 vssd1 vccd1 vccd1 _21251_/A
+ sky130_fd_sc_hd__nor4b_1
XFILLER_3_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22199_ _26184_/Q _22185_/X _22198_/X _22195_/X vssd1 vssd1 vccd1 vccd1 _26184_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_278_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16760_ _22511_/A _16756_/X _16757_/X _19046_/A vssd1 vssd1 vccd1 vccd1 _16760_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_281_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25958_ _26995_/CLK _25958_/D vssd1 vssd1 vccd1 vccd1 _25958_/Q sky130_fd_sc_hd__dfxtp_1
X_13972_ _26494_/Q _26366_/Q _14369_/S vssd1 vssd1 vccd1 vccd1 _13972_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15711_ _13558_/A _15709_/X _15710_/Y vssd1 vssd1 vccd1 vccd1 _15711_/Y sky130_fd_sc_hd__a21oi_1
X_24909_ _24938_/A vssd1 vssd1 vccd1 vccd1 _24909_/X sky130_fd_sc_hd__clkbuf_2
X_12923_ _25795_/Q vssd1 vssd1 vccd1 vccd1 _13748_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16691_ _16691_/A vssd1 vssd1 vccd1 vccd1 _16691_/X sky130_fd_sc_hd__clkbuf_1
X_25889_ _26609_/CLK _25889_/D vssd1 vssd1 vccd1 vccd1 _25889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18430_ _18544_/A _18427_/X _18429_/X vssd1 vssd1 vccd1 vccd1 _18430_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_262_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15642_ _15640_/X _15641_/X _16079_/S vssd1 vssd1 vccd1 vccd1 _15642_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _16657_/A _25793_/Q vssd1 vssd1 vccd1 vccd1 _12893_/A sky130_fd_sc_hd__nand2_2
XFILLER_73_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _19454_/A vssd1 vssd1 vccd1 vccd1 _18544_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _16439_/A _16122_/S _15244_/A _15572_/Y vssd1 vssd1 vccd1 vccd1 _17838_/A
+ sky130_fd_sc_hd__o22a_4
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _25687_/Q _25686_/Q _25685_/Q _25684_/Q vssd1 vssd1 vccd1 vccd1 _14580_/C
+ sky130_fd_sc_hd__or4_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _25523_/Q _25524_/Q _17312_/C vssd1 vssd1 vccd1 vccd1 _17314_/B sky130_fd_sc_hd__and3_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14524_ _13172_/A _14509_/X _14523_/X _13026_/A vssd1 vssd1 vccd1 vccd1 _16809_/C
+ sky130_fd_sc_hd__o31a_4
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18292_ _18292_/A vssd1 vssd1 vccd1 vccd1 _18816_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17243_ _17283_/A _17243_/B _17243_/C vssd1 vssd1 vccd1 vccd1 _25503_/D sky130_fd_sc_hd__nor3_1
X_14455_ _13337_/A _14452_/X _14454_/X _13827_/A vssd1 vssd1 vccd1 vccd1 _14455_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_174_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13406_ _27305_/Q _26562_/Q _13719_/A vssd1 vssd1 vccd1 vccd1 _13406_/X sky130_fd_sc_hd__mux2_1
X_17174_ _25484_/Q _17185_/B vssd1 vssd1 vccd1 vccd1 _17174_/X sky130_fd_sc_hd__or2_1
X_14386_ _14064_/X _14383_/X _14385_/X _13309_/B vssd1 vssd1 vccd1 vccd1 _14387_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16125_ _16125_/A _16124_/Y vssd1 vssd1 vccd1 vccd1 _19045_/B sky130_fd_sc_hd__nor2b_2
X_13337_ _13337_/A vssd1 vssd1 vccd1 vccd1 _13475_/A sky130_fd_sc_hd__buf_2
XFILLER_143_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16056_ _15384_/S _16053_/X _16055_/X _14659_/A vssd1 vssd1 vccd1 vccd1 _16056_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_170_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13268_ _13267_/X _26887_/Q _26759_/Q _16341_/S _13221_/A vssd1 vssd1 vccd1 vccd1
+ _13268_/X sky130_fd_sc_hd__a221o_1
XFILLER_29_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15007_ _14755_/A _15005_/X _15006_/X _14794_/A vssd1 vssd1 vccd1 vccd1 _15007_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_269_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13199_ _14043_/A vssd1 vssd1 vccd1 vccd1 _13336_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_269_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19815_ _27139_/Q _27073_/Q vssd1 vssd1 vccd1 vccd1 _19816_/B sky130_fd_sc_hd__nand2_1
XFILLER_285_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19746_ _27105_/Q _19722_/X _19724_/X _19745_/Y vssd1 vssd1 vccd1 vccd1 _19746_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16958_ _16855_/Y _16954_/X _16956_/X _16852_/X _16957_/Y vssd1 vssd1 vccd1 vccd1
+ _16959_/C sky130_fd_sc_hd__a221o_1
XFILLER_272_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15909_ _13876_/X _15885_/X _15893_/X _15908_/X vssd1 vssd1 vccd1 vccd1 _15909_/X
+ sky130_fd_sc_hd__a31o_2
X_19677_ _25662_/Q _19833_/A _20100_/A vssd1 vssd1 vccd1 vccd1 _19677_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_65_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16889_ _16889_/A _16927_/B vssd1 vssd1 vccd1 vccd1 _16889_/X sky130_fd_sc_hd__or2_2
XFILLER_253_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18628_ _19256_/A _16732_/X _18627_/X vssd1 vssd1 vccd1 vccd1 _18628_/X sky130_fd_sc_hd__a21bo_1
XFILLER_53_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18559_ _18559_/A vssd1 vssd1 vccd1 vccd1 _18559_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_252_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_19_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27314_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_178_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21570_ _21552_/X _21566_/X _21569_/Y _21518_/X vssd1 vssd1 vccd1 vccd1 _21570_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_177_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20521_ _23709_/A vssd1 vssd1 vccd1 vccd1 _20521_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23240_ _26564_/Q _23076_/X _23244_/S vssd1 vssd1 vccd1 vccd1 _23241_/A sky130_fd_sc_hd__mux2_1
X_20452_ _20452_/A _20452_/B _20471_/B vssd1 vssd1 vccd1 vccd1 _20452_/X sky130_fd_sc_hd__or3b_1
XFILLER_174_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23171_ _23171_/A vssd1 vssd1 vccd1 vccd1 _26533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20383_ _25686_/Q _20382_/C _22528_/A vssd1 vssd1 vccd1 vccd1 _20383_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_173_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22122_ _22122_/A vssd1 vssd1 vccd1 vccd1 _22122_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_284_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22053_ _26136_/Q _20897_/X _22055_/S vssd1 vssd1 vccd1 vccd1 _22054_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26930_ _27253_/CLK _26930_/D vssd1 vssd1 vccd1 vccd1 _26930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21004_ _25873_/Q _20884_/X _21004_/S vssd1 vssd1 vccd1 vccd1 _21005_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26861_ _26925_/CLK _26861_/D vssd1 vssd1 vccd1 vccd1 _26861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25812_ _27293_/CLK _25812_/D vssd1 vssd1 vccd1 vccd1 _25812_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26792_ _26920_/CLK _26792_/D vssd1 vssd1 vccd1 vccd1 _26792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25743_ _26282_/CLK _25743_/D vssd1 vssd1 vccd1 vccd1 _25743_/Q sky130_fd_sc_hd__dfxtp_4
X_22955_ _22955_/A vssd1 vssd1 vccd1 vccd1 _26452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21906_ _21906_/A vssd1 vssd1 vccd1 vccd1 _26070_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25674_ _27122_/CLK _25674_/D vssd1 vssd1 vccd1 vccd1 _25674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22886_ _26422_/Q _22739_/X _22888_/S vssd1 vssd1 vccd1 vccd1 _22887_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24625_ _24625_/A _24629_/B vssd1 vssd1 vccd1 vccd1 _24625_/Y sky130_fd_sc_hd__nand2_1
X_21837_ _21837_/A vssd1 vssd1 vccd1 vccd1 _26047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24556_ _24610_/A vssd1 vssd1 vccd1 vccd1 _24569_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_178_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21768_ _20575_/X _26017_/Q _21776_/S vssd1 vssd1 vccd1 vccd1 _21769_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20719_ _20787_/S vssd1 vssd1 vccd1 vccd1 _20728_/S sky130_fd_sc_hd__buf_2
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23507_ _23507_/A vssd1 vssd1 vccd1 vccd1 _26683_/D sky130_fd_sc_hd__clkbuf_1
X_27275_ _27275_/CLK _27275_/D vssd1 vssd1 vccd1 vccd1 _27275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21699_ _25988_/Q input200/X _21707_/S vssd1 vssd1 vccd1 vccd1 _21700_/A sky130_fd_sc_hd__mux2_1
X_24487_ _24732_/B vssd1 vssd1 vccd1 vccd1 _24605_/A sky130_fd_sc_hd__clkinv_2
XFILLER_200_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26226_ _27297_/CLK _26226_/D vssd1 vssd1 vccd1 vccd1 _26226_/Q sky130_fd_sc_hd__dfxtp_1
X_14240_ input140/X input135/X _14240_/S vssd1 vssd1 vccd1 vccd1 _14240_/X sky130_fd_sc_hd__mux2_8
X_23438_ _23506_/S vssd1 vssd1 vccd1 vccd1 _23447_/S sky130_fd_sc_hd__buf_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14171_ _14107_/X _14168_/X _14170_/X _14111_/X vssd1 vssd1 vccd1 vccd1 _14171_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_165_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23369_ _26621_/Q _23041_/X _23375_/S vssd1 vssd1 vccd1 vccd1 _23370_/A sky130_fd_sc_hd__mux2_1
X_26157_ _26453_/CLK _26157_/D vssd1 vssd1 vccd1 vccd1 _26157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13122_ _14331_/A vssd1 vssd1 vccd1 vccd1 _14111_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_164_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25108_ _20675_/A _25086_/X _25107_/X vssd1 vssd1 vccd1 vccd1 _25108_/Y sky130_fd_sc_hd__o21ai_1
X_26088_ _27287_/CLK _26088_/D vssd1 vssd1 vccd1 vccd1 _26088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13053_ _26791_/Q _26435_/Q _15566_/S vssd1 vssd1 vccd1 vccd1 _13053_/X sky130_fd_sc_hd__mux2_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17930_ _17928_/X _17929_/X _18042_/S vssd1 vssd1 vccd1 vccd1 _17930_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25039_ _25666_/Q _25038_/X _25033_/X _18424_/A _25024_/X vssd1 vssd1 vccd1 vccd1
+ _25039_/X sky130_fd_sc_hd__a221o_1
XFILLER_79_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17861_ _18597_/A vssd1 vssd1 vccd1 vccd1 _18899_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19600_ _19670_/A vssd1 vssd1 vccd1 vccd1 _19600_/X sky130_fd_sc_hd__buf_2
X_16812_ _16812_/A vssd1 vssd1 vccd1 vccd1 _16828_/A sky130_fd_sc_hd__clkbuf_1
X_17792_ _19121_/B _19122_/A _17791_/X vssd1 vssd1 vccd1 vccd1 _17792_/X sky130_fd_sc_hd__o21a_1
XFILLER_266_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19531_ _19525_/X _18958_/X _19530_/X _19528_/X vssd1 vssd1 vccd1 vccd1 _25646_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16743_ _16770_/A vssd1 vssd1 vccd1 vccd1 _16743_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13955_ _13955_/A vssd1 vssd1 vccd1 vccd1 _16006_/A sky130_fd_sc_hd__buf_2
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12906_ _15954_/B vssd1 vssd1 vccd1 vccd1 _14604_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_19462_ _27230_/Q _19462_/B vssd1 vssd1 vccd1 vccd1 _19462_/X sky130_fd_sc_hd__and2_1
X_16674_ _16674_/A vssd1 vssd1 vccd1 vccd1 _20978_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_34_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13886_ _25699_/Q _15808_/B vssd1 vssd1 vccd1 vccd1 _13886_/X sky130_fd_sc_hd__or2_1
XFILLER_35_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18413_ _18413_/A vssd1 vssd1 vccd1 vccd1 _18413_/Y sky130_fd_sc_hd__inv_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15625_ _15265_/X _15622_/X _15624_/X _15019_/A vssd1 vssd1 vccd1 vccd1 _15625_/X
+ sky130_fd_sc_hd__a211o_1
X_12837_ _12837_/A vssd1 vssd1 vccd1 vccd1 _12891_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19393_ _19393_/A _19393_/B vssd1 vssd1 vccd1 vccd1 _19393_/Y sky130_fd_sc_hd__nand2_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18344_ _18344_/A vssd1 vssd1 vccd1 vccd1 _18344_/Y sky130_fd_sc_hd__inv_2
X_15556_ _15554_/X _15555_/X _15567_/S vssd1 vssd1 vccd1 vccd1 _15556_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _12768_/A vssd1 vssd1 vccd1 vccd1 _12769_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14111_/X _14505_/X _14506_/X _13409_/A vssd1 vssd1 vccd1 vccd1 _14507_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_202_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18275_ _16707_/B _18603_/A _18214_/A vssd1 vssd1 vccd1 vccd1 _18275_/X sky130_fd_sc_hd__o21a_1
X_15487_ _13359_/X _15484_/X _15486_/X _15312_/A vssd1 vssd1 vccd1 vccd1 _15495_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_202_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12699_ _13630_/A vssd1 vssd1 vccd1 vccd1 _12700_/A sky130_fd_sc_hd__buf_2
X_17226_ _25501_/Q vssd1 vssd1 vccd1 vccd1 _17242_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14438_ _14436_/X _14437_/X _14515_/S vssd1 vssd1 vccd1 vccd1 _14438_/X sky130_fd_sc_hd__mux2_1
Xinput10 core_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput21 core_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_1
Xinput32 core_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
Xinput43 dout0[0] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_2
Xinput54 dout0[1] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_2
X_17157_ _17200_/A _17157_/B vssd1 vssd1 vccd1 vccd1 _17158_/A sky130_fd_sc_hd__and2_1
X_14369_ _26490_/Q _26362_/Q _14369_/S vssd1 vssd1 vccd1 vccd1 _14369_/X sky130_fd_sc_hd__mux2_1
Xinput65 dout0[2] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput76 dout0[3] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__clkbuf_2
Xinput87 dout0[4] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_137_wb_clk_i _25501_/CLK vssd1 vssd1 vccd1 vccd1 _27044_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput98 dout0[5] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_2
X_16108_ _14729_/A _16106_/X _16107_/X _14820_/A vssd1 vssd1 vccd1 vccd1 _16108_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17088_ _26192_/Q _22230_/B _22416_/B vssd1 vssd1 vccd1 vccd1 _17088_/X sky130_fd_sc_hd__a21o_1
XFILLER_6_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16039_ _18838_/A _18838_/B _18801_/S vssd1 vssd1 vccd1 vccd1 _18851_/B sky130_fd_sc_hd__a21boi_4
XFILLER_103_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19729_ _20252_/B _18288_/Y _19671_/A _19728_/X vssd1 vssd1 vccd1 vccd1 _19729_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_226_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22740_ _26358_/Q _22739_/X _22743_/S vssd1 vssd1 vccd1 vccd1 _22741_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22671_ _22671_/A vssd1 vssd1 vccd1 vccd1 _26336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24410_ _24494_/A vssd1 vssd1 vccd1 vccd1 _24434_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_21622_ _21620_/X _21621_/X _21589_/X vssd1 vssd1 vccd1 vccd1 _21622_/X sky130_fd_sc_hd__a21o_1
XFILLER_178_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25390_ _25390_/A vssd1 vssd1 vccd1 vccd1 _27293_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21553_ input58/X input93/X _21553_/S vssd1 vssd1 vccd1 vccd1 _21554_/A sky130_fd_sc_hd__mux2_8
X_24341_ _24341_/A _24900_/C vssd1 vssd1 vccd1 vccd1 _25206_/B sky130_fd_sc_hd__or2_1
XFILLER_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20504_ _23696_/A vssd1 vssd1 vccd1 vccd1 _20504_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_24272_ _26981_/Q _24275_/C _24271_/X vssd1 vssd1 vccd1 vccd1 _24272_/Y sky130_fd_sc_hd__a21oi_1
X_27060_ _27062_/CLK _27060_/D vssd1 vssd1 vccd1 vccd1 _27060_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_138_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21484_ _21430_/X _19030_/X _21431_/X _25815_/Q _21483_/X vssd1 vssd1 vccd1 vccd1
+ _21484_/X sky130_fd_sc_hd__a221o_1
XFILLER_148_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26011_ _26599_/CLK _26011_/D vssd1 vssd1 vccd1 vccd1 _26011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23223_ _23223_/A vssd1 vssd1 vccd1 vccd1 _26556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20435_ _20413_/A _20415_/B _20412_/Y vssd1 vssd1 vccd1 vccd1 _20435_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23154_ _23154_/A vssd1 vssd1 vccd1 vccd1 _26525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20366_ _20343_/A _20342_/B _20342_/A vssd1 vssd1 vccd1 vccd1 _20370_/A sky130_fd_sc_hd__a21boi_1
X_22105_ _26240_/Q _26239_/Q vssd1 vssd1 vccd1 vccd1 _22395_/A sky130_fd_sc_hd__nor2_1
X_23085_ _23558_/A vssd1 vssd1 vccd1 vccd1 _23085_/X sky130_fd_sc_hd__clkbuf_2
X_20297_ _20179_/X _20296_/X _20186_/X vssd1 vssd1 vccd1 vccd1 _20297_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22036_ _26128_/Q _20866_/X _22044_/S vssd1 vssd1 vccd1 vccd1 _22037_/A sky130_fd_sc_hd__mux2_1
X_26913_ _26913_/CLK _26913_/D vssd1 vssd1 vccd1 vccd1 _26913_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26844_ _26877_/CLK _26844_/D vssd1 vssd1 vccd1 vccd1 _26844_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_130_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26775_ _26900_/CLK _26775_/D vssd1 vssd1 vccd1 vccd1 _26775_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23987_ _26868_/Q _23587_/X _23987_/S vssd1 vssd1 vccd1 vccd1 _23988_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13740_ _15791_/A _14604_/B _15134_/A vssd1 vssd1 vccd1 vccd1 _13740_/Y sky130_fd_sc_hd__nor3_1
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25726_ _26264_/CLK _25726_/D vssd1 vssd1 vccd1 vccd1 _25726_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22938_ _22938_/A vssd1 vssd1 vccd1 vccd1 _26444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_250_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25657_ _25660_/CLK _25657_/D vssd1 vssd1 vccd1 vccd1 _25657_/Q sky130_fd_sc_hd__dfxtp_1
X_13671_ _14725_/A _13671_/B _13671_/C vssd1 vssd1 vccd1 vccd1 _13671_/X sky130_fd_sc_hd__or3_1
X_22869_ _26414_/Q _22714_/X _22873_/S vssd1 vssd1 vccd1 vccd1 _22870_/A sky130_fd_sc_hd__mux2_1
XFILLER_188_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15410_ _16273_/S vssd1 vssd1 vccd1 vccd1 _16440_/S sky130_fd_sc_hd__buf_4
XFILLER_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24608_ hold1/A _24608_/B vssd1 vssd1 vccd1 vccd1 _24608_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16390_ _14877_/S _16387_/X _16389_/X _14661_/A vssd1 vssd1 vccd1 vccd1 _16390_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25588_ _26843_/CLK _25588_/D vssd1 vssd1 vccd1 vccd1 _25588_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15341_ _17793_/A _15342_/B vssd1 vssd1 vccd1 vccd1 _19158_/S sky130_fd_sc_hd__and2_2
X_27327_ _27327_/CLK _27327_/D vssd1 vssd1 vccd1 vccd1 _27327_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24539_ _27036_/Q _24372_/A _24538_/Y _24523_/X vssd1 vssd1 vccd1 vccd1 _27036_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18060_ _18254_/A _18057_/X _18059_/X vssd1 vssd1 vccd1 vccd1 _18061_/A sky130_fd_sc_hd__a21oi_1
XFILLER_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27258_ _27258_/CLK _27258_/D vssd1 vssd1 vccd1 vccd1 _27258_/Q sky130_fd_sc_hd__dfxtp_1
X_15272_ _16161_/S vssd1 vssd1 vccd1 vccd1 _16399_/S sky130_fd_sc_hd__buf_4
X_17011_ _16810_/A _17008_/X _16873_/B _17006_/X input242/X vssd1 vssd1 vccd1 vccd1
+ _17011_/X sky130_fd_sc_hd__a32o_4
X_26209_ _26974_/CLK _26209_/D vssd1 vssd1 vccd1 vccd1 _26209_/Q sky130_fd_sc_hd__dfxtp_1
X_14223_ _14221_/X _14222_/X _14223_/S vssd1 vssd1 vccd1 vccd1 _14223_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27189_ _27196_/CLK _27189_/D vssd1 vssd1 vccd1 vccd1 _27189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14154_ _14153_/X _26880_/Q _26752_/Q _14103_/X _13611_/A vssd1 vssd1 vccd1 vccd1
+ _14154_/X sky130_fd_sc_hd__a221o_1
XFILLER_125_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13105_ _13269_/A _13105_/B vssd1 vssd1 vccd1 vccd1 _14100_/A sky130_fd_sc_hd__nand2_8
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14085_ _14344_/S vssd1 vssd1 vccd1 vccd1 _14095_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18962_ _18552_/X _18944_/X _18961_/Y _18779_/X vssd1 vssd1 vccd1 vccd1 _18962_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13036_ _15964_/S vssd1 vssd1 vccd1 vccd1 _15453_/A sky130_fd_sc_hd__buf_2
X_17913_ _17908_/X _17911_/X _18071_/S vssd1 vssd1 vccd1 vccd1 _17913_/X sky130_fd_sc_hd__mux2_1
X_18893_ _25738_/Q _18892_/C _25739_/Q vssd1 vssd1 vccd1 vccd1 _18894_/B sky130_fd_sc_hd__a21oi_1
XFILLER_239_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17844_ _19109_/A _19121_/B vssd1 vssd1 vccd1 vccd1 _17844_/X sky130_fd_sc_hd__or2_1
XFILLER_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17775_ _17767_/X _18474_/A _17774_/X vssd1 vssd1 vccd1 vccd1 _17775_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_226_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14987_ _16521_/A _14987_/B _14987_/C vssd1 vssd1 vccd1 vccd1 _14987_/Y sky130_fd_sc_hd__nor3_1
XFILLER_93_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19514_ _25640_/Q _19523_/B vssd1 vssd1 vccd1 vccd1 _19514_/X sky130_fd_sc_hd__or2_1
X_16726_ _20800_/B vssd1 vssd1 vccd1 vccd1 _16726_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13938_ _13937_/X _25835_/Q _26035_/Q _15938_/S _13337_/A vssd1 vssd1 vccd1 vccd1
+ _13938_/X sky130_fd_sc_hd__a221o_1
XFILLER_223_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_500 _16943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_511 _17067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_522 _17037_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19445_ _19196_/X _19443_/Y _19444_/X _25161_/A _18777_/X vssd1 vssd1 vccd1 vccd1
+ _19445_/X sky130_fd_sc_hd__o32a_1
XFILLER_207_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_533 _17049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16657_ _16657_/A _16676_/A _16676_/B vssd1 vssd1 vccd1 vccd1 _20796_/B sky130_fd_sc_hd__nor3b_4
X_13869_ _14269_/S vssd1 vssd1 vccd1 vccd1 _15879_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_222_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_544 _25728_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_555 _25731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15608_ _13254_/A _26861_/Q _25775_/Q _16113_/A _15924_/A vssd1 vssd1 vccd1 vccd1
+ _15608_/X sky130_fd_sc_hd__a221o_1
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19376_ _18775_/X _19374_/Y _18382_/A vssd1 vssd1 vccd1 vccd1 _19376_/X sky130_fd_sc_hd__o21ba_1
XFILLER_195_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16588_ _18035_/A vssd1 vssd1 vccd1 vccd1 _16589_/B sky130_fd_sc_hd__inv_2
X_18327_ _18327_/A _18327_/B vssd1 vssd1 vccd1 vccd1 _18328_/B sky130_fd_sc_hd__and2_1
X_15539_ _15031_/A _15535_/X _15537_/X _15538_/X vssd1 vssd1 vccd1 vccd1 _15539_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_175_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18258_ _18042_/X _18051_/X _18262_/S vssd1 vssd1 vccd1 vccd1 _18258_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17209_ _17209_/A vssd1 vssd1 vccd1 vccd1 _25495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18189_ _18210_/S _18045_/X _17981_/Y vssd1 vssd1 vccd1 vccd1 _18344_/A sky130_fd_sc_hd__o21ai_1
XFILLER_129_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20220_ _19993_/X _20217_/X _20218_/Y _20219_/Y vssd1 vssd1 vccd1 vccd1 _20220_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20151_ _25678_/Q _25677_/Q _20151_/C vssd1 vssd1 vccd1 vccd1 _20164_/B sky130_fd_sc_hd__and3_1
XFILLER_277_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20082_ _20082_/A _20082_/B vssd1 vssd1 vccd1 vccd1 _20082_/Y sky130_fd_sc_hd__nor2_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23910_ _23910_/A vssd1 vssd1 vccd1 vccd1 _26833_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_257_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24890_ _27130_/Q _24890_/B vssd1 vssd1 vccd1 vccd1 _24890_/Y sky130_fd_sc_hd__nand2_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23841_ _23760_/X _26803_/Q _23843_/S vssd1 vssd1 vccd1 vccd1 _23842_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27303_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26560_ _27303_/CLK _26560_/D vssd1 vssd1 vccd1 vccd1 _26560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20984_ _26586_/Q _20986_/B _25867_/D vssd1 vssd1 vccd1 vccd1 _20985_/A sky130_fd_sc_hd__and3_1
X_23772_ _23772_/A vssd1 vssd1 vccd1 vccd1 _26774_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25511_ _27014_/CLK _25511_/D vssd1 vssd1 vccd1 vccd1 _25511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22723_ _23766_/A vssd1 vssd1 vccd1 vccd1 _22723_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26491_ _27298_/CLK _26491_/D vssd1 vssd1 vccd1 vccd1 _26491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25442_ _23754_/X _27316_/Q _25448_/S vssd1 vssd1 vccd1 vccd1 _25443_/A sky130_fd_sc_hd__mux2_1
X_22654_ _26331_/Q _22653_/X _22657_/S vssd1 vssd1 vccd1 vccd1 _22655_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21605_ input62/X input97/X _21615_/S vssd1 vssd1 vccd1 vccd1 _21606_/A sky130_fd_sc_hd__mux2_8
XFILLER_139_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22585_ _22580_/X _22584_/Y _22574_/X vssd1 vssd1 vccd1 vccd1 _26309_/D sky130_fd_sc_hd__a21oi_1
X_25373_ _25373_/A vssd1 vssd1 vccd1 vccd1 _27285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27112_ _27198_/CLK _27112_/D vssd1 vssd1 vccd1 vccd1 _27112_/Q sky130_fd_sc_hd__dfxtp_2
X_24324_ _26999_/Q _24326_/C _24323_/Y vssd1 vssd1 vccd1 vccd1 _26999_/D sky130_fd_sc_hd__o21a_1
X_21536_ _20681_/A _21481_/X _21459_/A _21535_/X vssd1 vssd1 vccd1 vccd1 _21536_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_139_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27043_ _27044_/CLK _27043_/D vssd1 vssd1 vccd1 vccd1 _27043_/Q sky130_fd_sc_hd__dfxtp_1
X_24255_ _26975_/Q _24258_/C _24209_/X vssd1 vssd1 vccd1 vccd1 _24255_/Y sky130_fd_sc_hd__a21oi_1
X_21467_ _21597_/A vssd1 vssd1 vccd1 vccd1 _21467_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23206_ _23206_/A vssd1 vssd1 vccd1 vccd1 _26549_/D sky130_fd_sc_hd__clkbuf_1
X_20418_ _20420_/B _20003_/X _20410_/X _20417_/X _20346_/X vssd1 vssd1 vccd1 vccd1
+ _25688_/D sky130_fd_sc_hd__o221a_1
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24186_ _26952_/Q _24183_/A _24185_/Y vssd1 vssd1 vccd1 vccd1 _26952_/D sky130_fd_sc_hd__o21a_1
XFILLER_175_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21398_ _21394_/Y _21397_/X _21359_/X vssd1 vssd1 vccd1 vccd1 _21398_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_135_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20349_ _25686_/Q _20382_/C vssd1 vssd1 vccd1 vccd1 _20349_/X sky130_fd_sc_hd__or2_1
XFILLER_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23137_ _26519_/Q _23136_/X _23137_/S vssd1 vssd1 vccd1 vccd1 _23138_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23068_ _23068_/A vssd1 vssd1 vccd1 vccd1 _26497_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput200 localMemory_wb_adr_i[19] vssd1 vssd1 vccd1 vccd1 input200/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput211 localMemory_wb_adr_i[7] vssd1 vssd1 vccd1 vccd1 input211/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput222 localMemory_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input222/X sky130_fd_sc_hd__buf_6
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14910_ _14765_/A _14908_/X _14909_/X _14760_/A vssd1 vssd1 vccd1 vccd1 _14910_/X
+ sky130_fd_sc_hd__o211a_1
X_22019_ _26121_/Q _20951_/X _22027_/S vssd1 vssd1 vccd1 vccd1 _22020_/A sky130_fd_sc_hd__mux2_1
Xinput233 localMemory_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 input233/X sky130_fd_sc_hd__buf_8
XTAP_5444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15890_ _26633_/Q _26729_/Q _15890_/S vssd1 vssd1 vccd1 vccd1 _15890_/X sky130_fd_sc_hd__mux2_1
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput244 localMemory_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input244/X sky130_fd_sc_hd__buf_6
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput255 manufacturerID[1] vssd1 vssd1 vccd1 vccd1 input255/X sky130_fd_sc_hd__buf_2
XTAP_5466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput266 partID[11] vssd1 vssd1 vccd1 vccd1 input266/X sky130_fd_sc_hd__clkbuf_1
XTAP_5477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput277 partID[7] vssd1 vssd1 vccd1 vccd1 input277/X sky130_fd_sc_hd__clkbuf_1
XTAP_5488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26827_ _26827_/CLK _26827_/D vssd1 vssd1 vccd1 vccd1 _26827_/Q sky130_fd_sc_hd__dfxtp_1
X_14841_ _16053_/S vssd1 vssd1 vccd1 vccd1 _16396_/S sky130_fd_sc_hd__buf_4
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ _17592_/A vssd1 vssd1 vccd1 vccd1 _17560_/X sky130_fd_sc_hd__buf_2
X_26758_ _27276_/CLK _26758_/D vssd1 vssd1 vccd1 vccd1 _26758_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14772_ _14772_/A vssd1 vssd1 vccd1 vccd1 _14773_/A sky130_fd_sc_hd__buf_2
XFILLER_245_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16511_ _16533_/A vssd1 vssd1 vccd1 vccd1 _16523_/S sky130_fd_sc_hd__buf_2
XFILLER_244_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13723_ _13723_/A vssd1 vssd1 vccd1 vccd1 _15633_/S sky130_fd_sc_hd__clkbuf_4
X_25709_ _27280_/CLK _25709_/D vssd1 vssd1 vccd1 vccd1 _25709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_260_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17491_ _17691_/B _17683_/B vssd1 vssd1 vccd1 vccd1 _21218_/C sky130_fd_sc_hd__nor2_1
XFILLER_95_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26689_ _26908_/CLK _26689_/D vssd1 vssd1 vccd1 vccd1 _26689_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19230_ _18437_/A _19220_/X _19229_/X vssd1 vssd1 vccd1 vccd1 _19230_/X sky130_fd_sc_hd__a21o_4
XFILLER_16_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16442_ _16440_/X _16441_/X _16442_/S vssd1 vssd1 vccd1 vccd1 _16442_/X sky130_fd_sc_hd__mux2_1
X_13654_ _14452_/S vssd1 vssd1 vccd1 vccd1 _14221_/S sky130_fd_sc_hd__buf_2
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19161_ _18359_/X _19157_/X _19160_/X _18738_/A vssd1 vssd1 vccd1 vccd1 _19161_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16373_ _17846_/C vssd1 vssd1 vccd1 vccd1 _19277_/A sky130_fd_sc_hd__clkbuf_2
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _13585_/A vssd1 vssd1 vccd1 vccd1 _13585_/X sky130_fd_sc_hd__clkbuf_2
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ _18293_/A vssd1 vssd1 vccd1 vccd1 _19060_/A sky130_fd_sc_hd__buf_2
XFILLER_169_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15324_ _15321_/X _26414_/Q _14729_/A _15323_/X vssd1 vssd1 vccd1 vccd1 _15324_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19092_ _27121_/Q _18504_/A _19090_/X _19091_/X vssd1 vssd1 vccd1 vccd1 _19092_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_219_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18043_ _18041_/X _18042_/X _18209_/S vssd1 vssd1 vccd1 vccd1 _18043_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15255_ _15255_/A vssd1 vssd1 vccd1 vccd1 _16315_/S sky130_fd_sc_hd__buf_4
XFILLER_173_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14206_ _15490_/A _26880_/Q _26752_/Q _15842_/S _12738_/C vssd1 vssd1 vccd1 vccd1
+ _14206_/X sky130_fd_sc_hd__a221o_1
X_15186_ _15285_/A _15186_/B vssd1 vssd1 vccd1 vccd1 _15186_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14137_ _13911_/X _17592_/B _14136_/X _12902_/X _25914_/Q vssd1 vssd1 vccd1 vccd1
+ _14138_/B sky130_fd_sc_hd__o32a_1
XFILLER_141_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19994_ _27145_/Q _27079_/Q vssd1 vssd1 vccd1 vccd1 _19999_/A sky130_fd_sc_hd__and2_1
XFILLER_98_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14068_ _14064_/X _14065_/X _14066_/X _14067_/X vssd1 vssd1 vccd1 vccd1 _14069_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18945_ _18945_/A vssd1 vssd1 vccd1 vccd1 _18947_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13019_ _14169_/B vssd1 vssd1 vccd1 vccd1 _14253_/S sky130_fd_sc_hd__buf_2
XFILLER_67_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18876_ _18806_/X _18866_/X _18875_/X vssd1 vssd1 vccd1 vccd1 _18876_/X sky130_fd_sc_hd__a21o_4
XFILLER_67_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17827_ _17816_/X _17825_/Y _17826_/X vssd1 vssd1 vccd1 vccd1 _17827_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17758_ _18238_/A vssd1 vssd1 vccd1 vccd1 _18756_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16709_ _22476_/A _16703_/X _16705_/X _18230_/B vssd1 vssd1 vccd1 vccd1 _16709_/X
+ sky130_fd_sc_hd__a22o_2
X_17689_ _17704_/S _19798_/A vssd1 vssd1 vccd1 vccd1 _17689_/X sky130_fd_sc_hd__or2_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_330 input179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_341 _19609_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_352 _19612_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19428_ _14831_/A _17779_/A _18733_/X _19427_/X vssd1 vssd1 vccd1 vccd1 _19428_/X
+ sky130_fd_sc_hd__a22o_1
XINSDIODE2_363 input233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_374 _16992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_385 _17004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_396 _17034_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19359_ _16561_/B _18368_/A _18548_/A vssd1 vssd1 vccd1 vccd1 _19359_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22370_ _17085_/A _26227_/Q _22376_/S vssd1 vssd1 vccd1 vccd1 _22371_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_152_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27213_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_149_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21321_ _21346_/A vssd1 vssd1 vccd1 vccd1 _21547_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_176_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21252_ _21586_/A _18133_/X _21587_/A _25798_/Q _21346_/A vssd1 vssd1 vccd1 vccd1
+ _21252_/X sky130_fd_sc_hd__a221o_1
X_24040_ _26891_/Q _23558_/X _24048_/S vssd1 vssd1 vccd1 vccd1 _24041_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20203_ _20145_/X _20200_/Y _20202_/X vssd1 vssd1 vccd1 vccd1 _20206_/B sky130_fd_sc_hd__a21o_1
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21183_ _21183_/A vssd1 vssd1 vccd1 vccd1 _25931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20134_ _20134_/A _20134_/B vssd1 vssd1 vccd1 vccd1 _20135_/B sky130_fd_sc_hd__nand2_1
XFILLER_277_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25991_ _27000_/CLK _25991_/D vssd1 vssd1 vccd1 vccd1 _25991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24942_ _24585_/A _24941_/X _24938_/X vssd1 vssd1 vccd1 vccd1 _24942_/Y sky130_fd_sc_hd__a21oi_1
X_20065_ _25675_/Q _20098_/C _20015_/A vssd1 vssd1 vccd1 vccd1 _20065_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_225_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_12 _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_23 _19119_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_34 _19315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24873_ _27125_/Q _24873_/B vssd1 vssd1 vccd1 vccd1 _24873_/Y sky130_fd_sc_hd__nand2_1
XINSDIODE2_45 _20630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_56 _20643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_67 _20664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26612_ _27287_/CLK _26612_/D vssd1 vssd1 vccd1 vccd1 _26612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23824_ _23734_/X _26795_/Q _23832_/S vssd1 vssd1 vccd1 vccd1 _23825_/A sky130_fd_sc_hd__mux2_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_78 _20699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_89 _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26543_ _27329_/A _26543_/D vssd1 vssd1 vccd1 vccd1 _26543_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23755_ _23754_/X _26769_/Q _23764_/S vssd1 vssd1 vccd1 vccd1 _23756_/A sky130_fd_sc_hd__mux2_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ _23782_/A vssd1 vssd1 vccd1 vccd1 _20967_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22706_ _22706_/A vssd1 vssd1 vccd1 vccd1 _26347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26474_ _27281_/CLK _26474_/D vssd1 vssd1 vccd1 vccd1 _26474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23686_ _23767_/A vssd1 vssd1 vccd1 vccd1 _23786_/S sky130_fd_sc_hd__buf_4
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ _25837_/Q _20897_/X _20901_/S vssd1 vssd1 vccd1 vccd1 _20899_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25425_ _25425_/A vssd1 vssd1 vccd1 vccd1 _27308_/D sky130_fd_sc_hd__clkbuf_1
X_22637_ _26326_/Q _22631_/A _22632_/C _22636_/Y _22402_/X vssd1 vssd1 vccd1 vccd1
+ _26326_/D sky130_fd_sc_hd__o221a_1
XFILLER_201_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13370_ _13322_/X _13327_/X _13369_/Y vssd1 vssd1 vccd1 vccd1 _13370_/Y sky130_fd_sc_hd__o21bai_4
X_25356_ _25378_/A vssd1 vssd1 vccd1 vccd1 _25365_/S sky130_fd_sc_hd__buf_4
X_22568_ _22607_/A vssd1 vssd1 vccd1 vccd1 _22578_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_221_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24307_ _26993_/Q _24309_/C _24306_/Y vssd1 vssd1 vccd1 vccd1 _26993_/D sky130_fd_sc_hd__o21a_1
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21519_ _21488_/X _21462_/X _21517_/Y _21518_/X vssd1 vssd1 vccd1 vccd1 _21519_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_155_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25287_ _23738_/X _27247_/Q _25293_/S vssd1 vssd1 vccd1 vccd1 _25288_/A sky130_fd_sc_hd__mux2_1
X_22499_ _22499_/A vssd1 vssd1 vccd1 vccd1 _26274_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27026_ _27154_/CLK _27026_/D vssd1 vssd1 vccd1 vccd1 _27026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15040_ _15040_/A vssd1 vssd1 vccd1 vccd1 _15040_/X sky130_fd_sc_hd__clkbuf_4
X_24238_ _26969_/Q _24240_/C _24237_/Y vssd1 vssd1 vccd1 vccd1 _26969_/D sky130_fd_sc_hd__o21a_1
XFILLER_79_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24169_ _26947_/Q _26946_/Q _24169_/C vssd1 vssd1 vccd1 vccd1 _24175_/C sky130_fd_sc_hd__and3_1
XFILLER_269_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16991_ _22474_/A _16988_/X _16990_/X _18151_/B vssd1 vssd1 vccd1 vccd1 _16991_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_268_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15942_ _15491_/A _27276_/Q _26469_/Q _15501_/A _13775_/A vssd1 vssd1 vccd1 vccd1
+ _15942_/X sky130_fd_sc_hd__a221o_1
XFILLER_150_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18730_ _18896_/A _18318_/X _18729_/X _18343_/A vssd1 vssd1 vccd1 vccd1 _18730_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18661_ _25543_/Q _18459_/X _18660_/X _18154_/A _18466_/X vssd1 vssd1 vccd1 vccd1
+ _18661_/X sky130_fd_sc_hd__a221o_1
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ _15954_/A _15954_/B _15873_/C vssd1 vssd1 vccd1 vccd1 _15873_/Y sky130_fd_sc_hd__nor3_1
XFILLER_64_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14824_ _14776_/Y _14788_/Y _14790_/X _14823_/Y vssd1 vssd1 vccd1 vccd1 _14824_/X
+ sky130_fd_sc_hd__o211a_1
X_17612_ _17612_/A vssd1 vssd1 vccd1 vccd1 _17612_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18592_ _18593_/B _18593_/C _18593_/A vssd1 vssd1 vccd1 vccd1 _18634_/B sky130_fd_sc_hd__o21a_1
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17543_ _17548_/A _17543_/B vssd1 vssd1 vccd1 vccd1 _25569_/D sky130_fd_sc_hd__nor2_1
XFILLER_251_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14755_ _14755_/A vssd1 vssd1 vccd1 vccd1 _14755_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_251_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13706_ _13706_/A vssd1 vssd1 vccd1 vccd1 _15734_/S sky130_fd_sc_hd__buf_4
XFILLER_205_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17474_ _26244_/Q _17455_/X _21206_/A _25972_/Q vssd1 vssd1 vccd1 vccd1 _21208_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_189_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14686_ _15168_/A vssd1 vssd1 vccd1 vccd1 _15048_/A sky130_fd_sc_hd__buf_4
XFILLER_204_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19213_ _25747_/Q _19246_/C vssd1 vssd1 vccd1 vccd1 _20279_/A sky130_fd_sc_hd__xnor2_2
X_16425_ _27322_/Q _26579_/Q _16440_/S vssd1 vssd1 vccd1 vccd1 _16425_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13637_ _15482_/A _16846_/A _13636_/Y _15868_/B vssd1 vssd1 vccd1 vccd1 _13689_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_220_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19144_ _19482_/B _19142_/Y _19143_/X _19121_/Y _19076_/X vssd1 vssd1 vccd1 vccd1
+ _19144_/X sky130_fd_sc_hd__o32a_2
X_16356_ _15111_/X _26417_/Q _16360_/S _16355_/X vssd1 vssd1 vccd1 vccd1 _16356_/X
+ sky130_fd_sc_hd__o211a_1
X_13568_ _12913_/A _13567_/Y _12929_/X vssd1 vssd1 vccd1 vccd1 _13568_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15307_ _25851_/Q _26051_/Q _16262_/S vssd1 vssd1 vccd1 vccd1 _15307_/X sky130_fd_sc_hd__mux2_1
X_19075_ _18666_/A _19073_/Y _17774_/X vssd1 vssd1 vccd1 vccd1 _19075_/X sky130_fd_sc_hd__o21a_1
X_16287_ _17795_/A _16287_/B vssd1 vssd1 vccd1 vccd1 _16288_/B sky130_fd_sc_hd__nor2_1
X_13499_ _14542_/A vssd1 vssd1 vccd1 vccd1 _14777_/A sky130_fd_sc_hd__buf_6
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18026_ _18721_/A vssd1 vssd1 vccd1 vccd1 _18144_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15238_ _17782_/A _17781_/A vssd1 vssd1 vccd1 vccd1 _19240_/S sky130_fd_sc_hd__nor2_1
XFILLER_114_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_160_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15169_ _15169_/A vssd1 vssd1 vccd1 vccd1 _15169_/X sky130_fd_sc_hd__buf_4
XFILLER_114_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19977_ _19950_/A _19977_/B vssd1 vssd1 vccd1 vccd1 _19977_/X sky130_fd_sc_hd__and2b_1
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18928_ _18895_/X _18909_/X _18926_/Y _18927_/X vssd1 vssd1 vccd1 vccd1 _18928_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_228_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18859_ _18859_/A _18859_/B vssd1 vssd1 vccd1 vccd1 _18859_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21870_ _21870_/A _21870_/B _24455_/A vssd1 vssd1 vccd1 vccd1 _24456_/A sky130_fd_sc_hd__nor3_2
XFILLER_270_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20821_ _20821_/A vssd1 vssd1 vccd1 vccd1 _25806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_270_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23540_ _26693_/Q _23539_/X _23540_/S vssd1 vssd1 vccd1 vccd1 _23541_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20752_ _20774_/A vssd1 vssd1 vccd1 vccd1 _20761_/S sky130_fd_sc_hd__buf_4
XINSDIODE2_160 _15292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_171 _14449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_182 _17818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20683_ _20683_/A _20683_/B vssd1 vssd1 vccd1 vccd1 _20683_/X sky130_fd_sc_hd__or2_1
XINSDIODE2_193 _17856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23471_ _23493_/A vssd1 vssd1 vccd1 vccd1 _23480_/S sky130_fd_sc_hd__buf_4
XFILLER_210_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25210_ _27053_/Q _21874_/A input171/X _25209_/X _25199_/A vssd1 vssd1 vccd1 vccd1
+ _25210_/X sky130_fd_sc_hd__a41o_1
X_22422_ _26193_/Q _22418_/X _22421_/X _22348_/X vssd1 vssd1 vccd1 vccd1 _26241_/D
+ sky130_fd_sc_hd__o211a_1
X_26190_ _26238_/CLK _26190_/D vssd1 vssd1 vccd1 vccd1 _26190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25141_ _19283_/A _25138_/X _25140_/X vssd1 vssd1 vccd1 vccd1 _25141_/X sky130_fd_sc_hd__o21a_1
X_22353_ _22337_/X _26231_/Q _22356_/A vssd1 vssd1 vccd1 vccd1 _22353_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_176_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21304_ _21276_/X _21303_/X _21227_/X vssd1 vssd1 vccd1 vccd1 _21304_/Y sky130_fd_sc_hd__o21ai_1
X_22284_ _22315_/A vssd1 vssd1 vccd1 vccd1 _22284_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25072_ _20654_/A _25059_/X _25071_/X vssd1 vssd1 vccd1 vccd1 _25072_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_164_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21235_ _21235_/A vssd1 vssd1 vccd1 vccd1 _21581_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_24023_ _24023_/A vssd1 vssd1 vccd1 vccd1 _26883_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21166_ _21166_/A vssd1 vssd1 vccd1 vccd1 _21166_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20117_ _20204_/A _20205_/B vssd1 vssd1 vccd1 vccd1 _20118_/B sky130_fd_sc_hd__and2b_1
XFILLER_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25974_ _27058_/CLK _25974_/D vssd1 vssd1 vccd1 vccd1 _25974_/Q sky130_fd_sc_hd__dfxtp_4
X_21097_ _21100_/A _21097_/B vssd1 vssd1 vccd1 vccd1 _21098_/A sky130_fd_sc_hd__or2_1
XFILLER_172_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24925_ _24569_/A _24917_/X _24909_/X vssd1 vssd1 vccd1 vccd1 _24925_/Y sky130_fd_sc_hd__a21oi_1
X_20048_ _20046_/X _20047_/Y _20022_/Y _20024_/Y vssd1 vssd1 vccd1 vccd1 _20048_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_219_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12870_ _14025_/A _12868_/Y _12869_/X vssd1 vssd1 vccd1 vccd1 _12871_/A sky130_fd_sc_hd__a21o_1
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24856_ _27120_/Q _24856_/B vssd1 vssd1 vccd1 vccd1 _24856_/Y sky130_fd_sc_hd__nand2_1
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23807_ _23807_/A vssd1 vssd1 vccd1 vccd1 _26787_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24787_ _24785_/Y _24786_/X _22634_/X vssd1 vssd1 vccd1 vccd1 _27102_/D sky130_fd_sc_hd__a21oi_1
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21999_ _26112_/Q _20923_/X _22005_/S vssd1 vssd1 vccd1 vccd1 _22000_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14453_/X _26096_/Q _25997_/Q _16021_/S _14384_/X vssd1 vssd1 vccd1 vccd1
+ _14540_/X sky130_fd_sc_hd__a221o_1
XFILLER_214_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26526_ _27238_/CLK _26526_/D vssd1 vssd1 vccd1 vccd1 _26526_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23738_ _23738_/A vssd1 vssd1 vccd1 vccd1 _23738_/X sky130_fd_sc_hd__buf_2
XFILLER_230_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26457_ _27266_/CLK _26457_/D vssd1 vssd1 vccd1 vccd1 _26457_/Q sky130_fd_sc_hd__dfxtp_1
X_14471_ _26521_/Q _26129_/Q _14472_/S vssd1 vssd1 vccd1 vccd1 _14471_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23669_ _23669_/A vssd1 vssd1 vccd1 vccd1 _23678_/S sky130_fd_sc_hd__buf_6
XFILLER_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ _16612_/A _16612_/B _19123_/A _16209_/X vssd1 vssd1 vccd1 vccd1 _19156_/B
+ sky130_fd_sc_hd__o31ai_4
X_13422_ _14349_/S vssd1 vssd1 vccd1 vccd1 _14115_/S sky130_fd_sc_hd__buf_2
X_25408_ _25408_/A vssd1 vssd1 vccd1 vccd1 _27300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17190_ _20646_/A vssd1 vssd1 vccd1 vccd1 _17190_/X sky130_fd_sc_hd__clkbuf_4
X_26388_ _27321_/CLK _26388_/D vssd1 vssd1 vccd1 vccd1 _26388_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16141_ _15142_/X _16138_/X _16140_/X _14660_/A vssd1 vssd1 vccd1 vccd1 _16141_/X
+ sky130_fd_sc_hd__a211o_1
X_25339_ _27270_/Q _23709_/A _25343_/S vssd1 vssd1 vccd1 vccd1 _25340_/A sky130_fd_sc_hd__mux2_1
X_13353_ _14389_/S vssd1 vssd1 vccd1 vccd1 _14310_/S sky130_fd_sc_hd__buf_2
XFILLER_127_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16072_ _16068_/X _16071_/X _16072_/S vssd1 vssd1 vccd1 vccd1 _16072_/X sky130_fd_sc_hd__mux2_1
X_13284_ _13284_/A vssd1 vssd1 vccd1 vccd1 _13321_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27009_ _27044_/CLK _27009_/D vssd1 vssd1 vccd1 vccd1 _27009_/Q sky130_fd_sc_hd__dfxtp_1
X_15023_ _16135_/B vssd1 vssd1 vccd1 vccd1 _15030_/S sky130_fd_sc_hd__buf_4
X_19900_ _19895_/X _19896_/Y _19898_/Y _19787_/A vssd1 vssd1 vccd1 vccd1 _19900_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_268_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19831_ _19830_/A _19830_/B _19830_/C vssd1 vssd1 vccd1 vccd1 _19831_/X sky130_fd_sc_hd__a21o_1
XFILLER_150_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19762_ _25665_/Q _19762_/B vssd1 vssd1 vccd1 vccd1 _19834_/C sky130_fd_sc_hd__and2_1
X_16974_ _16873_/X _16954_/X _16956_/X _16872_/X _16973_/X vssd1 vssd1 vccd1 vccd1
+ _16975_/C sky130_fd_sc_hd__a221o_1
XFILLER_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18713_ _25609_/Q _18973_/A _18013_/X _18712_/X vssd1 vssd1 vccd1 vccd1 _18714_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_265_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15925_ _13284_/A _15922_/X _15924_/X _13762_/X vssd1 vssd1 vccd1 vccd1 _15925_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19693_ _25663_/Q _25662_/Q vssd1 vssd1 vccd1 vccd1 _19693_/X sky130_fd_sc_hd__xor2_1
XFILLER_77_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput8 coreIndex[7] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15856_ _16195_/S _15854_/X _15855_/X _13274_/A vssd1 vssd1 vccd1 vccd1 _15856_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_188_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18644_ _18734_/A vssd1 vssd1 vccd1 vccd1 _19192_/B sky130_fd_sc_hd__buf_2
XFILLER_65_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14807_ _14807_/A vssd1 vssd1 vccd1 vccd1 _14808_/A sky130_fd_sc_hd__buf_2
XFILLER_224_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18575_ _25509_/Q _18559_/X _18567_/X _18573_/X _18574_/X vssd1 vssd1 vccd1 vccd1
+ _18575_/X sky130_fd_sc_hd__o221a_1
XFILLER_149_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15787_ _17826_/A _15788_/B vssd1 vssd1 vccd1 vccd1 _18901_/S sky130_fd_sc_hd__and2_2
XFILLER_80_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12999_ _20868_/B _13062_/A vssd1 vssd1 vccd1 vccd1 _13005_/B sky130_fd_sc_hd__xnor2_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14738_ _14905_/S vssd1 vssd1 vccd1 vccd1 _14811_/S sky130_fd_sc_hd__buf_2
X_17526_ _25903_/Q _17517_/X _14404_/B _17525_/X vssd1 vssd1 vccd1 vccd1 _17526_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17457_ _21198_/A _21870_/B vssd1 vssd1 vccd1 vccd1 _21244_/A sky130_fd_sc_hd__or2_4
XFILLER_178_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14669_ _14963_/S vssd1 vssd1 vccd1 vccd1 _14699_/S sky130_fd_sc_hd__buf_2
XFILLER_189_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16408_ _14683_/X _16383_/X _16391_/X _16407_/X vssd1 vssd1 vccd1 vccd1 _16408_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_221_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17388_ _17384_/X _17389_/C _25548_/Q vssd1 vssd1 vccd1 vccd1 _17390_/B sky130_fd_sc_hd__a21oi_1
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19127_ _19123_/A _18368_/X _19125_/X _19126_/X vssd1 vssd1 vccd1 vccd1 _19127_/X
+ sky130_fd_sc_hd__o211a_1
X_16339_ _16336_/X _16337_/X _16338_/X vssd1 vssd1 vccd1 vccd1 _16339_/X sky130_fd_sc_hd__o21a_1
XFILLER_146_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19058_ _19058_/A vssd1 vssd1 vccd1 vccd1 _19058_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput301 _16999_/X vssd1 vssd1 vccd1 vccd1 addr1[7] sky130_fd_sc_hd__buf_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput312 _16752_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[16] sky130_fd_sc_hd__buf_2
XFILLER_160_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18009_ _18552_/A vssd1 vssd1 vccd1 vccd1 _18895_/A sky130_fd_sc_hd__buf_2
Xoutput323 _16779_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[26] sky130_fd_sc_hd__buf_2
Xoutput334 _16811_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[0] sky130_fd_sc_hd__buf_2
Xoutput345 _16815_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[1] sky130_fd_sc_hd__buf_2
X_21020_ _25880_/Q _20907_/X _21026_/S vssd1 vssd1 vccd1 vccd1 _21021_/A sky130_fd_sc_hd__mux2_1
Xoutput356 _16819_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[2] sky130_fd_sc_hd__buf_2
Xoutput367 _16793_/X vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[1] sky130_fd_sc_hd__buf_2
XFILLER_273_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput378 _17023_/X vssd1 vssd1 vccd1 vccd1 din0[11] sky130_fd_sc_hd__buf_2
XFILLER_99_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput389 _17037_/X vssd1 vssd1 vccd1 vccd1 din0[21] sky130_fd_sc_hd__buf_2
XFILLER_206_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22971_ _26459_/Q _22653_/X _22973_/S vssd1 vssd1 vccd1 vccd1 _22972_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24710_ _24948_/A vssd1 vssd1 vccd1 vccd1 _24711_/B sky130_fd_sc_hd__inv_2
X_21922_ _20550_/X _26078_/Q _21922_/S vssd1 vssd1 vccd1 vccd1 _21923_/A sky130_fd_sc_hd__mux2_1
X_25690_ _25690_/CLK _25690_/D vssd1 vssd1 vccd1 vccd1 _25690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24641_ _24641_/A _24740_/A vssd1 vssd1 vccd1 vccd1 _24744_/A sky130_fd_sc_hd__and2_1
XFILLER_282_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21853_ _21853_/A vssd1 vssd1 vccd1 vccd1 _26054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20804_ _25798_/Q vssd1 vssd1 vccd1 vccd1 _20805_/A sky130_fd_sc_hd__clkbuf_1
X_24572_ _24572_/A _24582_/B vssd1 vssd1 vccd1 vccd1 _24572_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21784_ _21784_/A vssd1 vssd1 vccd1 vccd1 _26024_/D sky130_fd_sc_hd__clkbuf_1
X_26311_ _26322_/CLK _26311_/D vssd1 vssd1 vccd1 vccd1 _26311_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_196_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23523_ _23523_/A vssd1 vssd1 vccd1 vccd1 _23523_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20735_ _20521_/X _25765_/Q _20739_/S vssd1 vssd1 vccd1 vccd1 _20736_/A sky130_fd_sc_hd__mux2_1
X_27291_ _27291_/CLK _27291_/D vssd1 vssd1 vccd1 vccd1 _27291_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26242_ _26248_/CLK _26242_/D vssd1 vssd1 vccd1 vccd1 _26242_/Q sky130_fd_sc_hd__dfxtp_1
X_23454_ _26659_/Q _23060_/X _23458_/S vssd1 vssd1 vccd1 vccd1 _23455_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20666_ _20666_/A _20670_/B vssd1 vssd1 vccd1 vccd1 _20666_/X sky130_fd_sc_hd__or2_1
XFILLER_52_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22405_ _22405_/A _22405_/B vssd1 vssd1 vccd1 vccd1 _22405_/X sky130_fd_sc_hd__and2_1
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26173_ _26238_/CLK _26173_/D vssd1 vssd1 vccd1 vccd1 _26173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23385_ _23385_/A vssd1 vssd1 vccd1 vccd1 _26628_/D sky130_fd_sc_hd__clkbuf_1
X_20597_ _20597_/A vssd1 vssd1 vccd1 vccd1 _20614_/S sky130_fd_sc_hd__buf_6
XFILLER_167_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25124_ _25124_/A vssd1 vssd1 vccd1 vccd1 _25124_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22336_ _17085_/C input188/X _22340_/S vssd1 vssd1 vccd1 vccd1 _22336_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25055_ _25109_/A vssd1 vssd1 vccd1 vccd1 _25055_/X sky130_fd_sc_hd__clkbuf_2
X_22267_ _26201_/Q _22264_/X _22255_/X _26302_/Q _22256_/X vssd1 vssd1 vccd1 vccd1
+ _22267_/X sky130_fd_sc_hd__a221o_1
XFILLER_2_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24006_ _24074_/S vssd1 vssd1 vccd1 vccd1 _24015_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21218_ _21221_/B _17683_/A _21218_/C _21218_/D vssd1 vssd1 vccd1 vccd1 _21285_/A
+ sky130_fd_sc_hd__and4bb_1
X_22198_ _26183_/Q _22186_/X _22115_/X _22197_/X _22187_/X vssd1 vssd1 vccd1 vccd1
+ _22198_/X sky130_fd_sc_hd__a221o_1
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21149_ _21167_/A vssd1 vssd1 vccd1 vccd1 _21149_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25957_ _26995_/CLK _25957_/D vssd1 vssd1 vccd1 vccd1 _25957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13971_ _14391_/S vssd1 vssd1 vccd1 vccd1 _14369_/S sky130_fd_sc_hd__buf_2
XFILLER_262_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15710_ _25645_/Q _15443_/B _14612_/A vssd1 vssd1 vccd1 vccd1 _15710_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_18_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24908_ _27134_/Q _24902_/X _24907_/Y vssd1 vssd1 vccd1 vccd1 _27134_/D sky130_fd_sc_hd__o21a_1
X_12922_ _17623_/B _12922_/B vssd1 vssd1 vccd1 vccd1 _12922_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16690_ _25757_/Q _20800_/B vssd1 vssd1 vccd1 vccd1 _16691_/A sky130_fd_sc_hd__and2_2
XFILLER_74_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25888_ _26796_/CLK _25888_/D vssd1 vssd1 vccd1 vccd1 _25888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15641_ _25845_/Q _26045_/Q _15643_/S vssd1 vssd1 vccd1 vccd1 _15641_/X sky130_fd_sc_hd__mux2_1
X_12853_ _12837_/A _12934_/A _17592_/C _12899_/A _25917_/Q vssd1 vssd1 vccd1 vccd1
+ _15708_/A sky130_fd_sc_hd__o32a_2
X_24839_ _24837_/Y _24838_/X _24835_/X vssd1 vssd1 vccd1 vccd1 _27115_/D sky130_fd_sc_hd__a21oi_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18360_ _19046_/B _19572_/A _18357_/X _18359_/X vssd1 vssd1 vccd1 vccd1 _18360_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _15659_/A _16896_/A vssd1 vssd1 vccd1 vccd1 _15572_/Y sky130_fd_sc_hd__nor2_1
X_12784_ _25691_/Q _25690_/Q _25689_/Q vssd1 vssd1 vccd1 vccd1 _16685_/B sky130_fd_sc_hd__or3_2
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _17308_/X _17312_/C _25524_/Q vssd1 vssd1 vccd1 vccd1 _17313_/B sky130_fd_sc_hd__a21oi_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14523_ _14523_/A _14523_/B vssd1 vssd1 vccd1 vccd1 _14523_/X sky130_fd_sc_hd__and2_1
XFILLER_202_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26509_ _27315_/CLK _26509_/D vssd1 vssd1 vccd1 vccd1 _26509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18291_ _27203_/Q _18813_/A vssd1 vssd1 vccd1 vccd1 _18291_/X sky130_fd_sc_hd__and2_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17242_/A _17242_/B _25503_/Q vssd1 vssd1 vccd1 vccd1 _17243_/C sky130_fd_sc_hd__and3_1
XFILLER_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14454_ _14453_/X _26589_/Q _14308_/S _26329_/Q _14552_/S vssd1 vssd1 vccd1 vccd1
+ _14454_/X sky130_fd_sc_hd__o221a_1
XFILLER_186_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13405_ _13589_/S vssd1 vssd1 vccd1 vccd1 _13719_/A sky130_fd_sc_hd__buf_4
XFILLER_174_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17173_ _16526_/S _17170_/X _17172_/X _17134_/X vssd1 vssd1 vccd1 vccd1 _25483_/D
+ sky130_fd_sc_hd__o211a_1
X_14385_ _12736_/A _25831_/Q _26031_/Q _14375_/S _14384_/X vssd1 vssd1 vccd1 vccd1
+ _14385_/X sky130_fd_sc_hd__a221o_1
XFILLER_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16124_ _16124_/A _17842_/B vssd1 vssd1 vccd1 vccd1 _16124_/Y sky130_fd_sc_hd__nand2_1
X_13336_ _13336_/A vssd1 vssd1 vccd1 vccd1 _13337_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16055_ _25816_/Q _16163_/S _15633_/S _16054_/X vssd1 vssd1 vccd1 vccd1 _16055_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13267_ _15331_/A vssd1 vssd1 vccd1 vccd1 _13267_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15006_ _14746_/A _26616_/Q _14905_/S _26356_/Q _14917_/X vssd1 vssd1 vccd1 vccd1
+ _15006_/X sky130_fd_sc_hd__o221a_1
XFILLER_155_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13198_ _13641_/A _25581_/Q vssd1 vssd1 vccd1 vccd1 _14043_/A sky130_fd_sc_hd__nand2_2
XFILLER_123_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19814_ _27139_/Q _27073_/Q vssd1 vssd1 vccd1 vccd1 _19814_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19745_ _19745_/A _19745_/B vssd1 vssd1 vccd1 vccd1 _19745_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16957_ _16957_/A _16957_/B vssd1 vssd1 vccd1 vccd1 _16957_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15908_ _15900_/X _15907_/X _13107_/A vssd1 vssd1 vccd1 vccd1 _15908_/X sky130_fd_sc_hd__o21a_1
XFILLER_237_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19676_ _19676_/A vssd1 vssd1 vccd1 vccd1 _19833_/A sky130_fd_sc_hd__buf_2
X_16888_ _16932_/B vssd1 vssd1 vccd1 vccd1 _16927_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_264_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18627_ _18027_/X _18590_/X _18607_/X _18721_/A _18626_/X vssd1 vssd1 vccd1 vccd1
+ _18627_/X sky130_fd_sc_hd__o2111a_1
X_15839_ _15488_/X _26890_/Q _26762_/Q _15671_/S _15401_/A vssd1 vssd1 vccd1 vccd1
+ _15839_/X sky130_fd_sc_hd__a221o_1
XFILLER_213_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18558_ _25509_/Q _18556_/X _18557_/X _17365_/X vssd1 vssd1 vccd1 vccd1 _18558_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17509_ _19583_/A _18182_/B vssd1 vssd1 vccd1 vccd1 _18088_/A sky130_fd_sc_hd__and2_1
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18489_ _18265_/X _18261_/X _18489_/S vssd1 vssd1 vccd1 vccd1 _18489_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20520_ _23533_/A vssd1 vssd1 vccd1 vccd1 _23709_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_166_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_59_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26601_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_220_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20451_ _20450_/A _20450_/B _20450_/C vssd1 vssd1 vccd1 vccd1 _20471_/B sky130_fd_sc_hd__a21o_1
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23170_ _26533_/Q _23079_/X _23172_/S vssd1 vssd1 vccd1 vccd1 _23171_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20382_ _25687_/Q _25686_/Q _20382_/C vssd1 vssd1 vccd1 vccd1 _20420_/C sky130_fd_sc_hd__and3_1
XFILLER_119_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22121_ _22121_/A _22170_/A vssd1 vssd1 vccd1 vccd1 _22122_/A sky130_fd_sc_hd__or2_1
XFILLER_173_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22052_ _22052_/A vssd1 vssd1 vccd1 vccd1 _26135_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21003_ _21003_/A vssd1 vssd1 vccd1 vccd1 _25872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26860_ _27311_/CLK _26860_/D vssd1 vssd1 vccd1 vccd1 _26860_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25811_ _26881_/CLK _25811_/D vssd1 vssd1 vccd1 vccd1 _25811_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_229_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26791_ _27330_/A _26791_/D vssd1 vssd1 vccd1 vccd1 _26791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25742_ _26282_/CLK _25742_/D vssd1 vssd1 vccd1 vccd1 _25742_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22954_ _26452_/Q _22733_/X _22956_/S vssd1 vssd1 vccd1 vccd1 _22955_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21905_ _20517_/X _26070_/Q _21911_/S vssd1 vssd1 vccd1 vccd1 _21906_/A sky130_fd_sc_hd__mux2_1
XFILLER_260_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25673_ _25673_/CLK _25673_/D vssd1 vssd1 vccd1 vccd1 _25673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22885_ _22885_/A vssd1 vssd1 vccd1 vccd1 _26421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24624_ _27065_/Q _24615_/X _24623_/Y _24619_/X vssd1 vssd1 vccd1 vccd1 _27065_/D
+ sky130_fd_sc_hd__o211a_1
X_21836_ _26047_/Q _20929_/X _21838_/S vssd1 vssd1 vccd1 vccd1 _21837_/A sky130_fd_sc_hd__mux2_1
XFILLER_270_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24555_ _24561_/A vssd1 vssd1 vccd1 vccd1 _24610_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_168_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21767_ _21778_/A vssd1 vssd1 vccd1 vccd1 _21776_/S sky130_fd_sc_hd__buf_4
XFILLER_200_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23506_ _26683_/Q _23136_/X _23506_/S vssd1 vssd1 vccd1 vccd1 _23507_/A sky130_fd_sc_hd__mux2_1
X_27274_ _27277_/CLK _27274_/D vssd1 vssd1 vccd1 vccd1 _27274_/Q sky130_fd_sc_hd__dfxtp_4
X_20718_ _20774_/A vssd1 vssd1 vccd1 vccd1 _20787_/S sky130_fd_sc_hd__buf_6
XFILLER_178_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24486_ _24472_/X _25619_/Q _24485_/X vssd1 vssd1 vccd1 vccd1 _24732_/B sky130_fd_sc_hd__o21a_4
XFILLER_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21698_ _21698_/A vssd1 vssd1 vccd1 vccd1 _21707_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_200_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26225_ _27297_/CLK _26225_/D vssd1 vssd1 vccd1 vccd1 _26225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23437_ _23493_/A vssd1 vssd1 vccd1 vccd1 _23506_/S sky130_fd_sc_hd__buf_6
X_20649_ _26270_/Q _20646_/X _20648_/X _20644_/X vssd1 vssd1 vccd1 vccd1 _25733_/D
+ sky130_fd_sc_hd__o211a_1
X_14170_ _14153_/X _26396_/Q _14178_/S _14169_/X vssd1 vssd1 vccd1 vccd1 _14170_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26156_ _26453_/CLK _26156_/D vssd1 vssd1 vccd1 vccd1 _26156_/Q sky130_fd_sc_hd__dfxtp_2
X_23368_ _23368_/A vssd1 vssd1 vccd1 vccd1 _26620_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13121_ _13185_/A _13121_/B vssd1 vssd1 vccd1 vccd1 _14331_/A sky130_fd_sc_hd__nand2_4
XFILLER_180_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25107_ _22511_/A _25092_/X _25087_/X _19046_/A _25106_/X vssd1 vssd1 vccd1 vccd1
+ _25107_/X sky130_fd_sc_hd__a221o_1
X_22319_ _22428_/A vssd1 vssd1 vccd1 vccd1 _22319_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26087_ _27287_/CLK _26087_/D vssd1 vssd1 vccd1 vccd1 _26087_/Q sky130_fd_sc_hd__dfxtp_1
X_23299_ _23299_/A vssd1 vssd1 vccd1 vccd1 _26590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13052_ _13038_/X _13045_/X _15168_/A vssd1 vssd1 vccd1 vccd1 _13052_/X sky130_fd_sc_hd__mux2_1
X_25038_ _25065_/A vssd1 vssd1 vccd1 vccd1 _25038_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17860_ _18076_/A _18194_/B vssd1 vssd1 vccd1 vccd1 _18597_/A sky130_fd_sc_hd__nand2_2
XFILLER_267_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16811_ _16811_/A vssd1 vssd1 vccd1 vccd1 _16811_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_266_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17791_ _17791_/A _16206_/B vssd1 vssd1 vccd1 vccd1 _17791_/X sky130_fd_sc_hd__or2b_1
XFILLER_47_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26989_ _26996_/CLK _26989_/D vssd1 vssd1 vccd1 vccd1 _26989_/Q sky130_fd_sc_hd__dfxtp_1
X_19530_ _25646_/Q _19536_/B vssd1 vssd1 vccd1 vccd1 _19530_/X sky130_fd_sc_hd__or2_1
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13954_ _14542_/A _13954_/B _13954_/C vssd1 vssd1 vccd1 vccd1 _13954_/X sky130_fd_sc_hd__or3_1
X_16742_ _16769_/A vssd1 vssd1 vccd1 vccd1 _16742_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_219_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12905_ _12911_/A _12911_/B _15706_/B _15706_/C vssd1 vssd1 vccd1 vccd1 _15954_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19461_ _17336_/X _18743_/X _18744_/X _25564_/Q vssd1 vssd1 vccd1 vccd1 _19461_/X
+ sky130_fd_sc_hd__a22o_1
X_16673_ _16673_/A _21603_/A _16673_/C _16673_/D vssd1 vssd1 vccd1 vccd1 _16674_/A
+ sky130_fd_sc_hd__nor4_4
XFILLER_235_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13885_ _13880_/X _13884_/X _15983_/S vssd1 vssd1 vccd1 vccd1 _13885_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18412_ _18412_/A vssd1 vssd1 vccd1 vccd1 _25603_/D sky130_fd_sc_hd__clkbuf_1
X_12836_ _25795_/Q vssd1 vssd1 vccd1 vccd1 _12837_/A sky130_fd_sc_hd__inv_2
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15624_ _15167_/A _26408_/Q _15141_/A _15623_/X vssd1 vssd1 vccd1 vccd1 _15624_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19392_ _19392_/A _19392_/B vssd1 vssd1 vccd1 vccd1 _19392_/Y sky130_fd_sc_hd__nor2_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15555_ _25846_/Q _26046_/Q _15555_/S vssd1 vssd1 vccd1 vccd1 _15555_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18343_ _18343_/A vssd1 vssd1 vccd1 vccd1 _18547_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _12767_/A vssd1 vssd1 vccd1 vccd1 _12768_/A sky130_fd_sc_hd__buf_2
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _12674_/A _26488_/Q _26360_/Q _15972_/B _13140_/A vssd1 vssd1 vccd1 vccd1
+ _14506_/X sky130_fd_sc_hd__o221a_1
XFILLER_188_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18274_ _18859_/A _18273_/Y _17988_/A vssd1 vssd1 vccd1 vccd1 _19358_/B sky130_fd_sc_hd__o21ai_2
X_15486_ _15486_/A _15486_/B vssd1 vssd1 vccd1 vccd1 _15486_/X sky130_fd_sc_hd__or2_1
XFILLER_175_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12698_ _13121_/B vssd1 vssd1 vccd1 vccd1 _13630_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_202_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14437_ _26521_/Q _26129_/Q _14514_/S vssd1 vssd1 vccd1 vccd1 _14437_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17225_ _17107_/X _17224_/Y _17120_/X vssd1 vssd1 vccd1 vccd1 _25500_/D sky130_fd_sc_hd__o21ai_1
Xinput11 core_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput22 core_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput33 core_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput44 dout0[10] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_2
X_17156_ _22817_/A _17151_/X _17146_/X _17669_/B vssd1 vssd1 vccd1 vccd1 _17157_/B
+ sky130_fd_sc_hd__a22o_1
X_14368_ _13653_/S _14365_/X _14367_/X _13278_/A vssd1 vssd1 vccd1 vccd1 _14368_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_156_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput55 dout0[20] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput66 dout0[30] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_2
Xinput77 dout0[40] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16107_ _15676_/X _26115_/Q _26016_/Q _16273_/S _15672_/A vssd1 vssd1 vccd1 vccd1
+ _16107_/X sky130_fd_sc_hd__a221o_1
XFILLER_116_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput88 dout0[50] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__clkbuf_1
X_13319_ _15841_/S vssd1 vssd1 vccd1 vccd1 _15671_/S sky130_fd_sc_hd__buf_4
XFILLER_7_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17087_ _17087_/A _17091_/C _17087_/C _17085_/C vssd1 vssd1 vccd1 vccd1 _22416_/B
+ sky130_fd_sc_hd__nor4b_2
XFILLER_182_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput99 dout0[60] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14299_ _14542_/A _14299_/B _14299_/C vssd1 vssd1 vccd1 vccd1 _14299_/X sky130_fd_sc_hd__or3_1
XFILLER_182_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16038_ _17829_/A _16038_/B vssd1 vssd1 vccd1 vccd1 _18801_/S sky130_fd_sc_hd__nand2_1
XFILLER_192_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_177_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25590_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_258_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_106_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26327_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_229_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17989_ _17967_/X _18898_/B _17988_/X vssd1 vssd1 vccd1 vccd1 _17989_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_123_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19728_ _19728_/A _19910_/A vssd1 vssd1 vccd1 vccd1 _19728_/X sky130_fd_sc_hd__or2_1
XFILLER_238_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19659_ _19659_/A _19659_/B vssd1 vssd1 vccd1 vccd1 _19659_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22670_ _26336_/Q _22669_/X _22673_/S vssd1 vssd1 vccd1 vccd1 _22671_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21621_ _21586_/X _19407_/X _21587_/X _25826_/Q _21346_/X vssd1 vssd1 vccd1 vccd1
+ _21621_/X sky130_fd_sc_hd__a221o_1
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24340_ _25488_/Q _21208_/A _24340_/S vssd1 vssd1 vccd1 vccd1 _24900_/C sky130_fd_sc_hd__mux2_2
X_21552_ _21552_/A vssd1 vssd1 vccd1 vccd1 _21552_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_240_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20503_ _23520_/A vssd1 vssd1 vccd1 vccd1 _23696_/A sky130_fd_sc_hd__clkbuf_4
X_24271_ _24938_/A vssd1 vssd1 vccd1 vccd1 _24271_/X sky130_fd_sc_hd__buf_2
X_21483_ _21547_/A vssd1 vssd1 vccd1 vccd1 _21483_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_194_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26010_ _27307_/CLK _26010_/D vssd1 vssd1 vccd1 vccd1 _26010_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_165_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23222_ _26556_/Q _23050_/X _23222_/S vssd1 vssd1 vccd1 vccd1 _23223_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20434_ _20434_/A _20434_/B vssd1 vssd1 vccd1 vccd1 _20434_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23153_ _26525_/Q _23053_/X _23161_/S vssd1 vssd1 vccd1 vccd1 _23154_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20365_ _20350_/X _20362_/X _20364_/X vssd1 vssd1 vccd1 vccd1 _20365_/X sky130_fd_sc_hd__o21a_1
X_22104_ _22104_/A vssd1 vssd1 vccd1 vccd1 _26159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23084_ _23084_/A vssd1 vssd1 vccd1 vccd1 _26502_/D sky130_fd_sc_hd__clkbuf_1
X_20296_ _19649_/A _20293_/Y _20294_/X _20295_/X vssd1 vssd1 vccd1 vccd1 _20296_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22035_ _22103_/S vssd1 vssd1 vccd1 vccd1 _22044_/S sky130_fd_sc_hd__buf_2
X_26912_ _26913_/CLK _26912_/D vssd1 vssd1 vccd1 vccd1 _26912_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26843_ _26843_/CLK _26843_/D vssd1 vssd1 vccd1 vccd1 _26843_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26774_ _27322_/CLK _26774_/D vssd1 vssd1 vccd1 vccd1 _26774_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23986_ _23986_/A vssd1 vssd1 vccd1 vccd1 _26867_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25725_ _25725_/CLK _25725_/D vssd1 vssd1 vccd1 vccd1 _25725_/Q sky130_fd_sc_hd__dfxtp_4
X_22937_ _26444_/Q _22707_/X _22945_/S vssd1 vssd1 vccd1 vccd1 _22938_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25656_ _26248_/CLK _25656_/D vssd1 vssd1 vccd1 vccd1 _25656_/Q sky130_fd_sc_hd__dfxtp_1
X_13670_ _13791_/A _13668_/X _13669_/X _12754_/A vssd1 vssd1 vccd1 vccd1 _13671_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22868_ _22868_/A vssd1 vssd1 vccd1 vccd1 _26413_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24607_ _27058_/Q _24602_/X _24605_/Y _24606_/X vssd1 vssd1 vccd1 vccd1 _27058_/D
+ sky130_fd_sc_hd__o211a_1
X_21819_ _26039_/Q _20903_/X _21827_/S vssd1 vssd1 vccd1 vccd1 _21820_/A sky130_fd_sc_hd__mux2_1
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25587_ _26684_/CLK _25587_/D vssd1 vssd1 vccd1 vccd1 _25587_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22799_ _22799_/A vssd1 vssd1 vccd1 vccd1 _26383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27326_ _27326_/CLK _27326_/D vssd1 vssd1 vccd1 vccd1 _27326_/Q sky130_fd_sc_hd__dfxtp_1
X_15340_ _25746_/Q _15339_/Y _16368_/S vssd1 vssd1 vccd1 vccd1 _15342_/B sky130_fd_sc_hd__mux2_2
XPHY_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24538_ _24538_/A _24629_/A vssd1 vssd1 vccd1 vccd1 _24538_/Y sky130_fd_sc_hd__nand2_1
XPHY_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15271_ _26674_/Q _25714_/Q _16325_/S vssd1 vssd1 vccd1 vccd1 _15271_/X sky130_fd_sc_hd__mux2_1
X_27257_ _27257_/CLK _27257_/D vssd1 vssd1 vccd1 vccd1 _27257_/Q sky130_fd_sc_hd__dfxtp_1
X_24469_ _24492_/A hold2/A vssd1 vssd1 vccd1 vccd1 _24469_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17010_ _16810_/A _17008_/X _16868_/B _17006_/X input241/X vssd1 vssd1 vccd1 vccd1
+ _17010_/X sky130_fd_sc_hd__a32o_4
X_26208_ _26322_/CLK _26208_/D vssd1 vssd1 vccd1 vccd1 _26208_/Q sky130_fd_sc_hd__dfxtp_1
X_14222_ _27267_/Q _26460_/Q _14289_/S vssd1 vssd1 vccd1 vccd1 _14222_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27188_ _27188_/CLK _27188_/D vssd1 vssd1 vccd1 vccd1 _27188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26139_ _26599_/CLK _26139_/D vssd1 vssd1 vccd1 vccd1 _26139_/Q sky130_fd_sc_hd__dfxtp_4
X_14153_ _14153_/A vssd1 vssd1 vccd1 vccd1 _14153_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_4_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_4_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27283_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13104_ _13080_/X _13093_/X _13103_/X _16072_/S _12702_/A vssd1 vssd1 vccd1 vccd1
+ _13104_/X sky130_fd_sc_hd__o221a_1
XFILLER_153_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14084_ _14431_/A _14082_/X _14083_/X vssd1 vssd1 vccd1 vccd1 _14084_/X sky130_fd_sc_hd__o21a_1
X_18961_ _19219_/A _18968_/B _18960_/X vssd1 vssd1 vccd1 vccd1 _18961_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13035_ _15725_/S vssd1 vssd1 vccd1 vccd1 _15964_/S sky130_fd_sc_hd__clkbuf_4
X_17912_ _17975_/A vssd1 vssd1 vccd1 vccd1 _18071_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_152_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18892_ _25739_/Q _25738_/Q _18892_/C vssd1 vssd1 vccd1 vccd1 _18964_/B sky130_fd_sc_hd__and3_1
XFILLER_67_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17843_ _19048_/A _17841_/Y _17842_/X vssd1 vssd1 vccd1 vccd1 _19109_/C sky130_fd_sc_hd__a21oi_2
XFILLER_78_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17774_ _18998_/A vssd1 vssd1 vccd1 vccd1 _17774_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_266_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14986_ _14766_/A _14984_/X _14985_/X _12757_/A vssd1 vssd1 vccd1 vccd1 _14987_/C
+ sky130_fd_sc_hd__o211a_1
X_19513_ _19568_/B vssd1 vssd1 vccd1 vccd1 _19523_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_19_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16725_ _25668_/Q vssd1 vssd1 vccd1 vccd1 _22487_/A sky130_fd_sc_hd__buf_4
X_13937_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13937_/X sky130_fd_sc_hd__buf_2
XFILLER_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_501 _16986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19444_ _18947_/A _19442_/Y _18998_/X vssd1 vssd1 vccd1 vccd1 _19444_/X sky130_fd_sc_hd__o21a_1
XINSDIODE2_512 _17067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13868_ _13866_/X _13867_/X _14254_/S vssd1 vssd1 vccd1 vccd1 _13868_/X sky130_fd_sc_hd__mux2_1
XFILLER_223_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16656_ _21195_/B _16989_/A vssd1 vssd1 vccd1 vccd1 _16676_/B sky130_fd_sc_hd__or2b_2
XINSDIODE2_523 _17040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_534 _17049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_545 _17052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_556 _25983_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12819_ _25474_/Q vssd1 vssd1 vccd1 vccd1 _21320_/A sky130_fd_sc_hd__clkbuf_2
X_15607_ _13254_/A _26925_/Q _26409_/Q _16113_/A _15916_/A vssd1 vssd1 vccd1 vccd1
+ _15607_/X sky130_fd_sc_hd__a221o_1
XFILLER_250_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19375_ _18608_/X _19373_/X _19374_/Y vssd1 vssd1 vccd1 vccd1 _19375_/Y sky130_fd_sc_hd__a21oi_1
X_16587_ _16962_/A _17998_/A vssd1 vssd1 vccd1 vccd1 _18035_/A sky130_fd_sc_hd__xor2_4
X_13799_ _14833_/A _19849_/A _13798_/X vssd1 vssd1 vccd1 vccd1 _17818_/B sky130_fd_sc_hd__o21a_4
XFILLER_210_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18326_ _18327_/A _18327_/B vssd1 vssd1 vccd1 vccd1 _18328_/A sky130_fd_sc_hd__nor2_2
X_15538_ _15538_/A vssd1 vssd1 vccd1 vccd1 _15538_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15469_ _25815_/Q _15561_/B _15473_/S _15468_/X vssd1 vssd1 vccd1 vccd1 _15469_/X
+ sky130_fd_sc_hd__o211a_1
X_18257_ _18052_/X _18048_/X _18262_/S vssd1 vssd1 vccd1 vccd1 _18257_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17208_ _17222_/A _17208_/B vssd1 vssd1 vccd1 vccd1 _17209_/A sky130_fd_sc_hd__and2_1
X_18188_ _18685_/S vssd1 vssd1 vccd1 vccd1 _18898_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17139_ _20978_/A vssd1 vssd1 vccd1 vccd1 _18338_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20150_ _19725_/X _20149_/X _20015_/X vssd1 vssd1 vccd1 vccd1 _20154_/A sky130_fd_sc_hd__a21o_1
XFILLER_170_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20081_ _20081_/A _20081_/B vssd1 vssd1 vccd1 vccd1 _20081_/X sky130_fd_sc_hd__or2_1
XFILLER_258_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23840_ _23840_/A vssd1 vssd1 vccd1 vccd1 _26802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23771_ _23770_/X _26774_/Q _23780_/S vssd1 vssd1 vccd1 vccd1 _23772_/A sky130_fd_sc_hd__mux2_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20983_ _20983_/A vssd1 vssd1 vccd1 vccd1 _25863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25510_ _27014_/CLK _25510_/D vssd1 vssd1 vccd1 vccd1 _25510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22722_ _22722_/A vssd1 vssd1 vccd1 vccd1 _26352_/D sky130_fd_sc_hd__clkbuf_1
X_26490_ _26520_/CLK _26490_/D vssd1 vssd1 vccd1 vccd1 _26490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_74_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27266_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_230_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25441_ _25441_/A vssd1 vssd1 vccd1 vccd1 _27315_/D sky130_fd_sc_hd__clkbuf_1
X_22653_ _23696_/A vssd1 vssd1 vccd1 vccd1 _22653_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21604_ _21544_/X _21602_/X _21603_/X vssd1 vssd1 vccd1 vccd1 _21604_/Y sky130_fd_sc_hd__o21ai_1
X_25372_ _27285_/Q _23757_/A _25376_/S vssd1 vssd1 vccd1 vccd1 _25373_/A sky130_fd_sc_hd__mux2_1
X_22584_ _26309_/Q _22591_/B vssd1 vssd1 vccd1 vccd1 _22584_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27111_ _27198_/CLK _27111_/D vssd1 vssd1 vccd1 vccd1 _27111_/Q sky130_fd_sc_hd__dfxtp_4
X_24323_ _26999_/Q _24326_/C _24314_/X vssd1 vssd1 vccd1 vccd1 _24323_/Y sky130_fd_sc_hd__a21oi_1
X_21535_ _21533_/X _21534_/X _21512_/X vssd1 vssd1 vccd1 vccd1 _21535_/X sky130_fd_sc_hd__a21o_1
XFILLER_138_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27042_ _27044_/CLK _27042_/D vssd1 vssd1 vccd1 vccd1 _27042_/Q sky130_fd_sc_hd__dfxtp_1
X_24254_ _26974_/Q _24252_/B _24253_/Y vssd1 vssd1 vccd1 vccd1 _26974_/D sky130_fd_sc_hd__o21a_1
XFILLER_181_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21466_ _21461_/Y _21465_/X _21425_/X vssd1 vssd1 vccd1 vccd1 _21466_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_175_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23205_ _26549_/Q _23130_/X _23205_/S vssd1 vssd1 vccd1 vccd1 _23206_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20417_ _19683_/X _20416_/X _19718_/X vssd1 vssd1 vccd1 vccd1 _20417_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24185_ _24188_/A _24191_/C vssd1 vssd1 vccd1 vccd1 _24185_/Y sky130_fd_sc_hd__nor2_1
X_21397_ _21354_/X _21355_/X _21396_/Y _21386_/X vssd1 vssd1 vccd1 vccd1 _21397_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_175_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23136_ _23609_/A vssd1 vssd1 vccd1 vccd1 _23136_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20348_ _22526_/A _20382_/C vssd1 vssd1 vccd1 vccd1 _20348_/Y sky130_fd_sc_hd__nand2_1
XFILLER_150_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23067_ _26497_/Q _23066_/X _23067_/S vssd1 vssd1 vccd1 vccd1 _23068_/A sky130_fd_sc_hd__mux2_1
XTAP_5401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20279_ _20279_/A vssd1 vssd1 vccd1 vccd1 _20279_/Y sky130_fd_sc_hd__inv_2
XTAP_5412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput201 localMemory_wb_adr_i[1] vssd1 vssd1 vccd1 vccd1 input201/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput212 localMemory_wb_adr_i[8] vssd1 vssd1 vccd1 vccd1 input212/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22018_ _22018_/A vssd1 vssd1 vccd1 vccd1 _22027_/S sky130_fd_sc_hd__buf_6
XTAP_5434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput223 localMemory_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input223/X sky130_fd_sc_hd__buf_6
Xinput234 localMemory_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 input234/X sky130_fd_sc_hd__buf_8
XTAP_5445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 localMemory_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input245/X sky130_fd_sc_hd__buf_6
XFILLER_88_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput256 manufacturerID[2] vssd1 vssd1 vccd1 vccd1 input256/X sky130_fd_sc_hd__clkbuf_2
XTAP_5467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_264_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput267 partID[12] vssd1 vssd1 vccd1 vccd1 input267/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26826_ _27309_/CLK _26826_/D vssd1 vssd1 vccd1 vccd1 _26826_/Q sky130_fd_sc_hd__dfxtp_1
X_14840_ _15653_/S vssd1 vssd1 vccd1 vccd1 _16053_/S sky130_fd_sc_hd__buf_4
Xinput278 partID[8] vssd1 vssd1 vccd1 vccd1 input278/X sky130_fd_sc_hd__clkbuf_1
XTAP_5489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ _14771_/A vssd1 vssd1 vccd1 vccd1 _14772_/A sky130_fd_sc_hd__buf_2
XFILLER_57_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26757_ _27304_/CLK _26757_/D vssd1 vssd1 vccd1 vccd1 _26757_/Q sky130_fd_sc_hd__dfxtp_1
X_23969_ _23969_/A vssd1 vssd1 vccd1 vccd1 _26859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13722_ _15141_/A _13718_/X _13721_/X _15039_/A vssd1 vssd1 vccd1 vccd1 _13722_/X
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_4_4_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_4_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
X_16510_ _16510_/A vssd1 vssd1 vccd1 vccd1 _16533_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_25708_ _26673_/CLK _25708_/D vssd1 vssd1 vccd1 vccd1 _25708_/Q sky130_fd_sc_hd__dfxtp_1
X_17490_ _26256_/Q _17454_/A _17461_/A _25984_/Q vssd1 vssd1 vccd1 vccd1 _17683_/B
+ sky130_fd_sc_hd__a22o_2
X_26688_ _26913_/CLK _26688_/D vssd1 vssd1 vccd1 vccd1 _26688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13653_ _13651_/X _13652_/X _13653_/S vssd1 vssd1 vccd1 vccd1 _13653_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16441_ _26123_/Q _26024_/Q _16441_/S vssd1 vssd1 vccd1 vccd1 _16441_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25639_ _26297_/CLK _25639_/D vssd1 vssd1 vccd1 vccd1 _25639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16372_ _16372_/A _19273_/A vssd1 vssd1 vccd1 vccd1 _17846_/C sky130_fd_sc_hd__nor2_1
X_19160_ _18936_/A _18600_/X _18601_/Y _18597_/X _19159_/X vssd1 vssd1 vccd1 vccd1
+ _19160_/X sky130_fd_sc_hd__o221a_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ _13890_/A vssd1 vssd1 vccd1 vccd1 _13585_/A sky130_fd_sc_hd__buf_4
XFILLER_9_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _18161_/A _18161_/B _18111_/C vssd1 vssd1 vccd1 vccd1 _18293_/A sky130_fd_sc_hd__nor3_2
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _26930_/Q _16186_/S vssd1 vssd1 vccd1 vccd1 _15323_/X sky130_fd_sc_hd__or2_1
X_27309_ _27309_/CLK _27309_/D vssd1 vssd1 vccd1 vccd1 _27309_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19091_ _27089_/Q _18508_/A _18509_/A _27187_/Q _18510_/A vssd1 vssd1 vccd1 vccd1
+ _19091_/X sky130_fd_sc_hd__a221o_1
XFILLER_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18042_ _17876_/X _17869_/X _18042_/S vssd1 vssd1 vccd1 vccd1 _18042_/X sky130_fd_sc_hd__mux2_2
X_15254_ _16386_/S _15251_/X _15253_/X _14649_/A vssd1 vssd1 vccd1 vccd1 _15254_/X
+ sky130_fd_sc_hd__a211o_1
X_14205_ _26656_/Q _25696_/Q _15858_/S vssd1 vssd1 vccd1 vccd1 _14205_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15185_ _15044_/X _15183_/X _15184_/X vssd1 vssd1 vccd1 vccd1 _15186_/B sky130_fd_sc_hd__o21ai_1
X_14136_ input110/X input145/X _14240_/S vssd1 vssd1 vccd1 vccd1 _14136_/X sky130_fd_sc_hd__mux2_8
XFILLER_152_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19993_ _20295_/B vssd1 vssd1 vccd1 vccd1 _19993_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14067_ _25584_/Q vssd1 vssd1 vccd1 vccd1 _14067_/X sky130_fd_sc_hd__clkbuf_2
X_18944_ _18738_/X _18936_/X _18940_/Y _18943_/X vssd1 vssd1 vccd1 vccd1 _18944_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13018_ _14514_/S vssd1 vssd1 vccd1 vccd1 _14169_/B sky130_fd_sc_hd__buf_2
XFILLER_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18875_ _25515_/Q _18810_/X _18872_/X _18874_/X _18832_/X vssd1 vssd1 vccd1 vccd1
+ _18875_/X sky130_fd_sc_hd__o221a_1
XFILLER_140_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17826_ _17826_/A _15788_/B vssd1 vssd1 vccd1 vccd1 _17826_/X sky130_fd_sc_hd__or2b_1
XFILLER_39_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17757_ _18116_/B _18161_/C vssd1 vssd1 vccd1 vccd1 _18238_/A sky130_fd_sc_hd__nor2_2
X_14969_ _14967_/X _14968_/X _14969_/S vssd1 vssd1 vccd1 vccd1 _14969_/X sky130_fd_sc_hd__mux2_1
XFILLER_223_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16708_ _16708_/A _18251_/A vssd1 vssd1 vccd1 vccd1 _18230_/B sky130_fd_sc_hd__xnor2_4
XFILLER_208_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17688_ _17688_/A vssd1 vssd1 vccd1 vccd1 _18436_/A sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_320 _19616_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_331 _19624_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_342 _19609_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19427_ _18213_/X _18734_/X _19427_/S vssd1 vssd1 vccd1 vccd1 _19427_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_353 _19612_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16639_ _16639_/A _16639_/B vssd1 vssd1 vccd1 vccd1 _16639_/Y sky130_fd_sc_hd__nor2_1
XFILLER_211_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_364 input235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_375 _16994_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_386 _17022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19358_ _19358_/A _19358_/B vssd1 vssd1 vccd1 vccd1 _19358_/Y sky130_fd_sc_hd__nor2_1
XINSDIODE2_397 _17034_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18309_ _18324_/A _18213_/X _18308_/Y _18861_/A vssd1 vssd1 vccd1 vccd1 _18309_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_176_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19289_ _19318_/B _19289_/B vssd1 vssd1 vccd1 vccd1 _19289_/X sky130_fd_sc_hd__or2_1
XFILLER_176_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21320_ _21320_/A _21332_/B vssd1 vssd1 vccd1 vccd1 _21320_/X sky130_fd_sc_hd__or2_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21251_ _21251_/A vssd1 vssd1 vccd1 vccd1 _21346_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_192_wb_clk_i _26681_/CLK vssd1 vssd1 vccd1 vccd1 _27257_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_209_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20202_ _20173_/A _20173_/B _20201_/Y vssd1 vssd1 vccd1 vccd1 _20202_/X sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_121_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25553_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21182_ _21188_/A _21182_/B vssd1 vssd1 vccd1 vccd1 _21183_/A sky130_fd_sc_hd__or2_1
XFILLER_171_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20133_ _27150_/Q _27084_/Q vssd1 vssd1 vccd1 vccd1 _20134_/B sky130_fd_sc_hd__or2_1
X_25990_ _27000_/CLK _25990_/D vssd1 vssd1 vccd1 vccd1 _25990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_277_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24941_ _24941_/A vssd1 vssd1 vccd1 vccd1 _24941_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20064_ _19879_/X _20063_/Y _19926_/X vssd1 vssd1 vccd1 vccd1 _20067_/B sky130_fd_sc_hd__a21oi_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_13 _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_24 _19144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24872_ _24869_/Y _24870_/X _24871_/X vssd1 vssd1 vccd1 vccd1 _27124_/D sky130_fd_sc_hd__a21oi_1
XFILLER_273_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_35 _19381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_46 _20630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_57 _21718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_68 _20666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26611_ _26611_/CLK _26611_/D vssd1 vssd1 vccd1 vccd1 _26611_/Q sky130_fd_sc_hd__dfxtp_1
X_23823_ _23845_/A vssd1 vssd1 vccd1 vccd1 _23832_/S sky130_fd_sc_hd__buf_4
XFILLER_245_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_79 _20699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26542_ _27317_/CLK _26542_/D vssd1 vssd1 vccd1 vccd1 _26542_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23754_ _23754_/A vssd1 vssd1 vccd1 vccd1 _23754_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20966_ _20966_/A vssd1 vssd1 vccd1 vccd1 _25858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22705_ _26347_/Q _22704_/X _22705_/S vssd1 vssd1 vccd1 vccd1 _22706_/A sky130_fd_sc_hd__mux2_1
X_26473_ _27280_/CLK _26473_/D vssd1 vssd1 vccd1 vccd1 _26473_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23685_ _24004_/A _23860_/A vssd1 vssd1 vccd1 vccd1 _23767_/A sky130_fd_sc_hd__or2_4
X_20897_ _23712_/A vssd1 vssd1 vccd1 vccd1 _20897_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_213_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25424_ _23728_/X _27308_/Q _25426_/S vssd1 vssd1 vccd1 vccd1 _25425_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22636_ _22633_/A _26224_/Q _22632_/B vssd1 vssd1 vccd1 vccd1 _22636_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25355_ _25355_/A vssd1 vssd1 vccd1 vccd1 _27277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22567_ _22567_/A vssd1 vssd1 vccd1 vccd1 _22567_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_194_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24306_ _26993_/Q _24309_/C _24271_/X vssd1 vssd1 vccd1 vccd1 _24306_/Y sky130_fd_sc_hd__a21oi_1
X_21518_ _21581_/A vssd1 vssd1 vccd1 vccd1 _21518_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25286_ _25286_/A vssd1 vssd1 vccd1 vccd1 _27246_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22498_ _22498_/A _22502_/B vssd1 vssd1 vccd1 vccd1 _22499_/A sky130_fd_sc_hd__and2_1
XFILLER_6_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27025_ _27058_/CLK _27025_/D vssd1 vssd1 vccd1 vccd1 _27025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24237_ _24237_/A _24237_/B vssd1 vssd1 vccd1 vccd1 _24237_/Y sky130_fd_sc_hd__nor2_1
X_21449_ input49/X input84/X _21489_/S vssd1 vssd1 vccd1 vccd1 _21450_/A sky130_fd_sc_hd__mux2_8
XFILLER_182_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24168_ _26946_/Q _24169_/C _26947_/Q vssd1 vssd1 vccd1 vccd1 _24170_/B sky130_fd_sc_hd__a21oi_1
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23119_ _26513_/Q _23117_/X _23131_/S vssd1 vssd1 vccd1 vccd1 _23120_/A sky130_fd_sc_hd__mux2_1
X_24099_ _24099_/A vssd1 vssd1 vccd1 vccd1 _26917_/D sky130_fd_sc_hd__clkbuf_1
X_16990_ _16990_/A vssd1 vssd1 vccd1 vccd1 _16990_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15941_ _15491_/A _26341_/Q _26601_/Q _15501_/A _15939_/A vssd1 vssd1 vccd1 vccd1
+ _15941_/X sky130_fd_sc_hd__a221o_1
XTAP_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18660_ _26951_/Q _18461_/X _18463_/X _26983_/Q vssd1 vssd1 vccd1 vccd1 _18660_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15872_ _12912_/A _15871_/Y _12929_/A vssd1 vssd1 vccd1 vccd1 _15872_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_264_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17611_ _17615_/A _17611_/B vssd1 vssd1 vccd1 vccd1 _25584_/D sky130_fd_sc_hd__nor2_1
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26809_ _26905_/CLK _26809_/D vssd1 vssd1 vccd1 vccd1 _26809_/Q sky130_fd_sc_hd__dfxtp_1
X_14823_ _14809_/X _14819_/X _17179_/A vssd1 vssd1 vccd1 vccd1 _14823_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_252_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18591_ _19290_/A vssd1 vssd1 vccd1 vccd1 _19354_/B sky130_fd_sc_hd__buf_2
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ _17504_/B _17529_/X _17540_/X _17541_/Y vssd1 vssd1 vccd1 vccd1 _17543_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_44_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14754_ _14754_/A vssd1 vssd1 vccd1 vccd1 _14755_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_91_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ _15895_/S vssd1 vssd1 vccd1 vccd1 _13706_/A sky130_fd_sc_hd__buf_6
XFILLER_232_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17473_ _25969_/Q _25970_/Q _17455_/X _17472_/X vssd1 vssd1 vccd1 vccd1 _17475_/C
+ sky130_fd_sc_hd__o31a_1
X_14685_ _26682_/Q _25722_/Q _14699_/S vssd1 vssd1 vccd1 vccd1 _14685_/X sky130_fd_sc_hd__mux2_1
XFILLER_233_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19212_ _18716_/X _19195_/X _19211_/X _19078_/X vssd1 vssd1 vccd1 vccd1 _19212_/X
+ sky130_fd_sc_hd__a22o_1
X_16424_ _15085_/X _16422_/X _16423_/X _14793_/A vssd1 vssd1 vccd1 vccd1 _16424_/X
+ sky130_fd_sc_hd__a211o_1
X_13636_ _19887_/A _13636_/B vssd1 vssd1 vccd1 vccd1 _13636_/Y sky130_fd_sc_hd__nand2_1
XFILLER_198_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19143_ _18912_/A _19141_/Y _18705_/X vssd1 vssd1 vccd1 vccd1 _19143_/X sky130_fd_sc_hd__o21ba_1
X_13567_ _15871_/A _13567_/B vssd1 vssd1 vccd1 vccd1 _13567_/Y sky130_fd_sc_hd__nand2_1
X_16355_ _26933_/Q _16441_/S vssd1 vssd1 vccd1 vccd1 _16355_/X sky130_fd_sc_hd__or2_1
XFILLER_200_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15306_ _26802_/Q _26446_/Q _16262_/S vssd1 vssd1 vccd1 vccd1 _15306_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16286_ _19192_/A vssd1 vssd1 vccd1 vccd1 _16288_/A sky130_fd_sc_hd__inv_2
X_19074_ _18554_/X _19072_/X _19073_/Y vssd1 vssd1 vccd1 vccd1 _19074_/Y sky130_fd_sc_hd__a21oi_1
X_13498_ _14076_/A vssd1 vssd1 vccd1 vccd1 _14542_/A sky130_fd_sc_hd__buf_2
XFILLER_8_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18025_ _18025_/A vssd1 vssd1 vccd1 vccd1 _25598_/D sky130_fd_sc_hd__clkbuf_2
X_15237_ _20687_/A _19231_/A _16284_/S vssd1 vssd1 vccd1 vccd1 _17781_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15168_ _15168_/A vssd1 vssd1 vccd1 vccd1 _15169_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14119_ _14107_/A _14116_/X _14118_/X _14111_/A vssd1 vssd1 vccd1 vccd1 _14119_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_119_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19976_ _19852_/A _19976_/B _19976_/C vssd1 vssd1 vccd1 vccd1 _19976_/Y sky130_fd_sc_hd__nand3b_1
X_15099_ _16348_/S vssd1 vssd1 vccd1 vccd1 _15120_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_99_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18927_ _18927_/A vssd1 vssd1 vccd1 vccd1 _18927_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18858_ _18416_/X _18414_/X _18858_/S vssd1 vssd1 vccd1 vccd1 _18858_/X sky130_fd_sc_hd__mux2_1
XFILLER_267_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17809_ _17809_/A _18059_/B vssd1 vssd1 vccd1 vccd1 _17975_/A sky130_fd_sc_hd__nand2_4
XFILLER_283_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18789_ _17995_/B _18720_/X _18784_/Y _18787_/Y _18788_/X vssd1 vssd1 vccd1 vccd1
+ _18789_/X sky130_fd_sc_hd__a221o_4
XFILLER_242_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20820_ _25806_/Q vssd1 vssd1 vccd1 vccd1 _20821_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_242_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20751_ _20751_/A vssd1 vssd1 vccd1 vccd1 _25772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_150 _19947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_161 _15292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_172 _14449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23470_ _23470_/A vssd1 vssd1 vccd1 vccd1 _26666_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_183 _19824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20682_ _26283_/Q _20673_/X _20681_/X _20671_/X vssd1 vssd1 vccd1 vccd1 _25746_/D
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_194 _19728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22421_ _26241_/Q _22430_/B vssd1 vssd1 vccd1 vccd1 _22421_/X sky130_fd_sc_hd__or2_1
XFILLER_210_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25140_ _22524_/A _24639_/A _25139_/X _19256_/B _12781_/X vssd1 vssd1 vccd1 vccd1
+ _25140_/X sky130_fd_sc_hd__a221o_1
X_22352_ _22335_/Y _22350_/X _22351_/X _22348_/X vssd1 vssd1 vccd1 vccd1 _26229_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_176_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21303_ _20635_/A _21278_/X _21279_/X _21302_/X vssd1 vssd1 vccd1 vccd1 _21303_/X
+ sky130_fd_sc_hd__o211a_1
X_25071_ _22496_/A _25065_/X _25060_/X _16635_/D _25052_/X vssd1 vssd1 vccd1 vccd1
+ _25071_/X sky130_fd_sc_hd__a221o_1
X_22283_ _26207_/Q _22269_/X _22282_/X _22273_/X vssd1 vssd1 vccd1 vccd1 _26207_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24022_ _26883_/Q _23533_/X _24026_/S vssd1 vssd1 vccd1 vccd1 _24023_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21234_ input43/X input68/X _21327_/S vssd1 vssd1 vccd1 vccd1 _21234_/X sky130_fd_sc_hd__mux2_8
XFILLER_163_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21165_ _21165_/A vssd1 vssd1 vccd1 vccd1 _25926_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20116_ _20666_/A _20355_/A _20093_/X _20357_/A _20095_/A vssd1 vssd1 vccd1 vccd1
+ _20118_/A sky130_fd_sc_hd__o221a_1
XFILLER_120_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25973_ _27058_/CLK _25973_/D vssd1 vssd1 vccd1 vccd1 _25973_/Q sky130_fd_sc_hd__dfxtp_4
X_21096_ _25907_/Q _21094_/X _21095_/X input37/X vssd1 vssd1 vccd1 vccd1 _21097_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24924_ _27139_/Q _24913_/X _24923_/Y _24921_/X vssd1 vssd1 vccd1 vccd1 _27139_/D
+ sky130_fd_sc_hd__o211a_1
X_20047_ _27147_/Q _27081_/Q vssd1 vssd1 vccd1 vccd1 _20047_/Y sky130_fd_sc_hd__nor2_1
XFILLER_274_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24855_ _24852_/Y _24853_/X _24854_/X vssd1 vssd1 vccd1 vccd1 _27119_/D sky130_fd_sc_hd__a21oi_1
XFILLER_283_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23806_ _23709_/X _26787_/Q _23810_/S vssd1 vssd1 vccd1 vccd1 _23807_/A sky130_fd_sc_hd__mux2_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24786_ _20626_/A _19642_/X _24645_/Y _24782_/X vssd1 vssd1 vccd1 vccd1 _24786_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21998_ _21998_/A vssd1 vssd1 vccd1 vccd1 _26111_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26525_ _26877_/CLK _26525_/D vssd1 vssd1 vccd1 vccd1 _26525_/Q sky130_fd_sc_hd__dfxtp_1
X_23737_ _23737_/A vssd1 vssd1 vccd1 vccd1 _26763_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20949_ _25853_/Q _20948_/X _20949_/S vssd1 vssd1 vccd1 vccd1 _20950_/A sky130_fd_sc_hd__mux2_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _13945_/A _14468_/X _14469_/X _25582_/Q vssd1 vssd1 vccd1 vccd1 _14470_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26456_ _27266_/CLK _26456_/D vssd1 vssd1 vccd1 vccd1 _26456_/Q sky130_fd_sc_hd__dfxtp_2
X_23668_ _23668_/A vssd1 vssd1 vccd1 vccd1 _26740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13421_ _27273_/Q _26466_/Q _13616_/S vssd1 vssd1 vccd1 vccd1 _13421_/X sky130_fd_sc_hd__mux2_1
X_22619_ _22606_/X _22618_/Y _22614_/X vssd1 vssd1 vccd1 vccd1 _26322_/D sky130_fd_sc_hd__a21oi_1
X_25407_ _23702_/X _27300_/Q _25415_/S vssd1 vssd1 vccd1 vccd1 _25408_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26387_ _26483_/CLK _26387_/D vssd1 vssd1 vccd1 vccd1 _26387_/Q sky130_fd_sc_hd__dfxtp_1
X_23599_ _23599_/A vssd1 vssd1 vccd1 vccd1 _26711_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16140_ _25818_/Q _16380_/B _16308_/S _16139_/X vssd1 vssd1 vccd1 vccd1 _16140_/X
+ sky130_fd_sc_hd__o211a_1
X_25338_ _25338_/A vssd1 vssd1 vccd1 vccd1 _27269_/D sky130_fd_sc_hd__clkbuf_1
X_13352_ _14054_/A vssd1 vssd1 vccd1 vccd1 _14389_/S sky130_fd_sc_hd__buf_2
XFILLER_10_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16071_ _16069_/X _16070_/X _16071_/S vssd1 vssd1 vccd1 vccd1 _16071_/X sky130_fd_sc_hd__mux2_1
X_13283_ _26075_/Q _25880_/Q _16277_/S vssd1 vssd1 vccd1 vccd1 _13283_/X sky130_fd_sc_hd__mux2_1
X_25269_ _23712_/X _27239_/Q _25271_/S vssd1 vssd1 vccd1 vccd1 _25270_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15022_ _16305_/A vssd1 vssd1 vccd1 vccd1 _16135_/B sky130_fd_sc_hd__buf_2
X_27008_ _27044_/CLK _27008_/D vssd1 vssd1 vccd1 vccd1 _27008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19830_ _19830_/A _19830_/B _19830_/C vssd1 vssd1 vccd1 vccd1 _19830_/Y sky130_fd_sc_hd__nand3_1
XFILLER_123_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19761_ _20276_/A vssd1 vssd1 vccd1 vccd1 _19761_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16973_ _16983_/A _16973_/B _16973_/C vssd1 vssd1 vccd1 vccd1 _16973_/X sky130_fd_sc_hd__and3_1
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18712_ _18712_/A _18712_/B _18711_/X vssd1 vssd1 vccd1 vccd1 _18712_/X sky130_fd_sc_hd__or3b_1
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15924_ _15924_/A _15924_/B vssd1 vssd1 vccd1 vccd1 _15924_/X sky130_fd_sc_hd__or2_1
XFILLER_7_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19692_ _19779_/A vssd1 vssd1 vccd1 vccd1 _20452_/A sky130_fd_sc_hd__buf_2
XFILLER_249_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 core_wb_ack_i vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_2
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18643_ _18643_/A vssd1 vssd1 vccd1 vccd1 _18686_/B sky130_fd_sc_hd__clkbuf_2
X_15855_ _15488_/X _26110_/Q _26011_/Q _15671_/S _15401_/A vssd1 vssd1 vccd1 vccd1
+ _15855_/X sky130_fd_sc_hd__a221o_1
XFILLER_225_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _14806_/A vssd1 vssd1 vccd1 vccd1 _14807_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_64_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18574_ _18574_/A vssd1 vssd1 vccd1 vccd1 _18574_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15786_ _16585_/A _20055_/A _15785_/Y vssd1 vssd1 vccd1 vccd1 _15788_/B sky130_fd_sc_hd__a21oi_2
XFILLER_217_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12998_ _14349_/S vssd1 vssd1 vccd1 vccd1 _13062_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17525_ _25794_/Q vssd1 vssd1 vccd1 vccd1 _17525_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_205_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14737_ _14891_/A vssd1 vssd1 vccd1 vccd1 _14905_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_233_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17456_ _17456_/A _17456_/B _17456_/C _21235_/A vssd1 vssd1 vccd1 vccd1 _21870_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_178_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14668_ _14846_/B vssd1 vssd1 vccd1 vccd1 _14963_/S sky130_fd_sc_hd__buf_2
XFILLER_220_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16407_ _12705_/A _16398_/X _16406_/X _14710_/A vssd1 vssd1 vccd1 vccd1 _16407_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13619_ _13585_/X _26105_/Q _26006_/Q _15800_/S _15970_/S vssd1 vssd1 vccd1 vccd1
+ _13619_/X sky130_fd_sc_hd__a221o_1
XFILLER_193_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17387_ _24291_/A vssd1 vssd1 vccd1 vccd1 _17428_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_220_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14599_ _14599_/A vssd1 vssd1 vccd1 vccd1 _14600_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19126_ _18936_/A _18641_/Y _18642_/Y _18899_/A vssd1 vssd1 vccd1 vccd1 _19126_/X
+ sky130_fd_sc_hd__o22a_1
X_16338_ _15111_/A _26901_/Q _26773_/Q _16361_/S _15210_/X vssd1 vssd1 vccd1 vccd1
+ _16338_/X sky130_fd_sc_hd__a221o_1
XFILLER_118_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19057_ _27218_/Q _19331_/B vssd1 vssd1 vccd1 vccd1 _19057_/X sky130_fd_sc_hd__and2_1
X_16269_ _14763_/A _16267_/X _16268_/X vssd1 vssd1 vccd1 vccd1 _16269_/X sky130_fd_sc_hd__o21a_1
XFILLER_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput302 _17000_/X vssd1 vssd1 vccd1 vccd1 addr1[8] sky130_fd_sc_hd__buf_2
X_18008_ _18008_/A vssd1 vssd1 vccd1 vccd1 _18552_/A sky130_fd_sc_hd__clkbuf_2
Xoutput313 _16754_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[17] sky130_fd_sc_hd__buf_2
Xoutput324 _16781_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[27] sky130_fd_sc_hd__buf_2
Xoutput335 _16858_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[10] sky130_fd_sc_hd__buf_2
Xoutput346 _16920_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[20] sky130_fd_sc_hd__buf_2
XFILLER_114_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput357 _16981_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[30] sky130_fd_sc_hd__buf_2
XFILLER_259_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput368 _16796_/Y vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[2] sky130_fd_sc_hd__buf_2
XFILLER_273_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput379 _17024_/X vssd1 vssd1 vccd1 vccd1 din0[12] sky130_fd_sc_hd__buf_2
XFILLER_113_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19959_ _19958_/Y _19933_/C _19933_/B vssd1 vssd1 vccd1 vccd1 _19959_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_141_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22970_ _22970_/A vssd1 vssd1 vccd1 vccd1 _26458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_256_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21921_ _21921_/A vssd1 vssd1 vccd1 vccd1 _26077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24640_ _25173_/A vssd1 vssd1 vccd1 vccd1 _24771_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21852_ _26054_/Q _20951_/X _21860_/S vssd1 vssd1 vccd1 vccd1 _21853_/A sky130_fd_sc_hd__mux2_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20803_ _20803_/A vssd1 vssd1 vccd1 vccd1 _25797_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24571_ _24610_/A vssd1 vssd1 vccd1 vccd1 _24582_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_169_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21783_ _20605_/X _26024_/Q _21787_/S vssd1 vssd1 vccd1 vccd1 _21784_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26310_ _26322_/CLK _26310_/D vssd1 vssd1 vccd1 vccd1 _26310_/Q sky130_fd_sc_hd__dfxtp_2
X_23522_ _23522_/A vssd1 vssd1 vccd1 vccd1 _26687_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20734_ _20734_/A vssd1 vssd1 vccd1 vccd1 _25764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27290_ _27322_/CLK _27290_/D vssd1 vssd1 vccd1 vccd1 _27290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26241_ _26248_/CLK _26241_/D vssd1 vssd1 vccd1 vccd1 _26241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23453_ _23453_/A vssd1 vssd1 vccd1 vccd1 _26658_/D sky130_fd_sc_hd__clkbuf_1
X_20665_ _26276_/Q _20660_/X _20664_/X _20658_/X vssd1 vssd1 vccd1 vccd1 _25739_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22404_ _22360_/C _22395_/B _22390_/B vssd1 vssd1 vccd1 vccd1 _22405_/B sky130_fd_sc_hd__a21o_1
XFILLER_149_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26172_ _26238_/CLK _26172_/D vssd1 vssd1 vccd1 vccd1 _26172_/Q sky130_fd_sc_hd__dfxtp_1
X_23384_ _26628_/Q _23063_/X _23386_/S vssd1 vssd1 vccd1 vccd1 _23385_/A sky130_fd_sc_hd__mux2_1
X_20596_ _23766_/A vssd1 vssd1 vccd1 vccd1 _20596_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25123_ _27188_/Q _25112_/X _25122_/X vssd1 vssd1 vccd1 vccd1 _27188_/D sky130_fd_sc_hd__o21ba_1
X_22335_ _22379_/A _22390_/B vssd1 vssd1 vccd1 vccd1 _22335_/Y sky130_fd_sc_hd__nand2_2
XFILLER_152_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25054_ _20648_/A _25031_/X _25053_/X vssd1 vssd1 vccd1 vccd1 _25054_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_279_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22266_ _26201_/Q _22254_/X _22265_/X _22258_/X vssd1 vssd1 vccd1 vccd1 _26201_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24005_ _24061_/A vssd1 vssd1 vccd1 vccd1 _24074_/S sky130_fd_sc_hd__buf_4
X_21217_ _25468_/Q _21247_/A vssd1 vssd1 vccd1 vccd1 _21217_/X sky130_fd_sc_hd__or2_1
XFILLER_151_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22197_ input1/X input267/X _22207_/S vssd1 vssd1 vccd1 vccd1 _22197_/X sky130_fd_sc_hd__mux2_1
XFILLER_278_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21148_ _21166_/A vssd1 vssd1 vccd1 vccd1 _21148_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_278_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25956_ _27000_/CLK _25956_/D vssd1 vssd1 vccd1 vccd1 _25956_/Q sky130_fd_sc_hd__dfxtp_1
X_13970_ _14054_/A vssd1 vssd1 vccd1 vccd1 _14391_/S sky130_fd_sc_hd__clkbuf_4
X_21079_ _21197_/A _21079_/B vssd1 vssd1 vccd1 vccd1 _21080_/A sky130_fd_sc_hd__or2_1
XFILLER_281_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12921_ input117/X input153/X _14240_/S vssd1 vssd1 vccd1 vccd1 _12922_/B sky130_fd_sc_hd__mux2_8
X_24907_ _24550_/A _24978_/B _24314_/X vssd1 vssd1 vccd1 vccd1 _24907_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25887_ _27281_/CLK _25887_/D vssd1 vssd1 vccd1 vccd1 _25887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15640_ _26796_/Q _26440_/Q _15643_/S vssd1 vssd1 vccd1 vccd1 _15640_/X sky130_fd_sc_hd__mux2_1
X_12852_ input113/X input148/X _25868_/Q vssd1 vssd1 vccd1 vccd1 _17592_/C sky130_fd_sc_hd__mux2_8
X_24838_ _20662_/A _24829_/X _24703_/Y _24830_/X vssd1 vssd1 vccd1 vccd1 _24838_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _15073_/A _23565_/A _15570_/X _15388_/A vssd1 vssd1 vccd1 vccd1 _16896_/A
+ sky130_fd_sc_hd__o211ai_4
X_12783_ _12783_/A vssd1 vssd1 vccd1 vccd1 _21195_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24769_ _27099_/Q _24701_/A _24768_/Y _24720_/A vssd1 vssd1 vccd1 vccd1 _24770_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _17308_/X _17312_/C _17309_/Y vssd1 vssd1 vccd1 vccd1 _25523_/D sky130_fd_sc_hd__o21a_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ _14516_/X _14521_/X _14522_/S vssd1 vssd1 vccd1 vccd1 _14523_/B sky130_fd_sc_hd__mux2_1
XFILLER_203_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26508_ _27315_/CLK _26508_/D vssd1 vssd1 vccd1 vccd1 _26508_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _25505_/Q _18807_/A _18808_/A _25537_/Q vssd1 vssd1 vccd1 vccd1 _18290_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _17242_/A _17242_/B _25503_/Q vssd1 vssd1 vccd1 vccd1 _17243_/B sky130_fd_sc_hd__a21oi_1
XFILLER_203_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14453_ _14453_/A vssd1 vssd1 vccd1 vccd1 _14453_/X sky130_fd_sc_hd__buf_2
X_26439_ _27281_/CLK _26439_/D vssd1 vssd1 vccd1 vccd1 _26439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13404_ _15816_/S vssd1 vssd1 vccd1 vccd1 _13589_/S sky130_fd_sc_hd__buf_2
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14384_ _14384_/A vssd1 vssd1 vccd1 vccd1 _14384_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17172_ _25483_/Q _17185_/B vssd1 vssd1 vccd1 vccd1 _17172_/X sky130_fd_sc_hd__or2_1
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13335_ _13335_/A _13335_/B vssd1 vssd1 vccd1 vccd1 _13335_/X sky130_fd_sc_hd__or2_1
X_16123_ _16124_/A _17842_/B vssd1 vssd1 vccd1 vccd1 _16125_/A sky130_fd_sc_hd__nor2_2
XFILLER_182_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13266_ _13266_/A vssd1 vssd1 vccd1 vccd1 _15331_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16054_ _27250_/Q _16073_/B vssd1 vssd1 vccd1 vccd1 _16054_/X sky130_fd_sc_hd__or2_1
XFILLER_142_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15005_ _26516_/Q _26388_/Q _15005_/S vssd1 vssd1 vccd1 vccd1 _15005_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13197_ _13197_/A vssd1 vssd1 vccd1 vccd1 _22817_/C sky130_fd_sc_hd__buf_2
XFILLER_97_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19813_ _27107_/Q _19722_/X _19761_/X _19812_/X vssd1 vssd1 vccd1 vccd1 _19813_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19744_ _19740_/X _19741_/Y _19762_/B _20248_/A vssd1 vssd1 vccd1 vccd1 _19745_/B
+ sky130_fd_sc_hd__o31a_1
X_16956_ _16956_/A vssd1 vssd1 vccd1 vccd1 _16956_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15907_ _13863_/A _15903_/X _15906_/X _13162_/A vssd1 vssd1 vccd1 vccd1 _15907_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19675_ _19675_/A _19675_/B vssd1 vssd1 vccd1 vccd1 _19675_/X sky130_fd_sc_hd__or2_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16887_ _16887_/A vssd1 vssd1 vccd1 vccd1 _16887_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_225_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18626_ _19196_/A _18626_/B _18626_/C vssd1 vssd1 vccd1 vccd1 _18626_/X sky130_fd_sc_hd__or3_2
XFILLER_266_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15838_ _15488_/X _26698_/Q _26826_/Q _15671_/S _15836_/A vssd1 vssd1 vccd1 vccd1
+ _15838_/X sky130_fd_sc_hd__a221o_1
XFILLER_225_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18557_ _18557_/A vssd1 vssd1 vccd1 vccd1 _18557_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_252_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15769_ _15769_/A _15769_/B vssd1 vssd1 vccd1 vccd1 _15769_/X sky130_fd_sc_hd__or2_1
XFILLER_75_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17508_ _18006_/C _17662_/A vssd1 vssd1 vccd1 vccd1 _18182_/B sky130_fd_sc_hd__nor2_4
XFILLER_162_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18488_ _17920_/X _18896_/B _18487_/X vssd1 vssd1 vccd1 vccd1 _18488_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17439_ _25563_/Q _17437_/B _17438_/Y vssd1 vssd1 vccd1 vccd1 _25563_/D sky130_fd_sc_hd__o21a_1
XFILLER_123_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20450_ _20450_/A _20450_/B _20450_/C vssd1 vssd1 vccd1 vccd1 _20452_/B sky130_fd_sc_hd__and3_1
XFILLER_119_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19109_ _19109_/A _19109_/B _19109_/C vssd1 vssd1 vccd1 vccd1 _19110_/B sky130_fd_sc_hd__nand3_1
XFILLER_146_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20381_ _19766_/X _20380_/Y _19780_/X vssd1 vssd1 vccd1 vccd1 _20385_/A sky130_fd_sc_hd__a21o_1
X_22120_ _26160_/Q _22110_/X _22119_/X _21878_/X vssd1 vssd1 vccd1 vccd1 _26160_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_99_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27264_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22051_ _26135_/Q _20894_/X _22055_/S vssd1 vssd1 vccd1 vccd1 _22052_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_28_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26843_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21002_ _25872_/Q _20881_/X _21004_/S vssd1 vssd1 vccd1 vccd1 _21003_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25810_ _27293_/CLK _25810_/D vssd1 vssd1 vccd1 vccd1 _25810_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_275_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26790_ _27276_/CLK _26790_/D vssd1 vssd1 vccd1 vccd1 _26790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25741_ _26282_/CLK _25741_/D vssd1 vssd1 vccd1 vccd1 _25741_/Q sky130_fd_sc_hd__dfxtp_4
X_22953_ _22953_/A vssd1 vssd1 vccd1 vccd1 _26451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_284_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21904_ _21904_/A vssd1 vssd1 vccd1 vccd1 _26069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22884_ _26421_/Q _22736_/X _22884_/S vssd1 vssd1 vccd1 vccd1 _22885_/A sky130_fd_sc_hd__mux2_1
X_25672_ _25673_/CLK _25672_/D vssd1 vssd1 vccd1 vccd1 _25672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24623_ _24978_/A _24629_/B vssd1 vssd1 vccd1 vccd1 _24623_/Y sky130_fd_sc_hd__nand2_1
X_21835_ _21835_/A vssd1 vssd1 vccd1 vccd1 _26046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24554_ _27039_/Q _24546_/X _24553_/Y _24551_/X vssd1 vssd1 vccd1 vccd1 _27039_/D
+ sky130_fd_sc_hd__o211a_1
X_21766_ _21766_/A vssd1 vssd1 vccd1 vccd1 _26016_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23505_ _23505_/A vssd1 vssd1 vccd1 vccd1 _26682_/D sky130_fd_sc_hd__clkbuf_1
X_20717_ _25249_/A _25249_/B _23860_/A vssd1 vssd1 vccd1 vccd1 _20774_/A sky130_fd_sc_hd__or3_4
X_27273_ _27277_/CLK _27273_/D vssd1 vssd1 vccd1 vccd1 _27273_/Q sky130_fd_sc_hd__dfxtp_1
X_24485_ _26314_/Q _24473_/X _24474_/X input228/X _24384_/X vssd1 vssd1 vccd1 vccd1
+ _24485_/X sky130_fd_sc_hd__a221o_2
X_21697_ _21697_/A vssd1 vssd1 vccd1 vccd1 _25987_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26224_ _26326_/CLK _26224_/D vssd1 vssd1 vccd1 vccd1 _26224_/Q sky130_fd_sc_hd__dfxtp_1
X_23436_ _24004_/A _25393_/A vssd1 vssd1 vccd1 vccd1 _23493_/A sky130_fd_sc_hd__nor2_4
X_20648_ _20648_/A _20656_/B vssd1 vssd1 vccd1 vccd1 _20648_/X sky130_fd_sc_hd__or2_1
XFILLER_11_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26155_ _26900_/CLK _26155_/D vssd1 vssd1 vccd1 vccd1 _26155_/Q sky130_fd_sc_hd__dfxtp_1
X_23367_ _26620_/Q _23034_/X _23375_/S vssd1 vssd1 vccd1 vccd1 _23368_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20579_ _23578_/A vssd1 vssd1 vccd1 vccd1 _23754_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_180_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13120_ _12772_/A _26403_/Q _15174_/A _13119_/X vssd1 vssd1 vccd1 vccd1 _13120_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22318_ _26217_/Q _22310_/X _22316_/X _26318_/Q _22317_/X vssd1 vssd1 vccd1 vccd1
+ _22318_/X sky130_fd_sc_hd__a221o_1
X_25106_ _25106_/A vssd1 vssd1 vccd1 vccd1 _25106_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26086_ _26610_/CLK _26086_/D vssd1 vssd1 vccd1 vccd1 _26086_/Q sky130_fd_sc_hd__dfxtp_1
X_23298_ _20500_/X _26590_/Q _23302_/S vssd1 vssd1 vccd1 vccd1 _23299_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13051_ _13051_/A vssd1 vssd1 vccd1 vccd1 _15168_/A sky130_fd_sc_hd__clkbuf_4
X_25037_ _27172_/Q _25030_/X _25036_/X vssd1 vssd1 vccd1 vccd1 _27172_/D sky130_fd_sc_hd__o21ba_1
X_22249_ _22249_/A vssd1 vssd1 vccd1 vccd1 _22249_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_180_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16810_ _16810_/A _16824_/B _16841_/B vssd1 vssd1 vccd1 vccd1 _16811_/A sky130_fd_sc_hd__and3_4
X_17790_ _17790_/A _15438_/B vssd1 vssd1 vccd1 vccd1 _19122_/A sky130_fd_sc_hd__or2b_1
X_26988_ _26996_/CLK _26988_/D vssd1 vssd1 vccd1 vccd1 _26988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16741_ _25673_/Q vssd1 vssd1 vccd1 vccd1 _22498_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_253_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13953_ _13941_/X _13951_/X _13952_/X _13939_/X vssd1 vssd1 vccd1 vccd1 _13954_/C
+ sky130_fd_sc_hd__o211a_1
X_25939_ _27154_/CLK _25939_/D vssd1 vssd1 vccd1 vccd1 _25939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12904_ _14834_/A _14834_/B _12904_/C vssd1 vssd1 vccd1 vccd1 _16409_/A sky130_fd_sc_hd__nor3_1
X_19460_ _18636_/X _19453_/X _19454_/X _19459_/X vssd1 vssd1 vccd1 vccd1 _19460_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16672_ _25989_/Q _25990_/Q _25991_/Q _25992_/Q vssd1 vssd1 vccd1 vccd1 _16673_/D
+ sky130_fd_sc_hd__or4_4
X_13884_ _13881_/X _13883_/X _13884_/S vssd1 vssd1 vccd1 vccd1 _13884_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18411_ _18630_/A _18411_/B vssd1 vssd1 vccd1 vccd1 _18412_/A sky130_fd_sc_hd__and2_1
XFILLER_62_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15623_ _26924_/Q _15623_/B vssd1 vssd1 vccd1 vccd1 _15623_/X sky130_fd_sc_hd__or2_1
X_12835_ _12862_/A _14131_/A vssd1 vssd1 vccd1 vccd1 _12835_/Y sky130_fd_sc_hd__nor2_1
X_19391_ _19049_/A _19389_/X _19390_/Y _18037_/X vssd1 vssd1 vccd1 vccd1 _19391_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _18342_/A vssd1 vssd1 vccd1 vccd1 _18495_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _26797_/Q _26441_/Q _15557_/S vssd1 vssd1 vccd1 vccd1 _15554_/X sky130_fd_sc_hd__mux2_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _13082_/A vssd1 vssd1 vccd1 vccd1 _12767_/A sky130_fd_sc_hd__buf_2
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14505_ _26064_/Q _25869_/Q _15902_/S vssd1 vssd1 vccd1 vccd1 _14505_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _18273_/A vssd1 vssd1 vccd1 vccd1 _18273_/Y sky130_fd_sc_hd__inv_2
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _25587_/Q vssd1 vssd1 vccd1 vccd1 _13121_/B sky130_fd_sc_hd__buf_2
X_15485_ _26638_/Q _26734_/Q _15485_/S vssd1 vssd1 vccd1 vccd1 _15486_/B sky130_fd_sc_hd__mux2_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17224_ _17224_/A _17224_/B vssd1 vssd1 vccd1 vccd1 _17224_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14436_ _26097_/Q _25998_/Q _14514_/S vssd1 vssd1 vccd1 vccd1 _14436_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput12 core_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_1
Xinput23 core_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_1
Xinput34 core_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17155_ _25479_/Q vssd1 vssd1 vccd1 vccd1 _22817_/A sky130_fd_sc_hd__buf_2
Xinput45 dout0[11] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_2
X_14367_ _26066_/Q _14289_/S _14366_/X _13644_/A vssd1 vssd1 vccd1 vccd1 _14367_/X
+ sky130_fd_sc_hd__o211a_1
Xinput56 dout0[21] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput67 dout0[31] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput78 dout0[41] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__clkbuf_1
X_16106_ _15676_/X _25848_/Q _26048_/Q _15674_/X _13281_/A vssd1 vssd1 vccd1 vccd1
+ _16106_/X sky130_fd_sc_hd__a221o_1
X_13318_ _15842_/S vssd1 vssd1 vccd1 vccd1 _15841_/S sky130_fd_sc_hd__buf_4
Xinput89 dout0[51] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_1
X_17086_ _17087_/A _26235_/Q _17086_/C vssd1 vssd1 vccd1 vccd1 _22230_/B sky130_fd_sc_hd__and3_1
X_14298_ _13484_/A _14296_/X _14297_/X _13939_/X vssd1 vssd1 vccd1 vccd1 _14299_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16037_ _16037_/A vssd1 vssd1 vccd1 vccd1 _16038_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_272_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13249_ _13249_/A vssd1 vssd1 vccd1 vccd1 _13250_/A sky130_fd_sc_hd__buf_2
XFILLER_257_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17988_ _17988_/A vssd1 vssd1 vccd1 vccd1 _17988_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_270_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19727_ _19727_/A vssd1 vssd1 vccd1 vccd1 _19727_/X sky130_fd_sc_hd__buf_2
XFILLER_284_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16939_ _16939_/A _16939_/B vssd1 vssd1 vccd1 vccd1 _16954_/A sky130_fd_sc_hd__nand2_1
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19658_ _19658_/A vssd1 vssd1 vccd1 vccd1 _19659_/A sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_146_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27173_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_281_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18609_ _25510_/Q _18439_/A _18441_/A _25542_/Q vssd1 vssd1 vccd1 vccd1 _18609_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19589_ _19589_/A _19589_/B vssd1 vssd1 vccd1 vccd1 _19887_/B sky130_fd_sc_hd__nor2_1
XFILLER_253_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21620_ _25497_/Q _21620_/B vssd1 vssd1 vccd1 vccd1 _21620_/X sky130_fd_sc_hd__or2_1
XFILLER_52_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21551_ _21544_/X _21550_/X _21537_/X vssd1 vssd1 vccd1 vccd1 _21551_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_179_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20502_ _20502_/A vssd1 vssd1 vccd1 vccd1 _25694_/D sky130_fd_sc_hd__clkbuf_1
X_24270_ _26980_/Q _24268_/B _24269_/Y vssd1 vssd1 vccd1 vccd1 _26980_/D sky130_fd_sc_hd__o21a_1
XFILLER_193_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21482_ _25486_/Q _21495_/B vssd1 vssd1 vccd1 vccd1 _21482_/X sky130_fd_sc_hd__or2_1
XFILLER_148_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23221_ _23221_/A vssd1 vssd1 vccd1 vccd1 _26555_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20433_ _20434_/A _20434_/B vssd1 vssd1 vccd1 vccd1 _20433_/X sky130_fd_sc_hd__or2_1
XFILLER_107_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23152_ _23209_/S vssd1 vssd1 vccd1 vccd1 _23161_/S sky130_fd_sc_hd__buf_6
XFILLER_107_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20364_ _27127_/Q _19691_/X _24765_/A vssd1 vssd1 vccd1 vccd1 _20364_/X sky130_fd_sc_hd__o21a_1
XFILLER_107_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22103_ _26159_/Q _20970_/X _22103_/S vssd1 vssd1 vccd1 vccd1 _22104_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23083_ _26502_/Q _23082_/X _23083_/S vssd1 vssd1 vccd1 vccd1 _23084_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20295_ _27156_/Q _20295_/B vssd1 vssd1 vccd1 vccd1 _20295_/X sky130_fd_sc_hd__and2_1
XFILLER_249_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26911_ _27269_/CLK _26911_/D vssd1 vssd1 vccd1 vccd1 _26911_/Q sky130_fd_sc_hd__dfxtp_1
X_22034_ _22090_/A vssd1 vssd1 vccd1 vccd1 _22103_/S sky130_fd_sc_hd__buf_8
XFILLER_0_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26842_ _27326_/CLK _26842_/D vssd1 vssd1 vccd1 vccd1 _26842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26773_ _26929_/CLK _26773_/D vssd1 vssd1 vccd1 vccd1 _26773_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23985_ _26867_/Q _23584_/X _23987_/S vssd1 vssd1 vccd1 vccd1 _23986_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25724_ _26264_/CLK _25724_/D vssd1 vssd1 vccd1 vccd1 _25724_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_228_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22936_ _22947_/A vssd1 vssd1 vccd1 vccd1 _22945_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_113_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25655_ _25660_/CLK _25655_/D vssd1 vssd1 vccd1 vccd1 _25655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22867_ _26413_/Q _22711_/X _22873_/S vssd1 vssd1 vccd1 vccd1 _22868_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24606_ _24619_/A vssd1 vssd1 vccd1 vccd1 _24606_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_21818_ _21864_/S vssd1 vssd1 vccd1 vccd1 _21827_/S sky130_fd_sc_hd__clkbuf_4
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25586_ _26684_/CLK _25586_/D vssd1 vssd1 vccd1 vccd1 _25586_/Q sky130_fd_sc_hd__dfxtp_2
X_22798_ _26383_/Q _22717_/X _22800_/S vssd1 vssd1 vccd1 vccd1 _22799_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27325_ _27326_/CLK _27325_/D vssd1 vssd1 vccd1 vccd1 _27325_/Q sky130_fd_sc_hd__dfxtp_1
X_21749_ _21749_/A vssd1 vssd1 vccd1 vccd1 _26008_/D sky130_fd_sc_hd__clkbuf_1
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24537_ _24772_/B vssd1 vssd1 vccd1 vccd1 _24629_/A sky130_fd_sc_hd__inv_2
XPHY_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15270_ _14622_/A _15254_/X _15260_/X _15269_/X _14683_/A vssd1 vssd1 vccd1 vccd1
+ _15270_/X sky130_fd_sc_hd__a311o_1
X_27256_ _27324_/CLK _27256_/D vssd1 vssd1 vccd1 vccd1 _27256_/Q sky130_fd_sc_hd__dfxtp_1
X_24468_ _24454_/X _25616_/Q _24467_/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__o21ai_4
XFILLER_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26207_ _26257_/CLK _26207_/D vssd1 vssd1 vccd1 vccd1 _26207_/Q sky130_fd_sc_hd__dfxtp_1
X_14221_ _26068_/Q _25873_/Q _14221_/S vssd1 vssd1 vccd1 vccd1 _14221_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23419_ _26644_/Q _23114_/X _23419_/S vssd1 vssd1 vccd1 vccd1 _23420_/A sky130_fd_sc_hd__mux2_1
X_24399_ _27010_/Q _24391_/X _24398_/Y _24379_/X vssd1 vssd1 vccd1 vccd1 _27010_/D
+ sky130_fd_sc_hd__o211a_1
X_27187_ _27196_/CLK _27187_/D vssd1 vssd1 vccd1 vccd1 _27187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14152_ _26656_/Q _25696_/Q _14497_/A vssd1 vssd1 vccd1 vccd1 _14152_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26138_ _26601_/CLK _26138_/D vssd1 vssd1 vccd1 vccd1 _26138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13103_ _13095_/X _13096_/X _15546_/S vssd1 vssd1 vccd1 vccd1 _13103_/X sky130_fd_sc_hd__mux2_2
X_14083_ _14153_/A _26881_/Q _26753_/Q _14518_/S _13610_/A vssd1 vssd1 vccd1 vccd1
+ _14083_/X sky130_fd_sc_hd__a221o_1
X_18960_ _18705_/X _18947_/Y _18959_/X _18010_/C vssd1 vssd1 vccd1 vccd1 _18960_/X
+ sky130_fd_sc_hd__o211a_2
X_26069_ _26593_/CLK _26069_/D vssd1 vssd1 vccd1 vccd1 _26069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13034_ _15714_/A vssd1 vssd1 vccd1 vccd1 _15725_/S sky130_fd_sc_hd__clkbuf_4
X_17911_ _17909_/X _17910_/X _18070_/S vssd1 vssd1 vccd1 vccd1 _17911_/X sky130_fd_sc_hd__mux2_1
X_18891_ _18891_/A vssd1 vssd1 vccd1 vccd1 _18891_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17842_ _16124_/A _17842_/B vssd1 vssd1 vccd1 vccd1 _17842_/X sky130_fd_sc_hd__and2b_1
XFILLER_67_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17773_ _18138_/B vssd1 vssd1 vccd1 vccd1 _18998_/A sky130_fd_sc_hd__buf_2
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14985_ _14747_/A _26712_/Q _26840_/Q _14811_/S _14773_/A vssd1 vssd1 vccd1 vccd1
+ _14985_/X sky130_fd_sc_hd__a221o_1
XFILLER_93_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19512_ _19512_/A vssd1 vssd1 vccd1 vccd1 _19512_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16724_ _22485_/A _16703_/X _16705_/X _18483_/A vssd1 vssd1 vccd1 vccd1 _16724_/X
+ sky130_fd_sc_hd__a22o_2
X_13936_ _26786_/Q _26430_/Q _14221_/S vssd1 vssd1 vccd1 vccd1 _13936_/X sky130_fd_sc_hd__mux2_1
XFILLER_208_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_502 _19583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19443_ _17673_/X _19441_/X _19442_/Y vssd1 vssd1 vccd1 vccd1 _19443_/Y sky130_fd_sc_hd__a21oi_1
XINSDIODE2_513 _17067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16655_ _20799_/B _16606_/Y _16638_/X _17514_/A _16654_/X vssd1 vssd1 vccd1 vccd1
+ _16676_/A sky130_fd_sc_hd__o32a_4
X_13867_ _26495_/Q _26367_/Q _14245_/S vssd1 vssd1 vccd1 vccd1 _13867_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_524 _17040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_535 _17049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_546 _25983_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15606_ _15606_/A vssd1 vssd1 vccd1 vccd1 _15606_/X sky130_fd_sc_hd__buf_6
XINSDIODE2_557 _26586_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12818_ _12959_/A vssd1 vssd1 vccd1 vccd1 _17224_/A sky130_fd_sc_hd__clkbuf_4
X_19374_ _19374_/A _19374_/B vssd1 vssd1 vccd1 vccd1 _19374_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16586_ _18079_/S _16586_/B vssd1 vssd1 vccd1 vccd1 _16962_/A sky130_fd_sc_hd__nand2_8
XFILLER_90_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13798_ _25732_/Q _15868_/B vssd1 vssd1 vccd1 vccd1 _13798_/X sky130_fd_sc_hd__or2_1
XFILLER_250_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18325_ _18325_/A _18325_/B vssd1 vssd1 vccd1 vccd1 _18327_/B sky130_fd_sc_hd__nor2_1
XFILLER_188_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15537_ _12772_/A _26409_/Q _15174_/A _15536_/X vssd1 vssd1 vccd1 vccd1 _15537_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _15044_/A vssd1 vssd1 vccd1 vccd1 _12750_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_231_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18256_ _18485_/A _17977_/X _18345_/S vssd1 vssd1 vccd1 vccd1 _18256_/X sky130_fd_sc_hd__mux2_1
X_15468_ _27249_/Q _15468_/B vssd1 vssd1 vccd1 vccd1 _15468_/X sky130_fd_sc_hd__or2_1
XFILLER_148_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17207_ _25495_/Q _17151_/X _17146_/A _17444_/A vssd1 vssd1 vccd1 vccd1 _17208_/B
+ sky130_fd_sc_hd__a22o_1
X_14419_ _13084_/A _26457_/Q _14001_/B _27264_/Q _14331_/X vssd1 vssd1 vccd1 vccd1
+ _14419_/X sky130_fd_sc_hd__o221a_1
XFILLER_147_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18187_ _19571_/C _18151_/B _19157_/S vssd1 vssd1 vccd1 vccd1 _18187_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15399_ _15399_/A _15399_/B vssd1 vssd1 vccd1 vccd1 _15399_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17138_ _17138_/A vssd1 vssd1 vccd1 vccd1 _25475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17069_ _25977_/Q _17061_/A _16998_/X _17015_/X vssd1 vssd1 vccd1 vccd1 _17069_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_170_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20080_ _20080_/A _20080_/B _20082_/A _20082_/B vssd1 vssd1 vccd1 vccd1 _20081_/B
+ sky130_fd_sc_hd__or4_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23770_ _23770_/A vssd1 vssd1 vccd1 vccd1 _23770_/X sky130_fd_sc_hd__buf_2
X_20982_ _26585_/Q _20986_/B _25867_/D vssd1 vssd1 vccd1 vccd1 _20983_/A sky130_fd_sc_hd__and3_1
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22721_ _26352_/Q _22720_/X _22721_/S vssd1 vssd1 vccd1 vccd1 _22722_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22652_ _22652_/A vssd1 vssd1 vccd1 vccd1 _26330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25440_ _23750_/X _27315_/Q _25448_/S vssd1 vssd1 vccd1 vccd1 _25441_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21603_ _21603_/A vssd1 vssd1 vccd1 vccd1 _21603_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22583_ _22580_/X _22582_/Y _22574_/X vssd1 vssd1 vccd1 vccd1 _26308_/D sky130_fd_sc_hd__a21oi_1
XFILLER_222_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25371_ _25371_/A vssd1 vssd1 vccd1 vccd1 _27284_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27110_ _27110_/CLK _27110_/D vssd1 vssd1 vccd1 vccd1 _27110_/Q sky130_fd_sc_hd__dfxtp_4
X_24322_ _26998_/Q _24320_/B _24321_/Y vssd1 vssd1 vccd1 vccd1 _26998_/D sky130_fd_sc_hd__o21a_1
XFILLER_221_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21534_ _21509_/X _19172_/X _21510_/X _25819_/Q _21483_/X vssd1 vssd1 vccd1 vccd1
+ _21534_/X sky130_fd_sc_hd__a221o_1
XFILLER_167_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24253_ _24269_/A _24258_/C vssd1 vssd1 vccd1 vccd1 _24253_/Y sky130_fd_sc_hd__nor2_1
X_27041_ _27044_/CLK _27041_/D vssd1 vssd1 vccd1 vccd1 _27041_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_43_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26797_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21465_ _21421_/X _21462_/X _21464_/Y _21451_/X vssd1 vssd1 vccd1 vccd1 _21465_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_5_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23204_ _23204_/A vssd1 vssd1 vccd1 vccd1 _26548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20416_ _27161_/Q _20415_/X _20461_/S vssd1 vssd1 vccd1 vccd1 _20416_/X sky130_fd_sc_hd__mux2_2
X_24184_ _26952_/Q _26951_/Q _24184_/C vssd1 vssd1 vccd1 vccd1 _24191_/C sky130_fd_sc_hd__and3_1
XFILLER_209_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21396_ _21396_/A vssd1 vssd1 vccd1 vccd1 _21396_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23135_ _23135_/A vssd1 vssd1 vccd1 vccd1 _26518_/D sky130_fd_sc_hd__clkbuf_1
X_20347_ _22524_/A _20225_/X _20338_/X _20345_/X _20346_/X vssd1 vssd1 vccd1 vccd1
+ _25685_/D sky130_fd_sc_hd__o221a_1
XFILLER_161_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23066_ _23539_/A vssd1 vssd1 vccd1 vccd1 _23066_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20278_ _20261_/A _20300_/C _20261_/B _20303_/B _20359_/A vssd1 vssd1 vccd1 vccd1
+ _20284_/A sky130_fd_sc_hd__o32a_1
XFILLER_68_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput202 localMemory_wb_adr_i[20] vssd1 vssd1 vccd1 vccd1 _17456_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22017_ _22017_/A vssd1 vssd1 vccd1 vccd1 _26120_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput213 localMemory_wb_adr_i[9] vssd1 vssd1 vccd1 vccd1 input213/X sky130_fd_sc_hd__clkbuf_1
XTAP_5435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput224 localMemory_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 input224/X sky130_fd_sc_hd__buf_6
XFILLER_76_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput235 localMemory_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 input235/X sky130_fd_sc_hd__buf_8
XFILLER_237_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput246 localMemory_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input246/X sky130_fd_sc_hd__buf_6
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput257 manufacturerID[3] vssd1 vssd1 vccd1 vccd1 input257/X sky130_fd_sc_hd__clkbuf_2
XTAP_5468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26825_ _26827_/CLK _26825_/D vssd1 vssd1 vccd1 vccd1 _26825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput268 partID[13] vssd1 vssd1 vccd1 vccd1 input268/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput279 partID[9] vssd1 vssd1 vccd1 vccd1 input279/X sky130_fd_sc_hd__clkbuf_1
XFILLER_276_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26756_ _26916_/CLK _26756_/D vssd1 vssd1 vccd1 vccd1 _26756_/Q sky130_fd_sc_hd__dfxtp_1
X_14770_ _14770_/A vssd1 vssd1 vccd1 vccd1 _14771_/A sky130_fd_sc_hd__buf_2
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23968_ _26859_/Q _23558_/X _23976_/S vssd1 vssd1 vccd1 vccd1 _23969_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25707_ _26531_/CLK _25707_/D vssd1 vssd1 vccd1 vccd1 _25707_/Q sky130_fd_sc_hd__dfxtp_1
X_13721_ _26072_/Q _15634_/S _13723_/A _13720_/X vssd1 vssd1 vccd1 vccd1 _13721_/X
+ sky130_fd_sc_hd__o211a_1
X_22919_ _26436_/Q _22682_/X _22923_/S vssd1 vssd1 vccd1 vccd1 _22920_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26687_ _26880_/CLK _26687_/D vssd1 vssd1 vccd1 vccd1 _26687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23899_ _23899_/A vssd1 vssd1 vccd1 vccd1 _26828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16440_ _26547_/Q _26155_/Q _16440_/S vssd1 vssd1 vccd1 vccd1 _16440_/X sky130_fd_sc_hd__mux2_1
X_25638_ _26250_/CLK _25638_/D vssd1 vssd1 vccd1 vccd1 _25638_/Q sky130_fd_sc_hd__dfxtp_1
X_13652_ _26917_/Q _26401_/Q _13652_/S vssd1 vssd1 vccd1 vccd1 _13652_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16371_ _17784_/A _17783_/A vssd1 vssd1 vccd1 vccd1 _19273_/A sky130_fd_sc_hd__nor2_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _14153_/A vssd1 vssd1 vccd1 vccd1 _13890_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_25569_ _25596_/CLK _25569_/D vssd1 vssd1 vccd1 vccd1 _25569_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18110_ _27070_/Q _19058_/A _19059_/A _27168_/Q vssd1 vssd1 vccd1 vccd1 _18110_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27308_ _27308_/CLK _27308_/D vssd1 vssd1 vccd1 vccd1 _27308_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _15322_/A vssd1 vssd1 vccd1 vccd1 _16186_/S sky130_fd_sc_hd__clkbuf_4
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19090_ _27219_/Q _19364_/B vssd1 vssd1 vccd1 vccd1 _19090_/X sky130_fd_sc_hd__and2_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18041_ _17870_/X _17890_/X _18044_/S vssd1 vssd1 vccd1 vccd1 _18041_/X sky130_fd_sc_hd__mux2_1
X_27239_ _27303_/CLK _27239_/D vssd1 vssd1 vccd1 vccd1 _27239_/Q sky130_fd_sc_hd__dfxtp_1
X_15253_ _15065_/X _26414_/Q _16397_/S _15252_/X vssd1 vssd1 vccd1 vccd1 _15253_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14204_ _14725_/A _14204_/B _14204_/C vssd1 vssd1 vccd1 vccd1 _14204_/X sky130_fd_sc_hd__or3_1
XFILLER_125_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15184_ _15167_/X _26708_/Q _26836_/Q _16223_/S _15048_/X vssd1 vssd1 vccd1 vccd1
+ _15184_/X sky130_fd_sc_hd__a221o_1
XFILLER_4_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14135_ _14237_/A _14237_/B _14237_/C _15345_/B vssd1 vssd1 vccd1 vccd1 _14135_/X
+ sky130_fd_sc_hd__or4_1
X_19992_ _20000_/A vssd1 vssd1 vccd1 vccd1 _20295_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14066_ _13250_/A _26689_/Q _26817_/Q _14544_/S _12731_/A vssd1 vssd1 vccd1 vccd1
+ _14066_/X sky130_fd_sc_hd__a221o_1
XFILLER_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18943_ _19049_/A _18941_/Y _18942_/Y _18636_/A vssd1 vssd1 vccd1 vccd1 _18943_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13017_ _14351_/S vssd1 vssd1 vccd1 vccd1 _14514_/S sky130_fd_sc_hd__buf_2
X_18874_ _17384_/X _18825_/X _18873_/X _18767_/X _18830_/X vssd1 vssd1 vccd1 vccd1
+ _18874_/X sky130_fd_sc_hd__a221o_1
XFILLER_95_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17825_ _17817_/D _17823_/Y _18724_/A vssd1 vssd1 vccd1 vccd1 _17825_/Y sky130_fd_sc_hd__a21oi_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__buf_2
XFILLER_95_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17756_ _18111_/C vssd1 vssd1 vccd1 vccd1 _18161_/C sky130_fd_sc_hd__clkbuf_2
X_14968_ _26516_/Q _26388_/Q _14970_/S vssd1 vssd1 vccd1 vccd1 _14968_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16707_ _16713_/A _16707_/B vssd1 vssd1 vccd1 vccd1 _18251_/A sky130_fd_sc_hd__nor2_2
XFILLER_223_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13919_ _13911_/A _17653_/B _13918_/X _12902_/X _25932_/Q vssd1 vssd1 vccd1 vccd1
+ _14606_/C sky130_fd_sc_hd__o32a_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17687_ _18172_/A vssd1 vssd1 vccd1 vccd1 _17688_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_310 _19620_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14899_ _15088_/S vssd1 vssd1 vccd1 vccd1 _15003_/S sky130_fd_sc_hd__buf_2
XFILLER_62_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_321 _19616_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_332 _19609_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19426_ _17853_/X _19423_/B _19425_/Y _18183_/X vssd1 vssd1 vccd1 vccd1 _19426_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_251_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_343 _19609_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16638_ _16638_/A _16638_/B _16762_/A _16638_/D vssd1 vssd1 vccd1 vccd1 _16638_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_223_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_354 _19612_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_365 input240/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_376 _16995_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_387 _17023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19357_ _19423_/B _19577_/C _18792_/A vssd1 vssd1 vccd1 vccd1 _19357_/X sky130_fd_sc_hd__a21o_1
XFILLER_204_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16569_ _19237_/A _16572_/B vssd1 vssd1 vccd1 vccd1 _16573_/A sky130_fd_sc_hd__and2_1
XFILLER_50_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_398 _17034_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18308_ _18324_/A _18308_/B vssd1 vssd1 vccd1 vccd1 _18308_/Y sky130_fd_sc_hd__nand2_1
XFILLER_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19288_ _19285_/Y _19286_/X _19287_/X _19185_/X vssd1 vssd1 vccd1 vccd1 _25623_/D
+ sky130_fd_sc_hd__o211a_1
X_18239_ _27136_/Q _18757_/A vssd1 vssd1 vccd1 vccd1 _18239_/X sky130_fd_sc_hd__or2_1
XFILLER_175_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21250_ _21285_/A vssd1 vssd1 vccd1 vccd1 _21587_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_144_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20201_ _20173_/A _20173_/B _20174_/A vssd1 vssd1 vccd1 vccd1 _20201_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_209_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21181_ _25931_/Q _21166_/X _21167_/X input31/X vssd1 vssd1 vccd1 vccd1 _21182_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20132_ _27150_/Q _27084_/Q vssd1 vssd1 vccd1 vccd1 _20134_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24940_ _27145_/Q _24927_/X _24939_/Y vssd1 vssd1 vccd1 vccd1 _27145_/D sky130_fd_sc_hd__o21a_1
X_20063_ _20082_/B _20063_/B vssd1 vssd1 vccd1 vccd1 _20063_/Y sky130_fd_sc_hd__xnor2_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_161_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27117_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_98_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_14 _18789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_25 _19144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_24871_ _24871_/A vssd1 vssd1 vccd1 vccd1 _24871_/X sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_36 _19381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_47 _20630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26610_ _26610_/CLK _26610_/D vssd1 vssd1 vccd1 vccd1 _26610_/Q sky130_fd_sc_hd__dfxtp_1
X_23822_ _23822_/A vssd1 vssd1 vccd1 vccd1 _26794_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_58 _21718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_69 _20668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26541_ _26673_/CLK _26541_/D vssd1 vssd1 vccd1 vccd1 _26541_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20965_ _25858_/Q _20964_/X _20965_/S vssd1 vssd1 vccd1 vccd1 _20966_/A sky130_fd_sc_hd__mux2_1
X_23753_ _23753_/A vssd1 vssd1 vccd1 vccd1 _26768_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22704_ _23747_/A vssd1 vssd1 vccd1 vccd1 _22704_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26472_ _26604_/CLK _26472_/D vssd1 vssd1 vccd1 vccd1 _26472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ _20896_/A vssd1 vssd1 vccd1 vccd1 _25836_/D sky130_fd_sc_hd__clkbuf_1
X_23684_ _23684_/A vssd1 vssd1 vccd1 vccd1 _23684_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_214_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25423_ _25423_/A vssd1 vssd1 vccd1 vccd1 _27307_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22635_ _22632_/X _22633_/X _22634_/X vssd1 vssd1 vccd1 vccd1 _26325_/D sky130_fd_sc_hd__a21oi_1
XFILLER_241_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25354_ _27277_/Q _23731_/A _25354_/S vssd1 vssd1 vccd1 vccd1 _25355_/A sky130_fd_sc_hd__mux2_1
X_22566_ _22553_/X _22565_/Y _22561_/X vssd1 vssd1 vccd1 vccd1 _26302_/D sky130_fd_sc_hd__a21oi_1
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24305_ _26992_/Q _24303_/B _24304_/Y vssd1 vssd1 vccd1 vccd1 _26992_/D sky130_fd_sc_hd__o21a_1
X_21517_ _21517_/A vssd1 vssd1 vccd1 vccd1 _21517_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25285_ _23734_/X _27246_/Q _25293_/S vssd1 vssd1 vccd1 vccd1 _25286_/A sky130_fd_sc_hd__mux2_1
X_22497_ _22497_/A vssd1 vssd1 vccd1 vccd1 _26273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27024_ _27058_/CLK _27024_/D vssd1 vssd1 vccd1 vccd1 _27024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24236_ _26969_/Q _24240_/C vssd1 vssd1 vccd1 vccd1 _24237_/B sky130_fd_sc_hd__and2_1
X_21448_ _21414_/X _21447_/X _21407_/X vssd1 vssd1 vccd1 vccd1 _21448_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_108_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24167_ _26946_/Q _24169_/C _24166_/Y vssd1 vssd1 vccd1 vccd1 _26946_/D sky130_fd_sc_hd__o21a_1
XFILLER_150_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21379_ _22817_/B _21416_/B vssd1 vssd1 vccd1 vccd1 _21379_/X sky130_fd_sc_hd__or2_1
XFILLER_269_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23118_ _23118_/A vssd1 vssd1 vccd1 vccd1 _23131_/S sky130_fd_sc_hd__buf_4
X_24098_ _26917_/Q _23539_/X _24098_/S vssd1 vssd1 vccd1 vccd1 _24099_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23049_ _23049_/A vssd1 vssd1 vccd1 vccd1 _26491_/D sky130_fd_sc_hd__clkbuf_1
X_15940_ _15486_/A _15937_/X _15939_/X _15311_/A vssd1 vssd1 vccd1 vccd1 _15940_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15871_ _15871_/A _15871_/B vssd1 vssd1 vccd1 vccd1 _15871_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ _14760_/X _17551_/X _17608_/X _17609_/X vssd1 vssd1 vccd1 vccd1 _17611_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_5298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14822_ _16350_/A vssd1 vssd1 vccd1 vccd1 _17179_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26808_ _26904_/CLK _26808_/D vssd1 vssd1 vccd1 vccd1 _26808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ _18650_/B _18590_/B vssd1 vssd1 vccd1 vccd1 _18590_/X sky130_fd_sc_hd__or2_2
XFILLER_92_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17541_ _17534_/X _17556_/B _14142_/X _17536_/X _25906_/Q vssd1 vssd1 vccd1 vccd1
+ _17541_/Y sky130_fd_sc_hd__o32ai_4
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26739_ _26739_/CLK _26739_/D vssd1 vssd1 vccd1 vccd1 _26739_/Q sky130_fd_sc_hd__dfxtp_1
X_14753_ _14753_/A vssd1 vssd1 vccd1 vccd1 _14754_/A sky130_fd_sc_hd__buf_2
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13704_ _13697_/X _13702_/X _14694_/A vssd1 vssd1 vccd1 vccd1 _13704_/X sky130_fd_sc_hd__o21a_1
XFILLER_233_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17472_ _26242_/Q _26241_/Q _17455_/X vssd1 vssd1 vccd1 vccd1 _17472_/X sky130_fd_sc_hd__or3b_4
XFILLER_204_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14684_ _17197_/A _14651_/X _14663_/X _14680_/X _14683_/X vssd1 vssd1 vccd1 vccd1
+ _14684_/X sky130_fd_sc_hd__a311o_1
XFILLER_60_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19211_ _19196_/X _19209_/Y _19210_/X _19187_/X _19076_/X vssd1 vssd1 vccd1 vccd1
+ _19211_/X sky130_fd_sc_hd__o32a_2
X_16423_ _15111_/X _26615_/Q _15221_/S _26355_/Q _15120_/S vssd1 vssd1 vccd1 vccd1
+ _16423_/X sky130_fd_sc_hd__o221a_1
XFILLER_32_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13635_ _25594_/Q vssd1 vssd1 vccd1 vccd1 _19887_/A sky130_fd_sc_hd__inv_6
XFILLER_204_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19142_ _18554_/X _19139_/X _19141_/Y vssd1 vssd1 vccd1 vccd1 _19142_/Y sky130_fd_sc_hd__a21oi_1
X_16354_ _27320_/Q _26577_/Q _16354_/S vssd1 vssd1 vccd1 vccd1 _16354_/X sky130_fd_sc_hd__mux2_1
X_13566_ _12892_/A _14133_/A _13565_/X _12915_/A _25919_/Q vssd1 vssd1 vccd1 vccd1
+ _13567_/B sky130_fd_sc_hd__o32a_2
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15305_ _14763_/A _15302_/X _15304_/X vssd1 vssd1 vccd1 vccd1 _15305_/X sky130_fd_sc_hd__o21a_1
X_19073_ _20168_/A _19268_/B vssd1 vssd1 vccd1 vccd1 _19073_/Y sky130_fd_sc_hd__nor2_1
XFILLER_185_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16285_ _17795_/A _16287_/B vssd1 vssd1 vccd1 vccd1 _19192_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13497_ _14725_/A _13497_/B _13497_/C vssd1 vssd1 vccd1 vccd1 _13497_/X sky130_fd_sc_hd__or3_1
XFILLER_8_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18024_ _18336_/A _18024_/B vssd1 vssd1 vccd1 vccd1 _18025_/A sky130_fd_sc_hd__and2_1
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15236_ _16204_/S vssd1 vssd1 vccd1 vccd1 _16284_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_60_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15167_ _15167_/A vssd1 vssd1 vccd1 vccd1 _15167_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14118_ _14153_/A _26397_/Q _13062_/A _14117_/X vssd1 vssd1 vccd1 vccd1 _14118_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_259_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19975_ _19977_/B _19950_/A vssd1 vssd1 vccd1 vccd1 _19982_/A sky130_fd_sc_hd__or2b_1
X_15098_ _16428_/S vssd1 vssd1 vccd1 vccd1 _15221_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14049_ _13337_/A _14046_/X _14048_/X _16006_/A vssd1 vssd1 vccd1 vccd1 _14049_/X
+ sky130_fd_sc_hd__a211o_1
X_18926_ _18340_/A _18932_/B _18925_/X vssd1 vssd1 vccd1 vccd1 _18926_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18857_ _18040_/X _18056_/X _18191_/X _18682_/A vssd1 vssd1 vccd1 vccd1 _18864_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17808_ _18079_/S _16586_/B _17871_/A _17807_/Y vssd1 vssd1 vccd1 vccd1 _18184_/B
+ sky130_fd_sc_hd__a22o_1
X_18788_ _18973_/A vssd1 vssd1 vccd1 vccd1 _18788_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17739_ _17703_/X _17739_/B _17739_/C vssd1 vssd1 vccd1 vccd1 _17740_/C sky130_fd_sc_hd__and3b_1
XFILLER_282_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20750_ _20550_/X _25772_/Q _20750_/S vssd1 vssd1 vccd1 vccd1 _20751_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_140 _16261_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_151 _19947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_162 _19912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19409_ _17673_/X _19407_/X _19408_/Y vssd1 vssd1 vccd1 vccd1 _19409_/Y sky130_fd_sc_hd__a21oi_1
XINSDIODE2_173 _14449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20681_ _20681_/A _20683_/B vssd1 vssd1 vccd1 vccd1 _20681_/X sky130_fd_sc_hd__or2_1
XINSDIODE2_184 _13921_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_195 _14240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22420_ _22460_/A vssd1 vssd1 vccd1 vccd1 _22430_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_148_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22351_ _22379_/A _22390_/B _26229_/Q vssd1 vssd1 vccd1 vccd1 _22351_/X sky130_fd_sc_hd__a21o_1
XFILLER_191_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21302_ _21300_/X _21301_/X _21290_/X vssd1 vssd1 vccd1 vccd1 _21302_/X sky130_fd_sc_hd__a21o_1
XFILLER_148_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25070_ _25124_/A vssd1 vssd1 vccd1 vccd1 _25070_/X sky130_fd_sc_hd__clkbuf_2
X_22282_ _26206_/Q _22279_/X _22270_/X _26307_/Q _22271_/X vssd1 vssd1 vccd1 vccd1
+ _22282_/X sky130_fd_sc_hd__a221o_1
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24021_ _24021_/A vssd1 vssd1 vccd1 vccd1 _26882_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21233_ _21356_/S vssd1 vssd1 vccd1 vccd1 _21327_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_105_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21164_ _21172_/A _21164_/B vssd1 vssd1 vccd1 vccd1 _21165_/A sky130_fd_sc_hd__or2_1
XFILLER_49_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20115_ _20115_/A vssd1 vssd1 vccd1 vccd1 _20357_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_252_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25972_ _27156_/CLK _25972_/D vssd1 vssd1 vccd1 vccd1 _25972_/Q sky130_fd_sc_hd__dfxtp_4
X_21095_ _21113_/A vssd1 vssd1 vccd1 vccd1 _21095_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_277_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24923_ _24923_/A _24923_/B vssd1 vssd1 vccd1 vccd1 _24923_/Y sky130_fd_sc_hd__nand2_1
X_20046_ _27147_/Q _27081_/Q vssd1 vssd1 vccd1 vccd1 _20046_/X sky130_fd_sc_hd__and2_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24854_ _24871_/A vssd1 vssd1 vccd1 vccd1 _24854_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23805_ _23805_/A vssd1 vssd1 vccd1 vccd1 _26786_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24785_ _27102_/Q _24798_/B vssd1 vssd1 vccd1 vccd1 _24785_/Y sky130_fd_sc_hd__nand2_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ _26111_/Q _20919_/X _22005_/S vssd1 vssd1 vccd1 vccd1 _21998_/A sky130_fd_sc_hd__mux2_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26524_ _26657_/CLK _26524_/D vssd1 vssd1 vccd1 vccd1 _26524_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23736_ _23734_/X _26763_/Q _23748_/S vssd1 vssd1 vccd1 vccd1 _23737_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ _23763_/A vssd1 vssd1 vccd1 vccd1 _20948_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26455_ _26913_/CLK _26455_/D vssd1 vssd1 vccd1 vccd1 _26455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23667_ _26740_/Q _23587_/X _23667_/S vssd1 vssd1 vccd1 vccd1 _23668_/A sky130_fd_sc_hd__mux2_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20879_ _25831_/Q _20878_/X _20885_/S vssd1 vssd1 vccd1 vccd1 _20880_/A sky130_fd_sc_hd__mux2_1
X_13420_ _26074_/Q _25879_/Q _13589_/S vssd1 vssd1 vccd1 vccd1 _13420_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25406_ _25463_/S vssd1 vssd1 vccd1 vccd1 _25415_/S sky130_fd_sc_hd__buf_2
X_22618_ _26322_/Q _22618_/B vssd1 vssd1 vccd1 vccd1 _22618_/Y sky130_fd_sc_hd__nand2_1
XFILLER_197_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26386_ _27292_/CLK _26386_/D vssd1 vssd1 vccd1 vccd1 _26386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23598_ _26711_/Q _23597_/X _23604_/S vssd1 vssd1 vccd1 vccd1 _23599_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25337_ _27269_/Q _23706_/A _25343_/S vssd1 vssd1 vccd1 vccd1 _25338_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13351_ _13351_/A vssd1 vssd1 vccd1 vccd1 _14741_/A sky130_fd_sc_hd__buf_4
X_22549_ _26296_/Q _22551_/B vssd1 vssd1 vccd1 vccd1 _22549_/Y sky130_fd_sc_hd__nand2_1
XFILLER_139_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16070_ _15063_/A _26703_/Q _26831_/Q _15634_/S vssd1 vssd1 vccd1 vccd1 _16070_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25268_ _25268_/A vssd1 vssd1 vccd1 vccd1 _27238_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13282_ _15662_/S vssd1 vssd1 vccd1 vccd1 _16277_/S sky130_fd_sc_hd__buf_6
XFILLER_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27007_ _27137_/CLK _27007_/D vssd1 vssd1 vccd1 vccd1 _27007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15021_ _14859_/X _15014_/X _15018_/X _15020_/X vssd1 vssd1 vccd1 vccd1 _15021_/X
+ sky130_fd_sc_hd__a211o_1
X_24219_ _26963_/Q _24221_/C _24218_/Y vssd1 vssd1 vccd1 vccd1 _26963_/D sky130_fd_sc_hd__o21a_1
XFILLER_108_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25199_ _25199_/A vssd1 vssd1 vccd1 vccd1 _25199_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19760_ _24706_/A vssd1 vssd1 vccd1 vccd1 _20276_/A sky130_fd_sc_hd__buf_6
X_16972_ _14886_/B _16952_/X _16887_/X vssd1 vssd1 vccd1 vccd1 _16975_/B sky130_fd_sc_hd__o21ai_2
XFILLER_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15923_ _25810_/Q _27244_/Q _15923_/S vssd1 vssd1 vccd1 vccd1 _15924_/B sky130_fd_sc_hd__mux2_1
X_18711_ _19482_/B _18704_/Y _18706_/X _18710_/Y _18027_/X vssd1 vssd1 vccd1 vccd1
+ _18711_/X sky130_fd_sc_hd__o32a_1
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19691_ _20100_/A vssd1 vssd1 vccd1 vccd1 _19691_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18642_ _18040_/X _18346_/X _18191_/X vssd1 vssd1 vccd1 vccd1 _18642_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_92_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15854_ _15488_/X _25843_/Q _26043_/Q _16087_/S _15836_/A vssd1 vssd1 vccd1 vccd1
+ _15854_/X sky130_fd_sc_hd__a221o_1
XFILLER_209_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14805_ _14755_/X _14798_/X _14799_/X _14804_/X vssd1 vssd1 vccd1 vccd1 _14805_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_264_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18573_ _17365_/X _18568_/X _18571_/X _18154_/A _18572_/X vssd1 vssd1 vccd1 vccd1
+ _18573_/X sky130_fd_sc_hd__a221o_1
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ _25739_/Q _16581_/A vssd1 vssd1 vccd1 vccd1 _15785_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12997_ _12992_/A _25586_/Q vssd1 vssd1 vccd1 vccd1 _14349_/S sky130_fd_sc_hd__and2b_2
XFILLER_206_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ _24335_/A vssd1 vssd1 vccd1 vccd1 _17548_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _16422_/S vssd1 vssd1 vccd1 vccd1 _14891_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ _17455_/A vssd1 vssd1 vccd1 vccd1 _17455_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14667_ _16387_/S vssd1 vssd1 vccd1 vccd1 _14846_/B sky130_fd_sc_hd__clkbuf_2
X_16406_ _16405_/A _16401_/X _16405_/Y _15187_/X vssd1 vssd1 vccd1 vccd1 _16406_/X
+ sky130_fd_sc_hd__o211a_1
X_13618_ _14495_/A vssd1 vssd1 vccd1 vccd1 _15970_/S sky130_fd_sc_hd__buf_2
X_17386_ _17384_/X _17389_/C _17385_/Y vssd1 vssd1 vccd1 vccd1 _25547_/D sky130_fd_sc_hd__o21a_1
X_14598_ _14602_/A _12868_/Y _12951_/X vssd1 vssd1 vccd1 vccd1 _14599_/A sky130_fd_sc_hd__a21o_1
XFILLER_220_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19125_ _16206_/Y _19192_/B _18366_/A _16207_/A _17503_/X vssd1 vssd1 vccd1 vccd1
+ _19125_/X sky130_fd_sc_hd__o221a_1
X_16337_ _26677_/Q _25717_/Q _16359_/S vssd1 vssd1 vccd1 vccd1 _16337_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13549_ _25734_/Q _16581_/A vssd1 vssd1 vccd1 vccd1 _13549_/X sky130_fd_sc_hd__or2_4
XFILLER_145_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19056_ _19056_/A vssd1 vssd1 vccd1 vccd1 _19056_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_195_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16268_ _13255_/X _26899_/Q _26771_/Q _16255_/S _14770_/A vssd1 vssd1 vccd1 vccd1
+ _16268_/X sky130_fd_sc_hd__a221o_1
X_18007_ _18010_/D vssd1 vssd1 vccd1 vccd1 _19218_/A sky130_fd_sc_hd__buf_2
Xoutput303 _27329_/X vssd1 vssd1 vccd1 vccd1 clk0 sky130_fd_sc_hd__clkbuf_1
X_15219_ _14744_/A _25782_/Q _15088_/S _26868_/Q _15120_/S vssd1 vssd1 vccd1 vccd1
+ _15219_/X sky130_fd_sc_hd__o221a_1
Xoutput314 _16758_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[18] sky130_fd_sc_hd__buf_2
X_16199_ _14801_/A _16195_/X _16198_/X _13314_/A vssd1 vssd1 vccd1 vccd1 _16199_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_273_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput325 _16701_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[2] sky130_fd_sc_hd__buf_2
Xoutput336 _16865_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[11] sky130_fd_sc_hd__buf_2
XFILLER_236_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput347 _16925_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[21] sky130_fd_sc_hd__buf_2
XFILLER_126_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput358 _16987_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[31] sky130_fd_sc_hd__buf_2
XFILLER_142_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput369 _16805_/X vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[3] sky130_fd_sc_hd__buf_2
XFILLER_113_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19958_ _27143_/Q _27077_/Q vssd1 vssd1 vccd1 vccd1 _19958_/Y sky130_fd_sc_hd__nor2_1
XFILLER_206_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18909_ _18738_/X _18899_/X _18903_/Y _18908_/X vssd1 vssd1 vccd1 vccd1 _18909_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_206_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19889_ _19889_/A _19980_/B vssd1 vssd1 vccd1 vccd1 _19889_/X sky130_fd_sc_hd__xor2_1
XFILLER_68_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21920_ _20546_/X _26077_/Q _21922_/S vssd1 vssd1 vccd1 vccd1 _21921_/A sky130_fd_sc_hd__mux2_1
XFILLER_255_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21851_ _21851_/A vssd1 vssd1 vccd1 vccd1 _21860_/S sky130_fd_sc_hd__buf_6
XFILLER_243_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20802_ _25797_/Q vssd1 vssd1 vccd1 vccd1 _20803_/A sky130_fd_sc_hd__clkbuf_1
X_24570_ _27044_/Q _24562_/X _24569_/Y _24567_/X vssd1 vssd1 vccd1 vccd1 _27044_/D
+ sky130_fd_sc_hd__o211a_1
X_21782_ _21782_/A vssd1 vssd1 vccd1 vccd1 _26023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23521_ _26687_/Q _23520_/X _23524_/S vssd1 vssd1 vccd1 vccd1 _23522_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20733_ _20517_/X _25764_/Q _20739_/S vssd1 vssd1 vccd1 vccd1 _20734_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26240_ _26240_/CLK _26240_/D vssd1 vssd1 vccd1 vccd1 _26240_/Q sky130_fd_sc_hd__dfxtp_1
X_23452_ _26658_/Q _23057_/X _23458_/S vssd1 vssd1 vccd1 vccd1 _23453_/A sky130_fd_sc_hd__mux2_1
X_20664_ _20664_/A _20670_/B vssd1 vssd1 vccd1 vccd1 _20664_/X sky130_fd_sc_hd__or2_1
XFILLER_196_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22403_ _22379_/X _22394_/A _22400_/Y _22401_/X _22402_/X vssd1 vssd1 vccd1 vccd1
+ _26238_/D sky130_fd_sc_hd__o221a_1
X_26171_ _26238_/CLK _26171_/D vssd1 vssd1 vccd1 vccd1 _26171_/Q sky130_fd_sc_hd__dfxtp_1
X_23383_ _23383_/A vssd1 vssd1 vccd1 vccd1 _26627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20595_ _23590_/A vssd1 vssd1 vccd1 vccd1 _23766_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25122_ _24732_/Y _25097_/X _25121_/Y _25109_/X vssd1 vssd1 vccd1 vccd1 _25122_/X
+ sky130_fd_sc_hd__a31o_1
X_22334_ _22337_/A vssd1 vssd1 vccd1 vccd1 _22379_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22265_ _26200_/Q _22264_/X _22255_/X _26301_/Q _22256_/X vssd1 vssd1 vccd1 vccd1
+ _22265_/X sky130_fd_sc_hd__a221o_1
X_25053_ _22489_/A _25038_/X _25033_/X _16732_/X _25052_/X vssd1 vssd1 vccd1 vccd1
+ _25053_/X sky130_fd_sc_hd__a221o_1
XFILLER_247_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21216_ _21219_/A _21219_/B _21221_/B _21208_/D vssd1 vssd1 vccd1 vccd1 _21247_/A
+ sky130_fd_sc_hd__or4b_1
X_24004_ _24004_/A _24004_/B vssd1 vssd1 vccd1 vccd1 _24061_/A sky130_fd_sc_hd__nor2_2
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22196_ _26183_/Q _22185_/X _22194_/X _22195_/X vssd1 vssd1 vccd1 vccd1 _26183_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_279_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21147_ _21147_/A vssd1 vssd1 vccd1 vccd1 _25921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25955_ _25992_/CLK _25955_/D vssd1 vssd1 vccd1 vccd1 _25955_/Q sky130_fd_sc_hd__dfxtp_1
X_21078_ _25902_/Q _21074_/X _21077_/X input10/X vssd1 vssd1 vccd1 vccd1 _21079_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_76_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12920_ _14320_/S vssd1 vssd1 vccd1 vccd1 _14240_/S sky130_fd_sc_hd__buf_4
X_24906_ _27133_/Q _24902_/X _24905_/Y vssd1 vssd1 vccd1 vccd1 _27133_/D sky130_fd_sc_hd__o21a_1
X_20029_ _22498_/A _19876_/X _20021_/X _20028_/X _19874_/X vssd1 vssd1 vccd1 vccd1
+ _25673_/D sky130_fd_sc_hd__o221a_1
XFILLER_74_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25886_ _27330_/A _25886_/D vssd1 vssd1 vccd1 vccd1 _25886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_274_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12851_ _25861_/Q _25791_/Q vssd1 vssd1 vccd1 vccd1 _12934_/A sky130_fd_sc_hd__nand2_2
X_24837_ _27115_/Q _24837_/B vssd1 vssd1 vccd1 vccd1 _24837_/Y sky130_fd_sc_hd__nand2_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _15553_/X _15569_/X _14590_/A vssd1 vssd1 vccd1 vccd1 _15570_/X sky130_fd_sc_hd__a21o_2
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _25935_/Q _25934_/Q vssd1 vssd1 vccd1 vccd1 _12783_/A sky130_fd_sc_hd__or2_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24768_ _24768_/A _24768_/B vssd1 vssd1 vccd1 vccd1 _24768_/Y sky130_fd_sc_hd__nand2_2
XFILLER_203_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14521_ _14517_/X _14518_/X _14519_/X _14520_/X _13048_/A _13630_/A vssd1 vssd1 vccd1
+ vccd1 _14521_/X sky130_fd_sc_hd__mux4_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26507_ _26796_/CLK _26507_/D vssd1 vssd1 vccd1 vccd1 _26507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23719_ _23786_/S vssd1 vssd1 vccd1 vccd1 _23732_/S sky130_fd_sc_hd__buf_6
XFILLER_159_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24699_ _24699_/A _24699_/B vssd1 vssd1 vccd1 vccd1 _27082_/D sky130_fd_sc_hd__nor2_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _24291_/A vssd1 vssd1 vccd1 vccd1 _17283_/A sky130_fd_sc_hd__buf_2
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26438_ _26467_/CLK _26438_/D vssd1 vssd1 vccd1 vccd1 _26438_/Q sky130_fd_sc_hd__dfxtp_2
X_14452_ _26489_/Q _26361_/Q _14452_/S vssd1 vssd1 vccd1 vccd1 _14452_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ _15904_/S vssd1 vssd1 vccd1 vccd1 _15816_/S sky130_fd_sc_hd__clkbuf_4
X_17171_ _17612_/A vssd1 vssd1 vccd1 vccd1 _17185_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_128_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26369_ _26465_/CLK _26369_/D vssd1 vssd1 vccd1 vccd1 _26369_/Q sky130_fd_sc_hd__dfxtp_2
X_14383_ _26782_/Q _26426_/Q _14553_/S vssd1 vssd1 vccd1 vccd1 _14383_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16122_ _25743_/Q _16121_/Y _16122_/S vssd1 vssd1 vccd1 vccd1 _17842_/B sky130_fd_sc_hd__mux2_2
XFILLER_128_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13334_ _25808_/Q _27242_/Q _15930_/S vssd1 vssd1 vccd1 vccd1 _13335_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16053_ _26863_/Q _25777_/Q _16053_/S vssd1 vssd1 vccd1 vccd1 _16053_/X sky130_fd_sc_hd__mux2_1
X_13265_ _13472_/A vssd1 vssd1 vccd1 vccd1 _13266_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15004_ _15002_/X _15003_/X _15004_/S vssd1 vssd1 vccd1 vccd1 _15004_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13196_ _13773_/A vssd1 vssd1 vccd1 vccd1 _13277_/A sky130_fd_sc_hd__clkbuf_4
X_19812_ _19793_/Y _19794_/X _20067_/A _19811_/Y vssd1 vssd1 vccd1 vccd1 _19812_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19743_ _20100_/A vssd1 vssd1 vccd1 vccd1 _20248_/A sky130_fd_sc_hd__clkbuf_2
X_16955_ _16983_/B _16955_/B vssd1 vssd1 vccd1 vccd1 _16956_/A sky130_fd_sc_hd__nor2_1
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15906_ _14107_/X _15904_/X _15905_/X _14111_/X vssd1 vssd1 vccd1 vccd1 _15906_/X
+ sky130_fd_sc_hd__a211o_1
X_19674_ _19675_/A _19675_/B vssd1 vssd1 vccd1 vccd1 _19674_/Y sky130_fd_sc_hd__nand2_1
X_16886_ _16886_/A vssd1 vssd1 vccd1 vccd1 _16886_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_265_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15837_ _16104_/A _15834_/X _15836_/X _15312_/A vssd1 vssd1 vccd1 vccd1 _15837_/X
+ sky130_fd_sc_hd__o211a_1
X_18625_ _18383_/A _18623_/X _18705_/A vssd1 vssd1 vccd1 vccd1 _18626_/C sky130_fd_sc_hd__o21ba_1
XFILLER_264_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18556_ _18556_/A vssd1 vssd1 vccd1 vccd1 _18556_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15768_ _26535_/Q _26143_/Q _15768_/S vssd1 vssd1 vccd1 vccd1 _15769_/B sky130_fd_sc_hd__mux2_1
XFILLER_280_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14719_ _16250_/A _14716_/X _14718_/X vssd1 vssd1 vccd1 vccd1 _14719_/Y sky130_fd_sc_hd__o21ai_1
X_17507_ _17679_/B vssd1 vssd1 vccd1 vccd1 _19583_/A sky130_fd_sc_hd__buf_4
X_18487_ _18487_/A _18487_/B vssd1 vssd1 vccd1 vccd1 _18487_/X sky130_fd_sc_hd__or2_1
X_15699_ _25740_/Q _15698_/Y _16122_/S vssd1 vssd1 vccd1 vccd1 _15701_/B sky130_fd_sc_hd__mux2_1
X_17438_ _24164_/A _17438_/B vssd1 vssd1 vccd1 vccd1 _17438_/Y sky130_fd_sc_hd__nor2_1
XFILLER_178_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17369_ _17365_/X _17370_/C _25542_/Q vssd1 vssd1 vccd1 vccd1 _17371_/B sky130_fd_sc_hd__a21oi_1
XFILLER_203_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19108_ _19109_/B _19109_/C _19109_/A vssd1 vssd1 vccd1 vccd1 _19122_/B sky130_fd_sc_hd__a21o_1
XFILLER_119_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20380_ _20380_/A _20398_/B vssd1 vssd1 vccd1 vccd1 _20380_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_107_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19039_ _19081_/B _19039_/B vssd1 vssd1 vccd1 vccd1 _19039_/X sky130_fd_sc_hd__or2_2
XFILLER_273_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22050_ _22050_/A vssd1 vssd1 vccd1 vccd1 _26134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21001_ _21001_/A vssd1 vssd1 vccd1 vccd1 _25871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_68_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26595_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_229_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25740_ _26282_/CLK _25740_/D vssd1 vssd1 vccd1 vccd1 _25740_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_233_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22952_ _26451_/Q _22730_/X _22956_/S vssd1 vssd1 vccd1 vccd1 _22953_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21903_ _20512_/X _26069_/Q _21911_/S vssd1 vssd1 vccd1 vccd1 _21904_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25671_ _27132_/CLK _25671_/D vssd1 vssd1 vccd1 vccd1 _25671_/Q sky130_fd_sc_hd__dfxtp_2
X_22883_ _22883_/A vssd1 vssd1 vccd1 vccd1 _26420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24622_ _27064_/Q _24615_/X _24621_/Y _24619_/X vssd1 vssd1 vccd1 vccd1 _27064_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_243_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21834_ _26046_/Q _20926_/X _21838_/S vssd1 vssd1 vccd1 vccd1 _21835_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24553_ _24553_/A _24553_/B vssd1 vssd1 vccd1 vccd1 _24553_/Y sky130_fd_sc_hd__nand2_1
XFILLER_169_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21765_ _20571_/X _26016_/Q _21765_/S vssd1 vssd1 vccd1 vccd1 _21766_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23504_ _26682_/Q _23133_/X _23506_/S vssd1 vssd1 vccd1 vccd1 _23505_/A sky130_fd_sc_hd__mux2_1
X_27272_ _27272_/CLK _27272_/D vssd1 vssd1 vccd1 vccd1 _27272_/Q sky130_fd_sc_hd__dfxtp_1
X_20716_ _25476_/Q _21793_/B vssd1 vssd1 vccd1 vccd1 _23860_/A sky130_fd_sc_hd__nand2_2
X_24484_ _27025_/Q _24480_/X _24483_/Y _24470_/X vssd1 vssd1 vccd1 vccd1 _27025_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21696_ _25987_/Q input199/X _21696_/S vssd1 vssd1 vccd1 vccd1 _21697_/A sky130_fd_sc_hd__mux2_1
X_26223_ _26326_/CLK _26223_/D vssd1 vssd1 vccd1 vccd1 _26223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23435_ _23435_/A vssd1 vssd1 vccd1 vccd1 _26651_/D sky130_fd_sc_hd__clkbuf_1
X_20647_ _20674_/A vssd1 vssd1 vccd1 vccd1 _20656_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26154_ _27292_/CLK _26154_/D vssd1 vssd1 vccd1 vccd1 _26154_/Q sky130_fd_sc_hd__dfxtp_1
X_23366_ _23434_/S vssd1 vssd1 vccd1 vccd1 _23375_/S sky130_fd_sc_hd__clkbuf_4
X_20578_ _20578_/A vssd1 vssd1 vccd1 vccd1 _25712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25105_ _27185_/Q _25085_/X _25104_/X vssd1 vssd1 vccd1 vccd1 _27185_/D sky130_fd_sc_hd__o21ba_1
X_22317_ _22317_/A vssd1 vssd1 vccd1 vccd1 _22317_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26085_ _26609_/CLK _26085_/D vssd1 vssd1 vccd1 vccd1 _26085_/Q sky130_fd_sc_hd__dfxtp_1
X_23297_ _23297_/A vssd1 vssd1 vccd1 vccd1 _26589_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13050_ _13050_/A vssd1 vssd1 vccd1 vccd1 _13051_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_152_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25036_ _24664_/Y _25014_/X _25035_/Y _25027_/X vssd1 vssd1 vccd1 vccd1 _25036_/X
+ sky130_fd_sc_hd__a31o_1
X_22248_ _26195_/Q _22235_/X _22247_/X _22243_/X vssd1 vssd1 vccd1 vccd1 _26195_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_274_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22179_ _22179_/A vssd1 vssd1 vccd1 vccd1 _22179_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_239_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26987_ _26987_/CLK _26987_/D vssd1 vssd1 vccd1 vccd1 _26987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16740_ _22496_/A _16726_/X _16727_/X _16635_/D vssd1 vssd1 vccd1 vccd1 _16740_/X
+ sky130_fd_sc_hd__a22o_1
X_13952_ _13937_/X _26102_/Q _26003_/Q _15759_/S _13943_/X vssd1 vssd1 vccd1 vccd1
+ _13952_/X sky130_fd_sc_hd__a221o_1
X_25938_ _27154_/CLK _25938_/D vssd1 vssd1 vccd1 vccd1 _25938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12903_ _13911_/A _17653_/B _12898_/X _12902_/X _25929_/Q vssd1 vssd1 vccd1 vccd1
+ _12904_/C sky130_fd_sc_hd__o32a_1
X_16671_ _25986_/Q _25987_/Q _25988_/Q _21562_/B vssd1 vssd1 vccd1 vccd1 _16673_/C
+ sky130_fd_sc_hd__o31a_4
X_25869_ _27265_/CLK _25869_/D vssd1 vssd1 vccd1 vccd1 _25869_/Q sky130_fd_sc_hd__dfxtp_1
X_13883_ _12768_/A _26691_/Q _26819_/Q _15890_/S vssd1 vssd1 vccd1 vccd1 _13883_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18410_ _14080_/X _18285_/X _18408_/X _18409_/X _25603_/Q vssd1 vssd1 vccd1 vccd1
+ _18411_/B sky130_fd_sc_hd__a32o_1
X_15622_ _27311_/Q _26568_/Q _16143_/S vssd1 vssd1 vccd1 vccd1 _15622_/X sky130_fd_sc_hd__mux2_1
X_12834_ _25598_/Q vssd1 vssd1 vccd1 vccd1 _14131_/A sky130_fd_sc_hd__clkbuf_2
X_19390_ _19389_/B _19389_/C _19392_/B vssd1 vssd1 vccd1 vccd1 _19390_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18341_ _18899_/A vssd1 vssd1 vccd1 vccd1 _18342_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15553_ _14621_/A _15539_/X _15543_/X _15552_/X _14681_/A vssd1 vssd1 vccd1 vccd1
+ _15553_/X sky130_fd_sc_hd__a311o_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _13582_/A vssd1 vssd1 vccd1 vccd1 _13082_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _13585_/A _26456_/Q _15726_/S _27263_/Q _13124_/A vssd1 vssd1 vccd1 vccd1
+ _14504_/X sky130_fd_sc_hd__o221a_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18272_ _18729_/A _18270_/X _18271_/X vssd1 vssd1 vccd1 vccd1 _18273_/A sky130_fd_sc_hd__o21ai_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15484_ _26670_/Q _25710_/Q _15484_/S vssd1 vssd1 vccd1 vccd1 _15484_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _13105_/B vssd1 vssd1 vccd1 vccd1 _17738_/B sky130_fd_sc_hd__buf_6
XFILLER_30_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17223_ _17223_/A vssd1 vssd1 vccd1 vccd1 _25499_/D sky130_fd_sc_hd__clkbuf_1
X_14435_ _14178_/S _14433_/X _14434_/X vssd1 vssd1 vccd1 vccd1 _14435_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 core_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17154_ _17154_/A vssd1 vssd1 vccd1 vccd1 _25478_/D sky130_fd_sc_hd__clkbuf_1
Xinput24 core_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_1
X_14366_ _25871_/Q _16419_/B vssd1 vssd1 vccd1 vccd1 _14366_/X sky130_fd_sc_hd__or2_1
Xinput35 core_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput46 dout0[12] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput57 dout0[22] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16105_ _15318_/A _16102_/X _16104_/X _15313_/A vssd1 vssd1 vccd1 vccd1 _16105_/X
+ sky130_fd_sc_hd__o211a_1
Xinput68 dout0[32] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_1
X_13317_ _13652_/S vssd1 vssd1 vccd1 vccd1 _15842_/S sky130_fd_sc_hd__buf_4
X_17085_ _17085_/A _17087_/C _17085_/C vssd1 vssd1 vccd1 vccd1 _17086_/C sky130_fd_sc_hd__and3_1
Xinput79 dout0[42] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__clkbuf_1
X_14297_ _13252_/A _26099_/Q _26000_/Q _16014_/S _13943_/X vssd1 vssd1 vccd1 vccd1
+ _14297_/X sky130_fd_sc_hd__a221o_1
X_16036_ _16633_/B _18726_/B _18735_/S vssd1 vssd1 vccd1 vccd1 _18838_/B sky130_fd_sc_hd__o21ai_4
X_13248_ _16261_/S vssd1 vssd1 vccd1 vccd1 _16348_/S sky130_fd_sc_hd__buf_4
XFILLER_108_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13179_ _13179_/A vssd1 vssd1 vccd1 vccd1 _13180_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17987_ _18364_/A vssd1 vssd1 vccd1 vccd1 _17988_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19726_ _25728_/Q vssd1 vssd1 vccd1 vccd1 _20635_/A sky130_fd_sc_hd__buf_6
XFILLER_78_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16938_ _16983_/B _16938_/B vssd1 vssd1 vccd1 vccd1 _16938_/X sky130_fd_sc_hd__or2_1
XFILLER_226_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19657_ _19676_/A vssd1 vssd1 vccd1 vccd1 _19657_/X sky130_fd_sc_hd__buf_2
XFILLER_226_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16869_ _16836_/X _16867_/X _16868_/X _16842_/X vssd1 vssd1 vccd1 vccd1 _16870_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_37_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18608_ _18741_/A vssd1 vssd1 vccd1 vccd1 _18608_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_252_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19588_ _19670_/A vssd1 vssd1 vccd1 vccd1 _19589_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_252_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18539_ _18539_/A _18539_/B _18539_/C _18539_/D vssd1 vssd1 vccd1 vccd1 _18540_/B
+ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_186_wb_clk_i _26681_/CLK vssd1 vssd1 vccd1 vccd1 _26453_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21550_ _20683_/A _21545_/X _21459_/A _21549_/X vssd1 vssd1 vccd1 vccd1 _21550_/X
+ sky130_fd_sc_hd__o211a_2
Xclkbuf_leaf_115_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26996_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_33_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20501_ _20500_/X _25694_/Q _20509_/S vssd1 vssd1 vccd1 vccd1 _20502_/A sky130_fd_sc_hd__mux2_1
X_21481_ _21545_/A vssd1 vssd1 vccd1 vccd1 _21481_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23220_ _26555_/Q _23047_/X _23222_/S vssd1 vssd1 vccd1 vccd1 _23221_/A sky130_fd_sc_hd__mux2_1
X_20432_ _27096_/Q vssd1 vssd1 vccd1 vccd1 _20434_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23151_ _23151_/A vssd1 vssd1 vccd1 vccd1 _26524_/D sky130_fd_sc_hd__clkbuf_1
X_20363_ _24641_/A vssd1 vssd1 vccd1 vccd1 _24765_/A sky130_fd_sc_hd__buf_6
XFILLER_146_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22102_ _22102_/A vssd1 vssd1 vccd1 vccd1 _26158_/D sky130_fd_sc_hd__clkbuf_1
X_23082_ _23555_/A vssd1 vssd1 vccd1 vccd1 _23082_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20294_ _20291_/Y _20292_/X _20268_/X _20271_/Y vssd1 vssd1 vccd1 vccd1 _20294_/X
+ sky130_fd_sc_hd__a211o_1
X_26910_ _27297_/CLK _26910_/D vssd1 vssd1 vccd1 vccd1 _26910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22033_ _23211_/A _23139_/A vssd1 vssd1 vccd1 vccd1 _22090_/A sky130_fd_sc_hd__nor2_4
XFILLER_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26841_ _26905_/CLK _26841_/D vssd1 vssd1 vccd1 vccd1 _26841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26772_ _26900_/CLK _26772_/D vssd1 vssd1 vccd1 vccd1 _26772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_263_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23984_ _23984_/A vssd1 vssd1 vccd1 vccd1 _26866_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25723_ _26843_/CLK _25723_/D vssd1 vssd1 vccd1 vccd1 _25723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22935_ _22935_/A vssd1 vssd1 vccd1 vccd1 _26443_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25654_ _25660_/CLK _25654_/D vssd1 vssd1 vccd1 vccd1 _25654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22866_ _22866_/A vssd1 vssd1 vccd1 vccd1 _26412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_271_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24605_ _24605_/A _24608_/B vssd1 vssd1 vccd1 vccd1 _24605_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21817_ _21817_/A vssd1 vssd1 vccd1 vccd1 _26038_/D sky130_fd_sc_hd__clkbuf_1
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25585_ _26684_/CLK _25585_/D vssd1 vssd1 vccd1 vccd1 _25585_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22797_ _22797_/A vssd1 vssd1 vccd1 vccd1 _26382_/D sky130_fd_sc_hd__clkbuf_1
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27324_ _27324_/CLK _27324_/D vssd1 vssd1 vccd1 vccd1 _27324_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24536_ _24472_/X _25629_/Q _24535_/X vssd1 vssd1 vccd1 vccd1 _24772_/B sky130_fd_sc_hd__o21a_4
XFILLER_169_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21748_ _20538_/X _26008_/Q _21754_/S vssd1 vssd1 vccd1 vccd1 _21749_/A sky130_fd_sc_hd__mux2_1
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27255_ _27319_/CLK _27255_/D vssd1 vssd1 vccd1 vccd1 _27255_/Q sky130_fd_sc_hd__dfxtp_1
X_24467_ _26311_/Q _24455_/X _24456_/X input224/X _24457_/X vssd1 vssd1 vccd1 vccd1
+ _24467_/X sky130_fd_sc_hd__a221o_1
XFILLER_157_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21679_ _25979_/Q input191/X _21685_/S vssd1 vssd1 vccd1 vccd1 _21680_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26206_ _26307_/CLK _26206_/D vssd1 vssd1 vccd1 vccd1 _26206_/Q sky130_fd_sc_hd__dfxtp_1
X_14220_ _15509_/A _14216_/X _14219_/X _14806_/A vssd1 vssd1 vccd1 vccd1 _14220_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_200_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23418_ _23418_/A vssd1 vssd1 vccd1 vccd1 _26643_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27186_ _27188_/CLK _27186_/D vssd1 vssd1 vccd1 vccd1 _27186_/Q sky130_fd_sc_hd__dfxtp_1
X_24398_ _24408_/A _24920_/A vssd1 vssd1 vccd1 vccd1 _24398_/Y sky130_fd_sc_hd__nand2_1
XFILLER_153_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26137_ _26595_/CLK _26137_/D vssd1 vssd1 vccd1 vccd1 _26137_/Q sky130_fd_sc_hd__dfxtp_2
X_14151_ _14433_/S vssd1 vssd1 vccd1 vccd1 _14497_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23349_ _20596_/X _26613_/Q _23357_/S vssd1 vssd1 vccd1 vccd1 _23350_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13102_ _13402_/A vssd1 vssd1 vccd1 vccd1 _15546_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_152_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26068_ _27269_/CLK _26068_/D vssd1 vssd1 vccd1 vccd1 _26068_/Q sky130_fd_sc_hd__dfxtp_1
X_14082_ _26657_/Q _25697_/Q _14433_/S vssd1 vssd1 vccd1 vccd1 _14082_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13033_ _14176_/S vssd1 vssd1 vccd1 vccd1 _15714_/A sky130_fd_sc_hd__clkbuf_4
X_17910_ _17821_/B _16206_/B _17954_/S vssd1 vssd1 vccd1 vccd1 _17910_/X sky130_fd_sc_hd__mux2_1
X_25019_ _27169_/Q _25000_/X _25018_/X vssd1 vssd1 vccd1 vccd1 _27169_/D sky130_fd_sc_hd__o21ba_1
XFILLER_106_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18890_ _19218_/A vssd1 vssd1 vccd1 vccd1 _18890_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17841_ _19011_/A _17839_/X _17840_/X vssd1 vssd1 vccd1 vccd1 _17841_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14984_ _26648_/Q _26744_/Q _14984_/S vssd1 vssd1 vccd1 vccd1 _14984_/X sky130_fd_sc_hd__mux2_1
X_17772_ _18076_/B _17772_/B vssd1 vssd1 vccd1 vccd1 _18138_/B sky130_fd_sc_hd__or2_1
XFILLER_219_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19511_ _19499_/X _18622_/X _19510_/X _19502_/X vssd1 vssd1 vccd1 vccd1 _25639_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_75_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13935_ _16639_/A _13932_/X _13934_/X vssd1 vssd1 vccd1 vccd1 _23530_/A sky130_fd_sc_hd__a21o_4
X_16723_ _17813_/A _16723_/B vssd1 vssd1 vccd1 vccd1 _18483_/A sky130_fd_sc_hd__xnor2_4
XFILLER_263_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16654_ _20798_/B _16654_/B _16654_/C _16654_/D vssd1 vssd1 vccd1 vccd1 _16654_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_35_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19442_ _19442_/A _19442_/B vssd1 vssd1 vccd1 vccd1 _19442_/Y sky130_fd_sc_hd__nor2_1
X_13866_ _26335_/Q _26595_/Q _14245_/S vssd1 vssd1 vccd1 vccd1 _13866_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_503 _25798_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_514 _17067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_525 _17040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15605_ _13284_/A _15602_/X _15604_/X _13762_/X vssd1 vssd1 vccd1 vccd1 _15610_/A
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_536 _17010_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12817_ _12822_/A vssd1 vssd1 vccd1 vccd1 _12959_/A sky130_fd_sc_hd__clkbuf_2
X_19373_ _18437_/A _19363_/X _19372_/X vssd1 vssd1 vccd1 vccd1 _19373_/X sky130_fd_sc_hd__a21o_4
XINSDIODE2_547 _20664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16585_ _16585_/A _18059_/B _17810_/B vssd1 vssd1 vccd1 vccd1 _18079_/S sky130_fd_sc_hd__nand3_4
XFILLER_222_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13797_ _13466_/X _23536_/A _13796_/X _13214_/A vssd1 vssd1 vccd1 vccd1 _19849_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15536_ _26925_/Q _16069_/S vssd1 vssd1 vccd1 vccd1 _15536_/X sky130_fd_sc_hd__or2_1
XFILLER_15_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18324_ _18324_/A _18324_/B vssd1 vssd1 vccd1 vccd1 _18327_/A sky130_fd_sc_hd__nor2_1
XFILLER_176_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _15376_/S vssd1 vssd1 vccd1 vccd1 _15044_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18255_ _18044_/X _18041_/X _18262_/S vssd1 vssd1 vccd1 vccd1 _18485_/A sky130_fd_sc_hd__mux2_1
X_15467_ _26862_/Q _25776_/Q _15467_/S vssd1 vssd1 vccd1 vccd1 _15467_/X sky130_fd_sc_hd__mux2_1
X_12679_ _25597_/Q vssd1 vssd1 vccd1 vccd1 _13001_/A sky130_fd_sc_hd__inv_2
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17206_ _19828_/A vssd1 vssd1 vccd1 vccd1 _17444_/A sky130_fd_sc_hd__buf_4
X_14418_ _12768_/A _26589_/Q _15890_/S _26329_/Q _13140_/A vssd1 vssd1 vccd1 vccd1
+ _14418_/X sky130_fd_sc_hd__o221a_1
XFILLER_147_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18186_ _18186_/A vssd1 vssd1 vccd1 vccd1 _19157_/S sky130_fd_sc_hd__buf_2
XFILLER_128_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15398_ _15227_/S _15396_/X _15397_/X _16185_/A vssd1 vssd1 vccd1 vccd1 _15399_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17137_ _17137_/A _17137_/B vssd1 vssd1 vccd1 vccd1 _17138_/A sky130_fd_sc_hd__and2_1
XFILLER_116_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14349_ _14347_/X _14348_/X _14349_/S vssd1 vssd1 vccd1 vccd1 _14349_/X sky130_fd_sc_hd__mux2_1
XFILLER_265_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17068_ _25976_/Q _17061_/A _16997_/X _17063_/X vssd1 vssd1 vccd1 vccd1 _17068_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16019_ _13346_/A _16017_/X _16018_/X _13976_/X vssd1 vssd1 vccd1 vccd1 _16019_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_170_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19709_ _19709_/A vssd1 vssd1 vccd1 vccd1 _20628_/A sky130_fd_sc_hd__buf_4
XFILLER_84_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20981_ _20981_/A vssd1 vssd1 vccd1 vccd1 _25862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22720_ _23763_/A vssd1 vssd1 vccd1 vccd1 _22720_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22651_ _26330_/Q _22650_/X _22657_/S vssd1 vssd1 vccd1 vccd1 _22652_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21602_ _20694_/A _21545_/X _21563_/X _21601_/X vssd1 vssd1 vccd1 vccd1 _21602_/X
+ sky130_fd_sc_hd__o211a_2
X_25370_ _27284_/Q _23754_/A _25376_/S vssd1 vssd1 vccd1 vccd1 _25371_/A sky130_fd_sc_hd__mux2_1
X_22582_ _26308_/Q _22591_/B vssd1 vssd1 vccd1 vccd1 _22582_/Y sky130_fd_sc_hd__nand2_1
XFILLER_179_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24321_ _24335_/A _24326_/C vssd1 vssd1 vccd1 vccd1 _24321_/Y sky130_fd_sc_hd__nor2_1
XFILLER_179_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21533_ _25490_/Q _21574_/B vssd1 vssd1 vccd1 vccd1 _21533_/X sky130_fd_sc_hd__or2_1
X_27040_ _27044_/CLK _27040_/D vssd1 vssd1 vccd1 vccd1 _27040_/Q sky130_fd_sc_hd__dfxtp_1
X_24252_ _26974_/Q _24252_/B vssd1 vssd1 vccd1 vccd1 _24258_/C sky130_fd_sc_hd__and2_1
XFILLER_182_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21464_ _21464_/A vssd1 vssd1 vccd1 vccd1 _21464_/Y sky130_fd_sc_hd__inv_2
XFILLER_239_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23203_ _26548_/Q _23127_/X _23205_/S vssd1 vssd1 vccd1 vccd1 _23204_/A sky130_fd_sc_hd__mux2_1
X_20415_ _20415_/A _20415_/B vssd1 vssd1 vccd1 vccd1 _20415_/X sky130_fd_sc_hd__xor2_1
X_24183_ _24183_/A _24183_/B vssd1 vssd1 vccd1 vccd1 _26951_/D sky130_fd_sc_hd__nor2_1
X_21395_ input45/X input80/X _21422_/S vssd1 vssd1 vccd1 vccd1 _21396_/A sky130_fd_sc_hd__mux2_8
XFILLER_135_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_83_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26877_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_161_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23134_ _26518_/Q _23133_/X _23137_/S vssd1 vssd1 vccd1 vccd1 _23135_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20346_ _22638_/B vssd1 vssd1 vccd1 vccd1 _20346_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_12_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26673_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23065_ _23065_/A vssd1 vssd1 vccd1 vccd1 _26496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20277_ _20277_/A vssd1 vssd1 vccd1 vccd1 _20359_/A sky130_fd_sc_hd__buf_2
XFILLER_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22016_ _26120_/Q _20948_/X _22016_/S vssd1 vssd1 vccd1 vccd1 _22017_/A sky130_fd_sc_hd__mux2_1
Xinput203 localMemory_wb_adr_i[21] vssd1 vssd1 vccd1 vccd1 _17456_/A sky130_fd_sc_hd__clkbuf_1
XTAP_5425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput214 localMemory_wb_cyc_i vssd1 vssd1 vccd1 vccd1 _21654_/C sky130_fd_sc_hd__clkbuf_1
XTAP_5436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput225 localMemory_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 input225/X sky130_fd_sc_hd__buf_6
Xinput236 localMemory_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 input236/X sky130_fd_sc_hd__buf_8
XTAP_5447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput247 localMemory_wb_sel_i[0] vssd1 vssd1 vccd1 vccd1 input247/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26824_ _27307_/CLK _26824_/D vssd1 vssd1 vccd1 vccd1 _26824_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput258 manufacturerID[4] vssd1 vssd1 vccd1 vccd1 input258/X sky130_fd_sc_hd__clkbuf_2
XTAP_5469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput269 partID[14] vssd1 vssd1 vccd1 vccd1 input269/X sky130_fd_sc_hd__clkbuf_2
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26755_ _27304_/CLK _26755_/D vssd1 vssd1 vccd1 vccd1 _26755_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23967_ _23989_/A vssd1 vssd1 vccd1 vccd1 _23976_/S sky130_fd_sc_hd__buf_2
XFILLER_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25706_ _27305_/CLK _25706_/D vssd1 vssd1 vccd1 vccd1 _25706_/Q sky130_fd_sc_hd__dfxtp_1
X_13720_ _25877_/Q _16061_/B vssd1 vssd1 vccd1 vccd1 _13720_/X sky130_fd_sc_hd__or2_1
X_22918_ _22918_/A vssd1 vssd1 vccd1 vccd1 _26435_/D sky130_fd_sc_hd__clkbuf_1
X_26686_ _26877_/CLK _26686_/D vssd1 vssd1 vccd1 vccd1 _26686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23898_ _23738_/X _26828_/Q _23904_/S vssd1 vssd1 vccd1 vccd1 _23899_/A sky130_fd_sc_hd__mux2_1
X_25637_ _26520_/CLK _25637_/D vssd1 vssd1 vccd1 vccd1 _25637_/Q sky130_fd_sc_hd__dfxtp_1
X_13651_ _27304_/Q _26561_/Q _13652_/S vssd1 vssd1 vccd1 vccd1 _13651_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22849_ _26405_/Q _22685_/X _22851_/S vssd1 vssd1 vccd1 vccd1 _22850_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16370_ _16370_/A vssd1 vssd1 vccd1 vccd1 _16372_/A sky130_fd_sc_hd__inv_2
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _13582_/A vssd1 vssd1 vccd1 vccd1 _14153_/A sky130_fd_sc_hd__clkbuf_4
X_25568_ _25596_/CLK _25568_/D vssd1 vssd1 vccd1 vccd1 _25568_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_185_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27307_ _27307_/CLK _27307_/D vssd1 vssd1 vccd1 vccd1 _27307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15321_ _15321_/A vssd1 vssd1 vccd1 vccd1 _15321_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_240_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24519_ _27032_/Q _24506_/X _24518_/Y _24499_/X vssd1 vssd1 vccd1 vccd1 _27032_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25499_ _26940_/CLK _25499_/D vssd1 vssd1 vccd1 vccd1 _25499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18040_ _18362_/A vssd1 vssd1 vccd1 vccd1 _18040_/X sky130_fd_sc_hd__clkbuf_2
X_27238_ _27238_/CLK _27238_/D vssd1 vssd1 vccd1 vccd1 _27238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15252_ _26930_/Q _16134_/S vssd1 vssd1 vccd1 vccd1 _15252_/X sky130_fd_sc_hd__or2_1
XFILLER_200_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14203_ _13941_/X _14201_/X _14202_/X _12754_/A vssd1 vssd1 vccd1 vccd1 _14204_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15183_ _26644_/Q _26740_/Q _16402_/S vssd1 vssd1 vccd1 vccd1 _15183_/X sky130_fd_sc_hd__mux2_1
X_27169_ _27173_/CLK _27169_/D vssd1 vssd1 vccd1 vccd1 _27169_/Q sky130_fd_sc_hd__dfxtp_1
X_14134_ _25922_/Q _14029_/B _14133_/Y _13748_/A vssd1 vssd1 vccd1 vccd1 _15345_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19991_ _24768_/A vssd1 vssd1 vccd1 vccd1 _19991_/X sky130_fd_sc_hd__buf_2
XFILLER_98_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14065_ _26625_/Q _26721_/Q _14459_/S vssd1 vssd1 vccd1 vccd1 _14065_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18942_ _18968_/B _18942_/B vssd1 vssd1 vccd1 vccd1 _18942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13016_ _14348_/S vssd1 vssd1 vccd1 vccd1 _14351_/S sky130_fd_sc_hd__clkbuf_2
X_18873_ _26955_/Q _18826_/X _18827_/X _26987_/Q vssd1 vssd1 vccd1 vccd1 _18873_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_239_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17824_ _17824_/A _17824_/B vssd1 vssd1 vccd1 vccd1 _18724_/A sky130_fd_sc_hd__and2_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__buf_2
XFILLER_282_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14967_ _26356_/Q _26616_/Q _14970_/S vssd1 vssd1 vccd1 vccd1 _14967_/X sky130_fd_sc_hd__mux2_1
X_17755_ _27069_/Q _18815_/A vssd1 vssd1 vccd1 vccd1 _17755_/X sky130_fd_sc_hd__or2b_4
XFILLER_282_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16706_ _16706_/A _16706_/B vssd1 vssd1 vccd1 vccd1 _16708_/A sky130_fd_sc_hd__nand2_2
X_13918_ input130/X input165/X _14488_/S vssd1 vssd1 vccd1 vccd1 _13918_/X sky130_fd_sc_hd__mux2_8
XINSDIODE2_300 _26464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17686_ _21203_/A _19552_/A _21283_/A vssd1 vssd1 vccd1 vccd1 _18172_/A sky130_fd_sc_hd__a21o_4
X_14898_ _16354_/S vssd1 vssd1 vccd1 vccd1 _15088_/S sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_311 _19620_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_322 _19616_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19425_ _19392_/B _19389_/B _19424_/X _16462_/A vssd1 vssd1 vccd1 vccd1 _19425_/Y
+ sky130_fd_sc_hd__o211ai_1
X_13849_ _13844_/X _13848_/X _13530_/X vssd1 vssd1 vccd1 vccd1 _13849_/Y sky130_fd_sc_hd__o21ai_4
XINSDIODE2_333 _19609_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16637_ _19046_/A _16637_/B _16637_/C _16637_/D vssd1 vssd1 vccd1 vccd1 _16638_/D
+ sky130_fd_sc_hd__or4_1
XINSDIODE2_344 _19609_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_355 _19612_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_366 _20487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19356_ _19356_/A _19356_/B vssd1 vssd1 vccd1 vccd1 _19577_/C sky130_fd_sc_hd__xor2_2
XINSDIODE2_377 _16997_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_388 _17024_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16568_ _19318_/B vssd1 vssd1 vccd1 vccd1 _16575_/C sky130_fd_sc_hd__inv_2
XFILLER_210_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_399 _17034_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18307_ _18307_/A vssd1 vssd1 vccd1 vccd1 _18738_/A sky130_fd_sc_hd__clkbuf_2
X_15519_ _15488_/A _26862_/Q _25776_/Q _15596_/S _15516_/A vssd1 vssd1 vccd1 vccd1
+ _15519_/X sky130_fd_sc_hd__a221o_1
XFILLER_149_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19287_ _25623_/Q _19287_/B vssd1 vssd1 vccd1 vccd1 _19287_/X sky130_fd_sc_hd__or2_1
X_16499_ _16497_/X _16498_/X _16499_/S vssd1 vssd1 vccd1 vccd1 _16499_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18238_ _18238_/A vssd1 vssd1 vccd1 vccd1 _19063_/A sky130_fd_sc_hd__buf_2
XFILLER_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18169_ _18460_/A vssd1 vssd1 vccd1 vccd1 _18826_/A sky130_fd_sc_hd__clkbuf_2
X_20200_ _20200_/A _20200_/B vssd1 vssd1 vccd1 vccd1 _20200_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21180_ _21180_/A vssd1 vssd1 vccd1 vccd1 _25930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20131_ _20131_/A _20131_/B vssd1 vssd1 vccd1 vccd1 _20135_/A sky130_fd_sc_hd__or2_1
XFILLER_116_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20062_ _20082_/A _20042_/B _20061_/X vssd1 vssd1 vccd1 vccd1 _20063_/B sky130_fd_sc_hd__o21ba_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_15 _18840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24870_ _20683_/A _19963_/X _24739_/Y _24779_/A vssd1 vssd1 vccd1 vccd1 _24870_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_85_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_26 _19150_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_37 _19433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23821_ _23731_/X _26794_/Q _23821_/S vssd1 vssd1 vccd1 vccd1 _23822_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_48 _20628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_59 _21718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26540_ _27283_/CLK _26540_/D vssd1 vssd1 vccd1 vccd1 _26540_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23752_ _23750_/X _26768_/Q _23764_/S vssd1 vssd1 vccd1 vccd1 _23753_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_130_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27156_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20964_ _23779_/A vssd1 vssd1 vccd1 vccd1 _20964_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22703_ _22703_/A vssd1 vssd1 vccd1 vccd1 _26346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26471_ _27278_/CLK _26471_/D vssd1 vssd1 vccd1 vccd1 _26471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23683_ _23683_/A vssd1 vssd1 vccd1 vccd1 _26747_/D sky130_fd_sc_hd__clkbuf_1
X_20895_ _25836_/Q _20894_/X _20901_/S vssd1 vssd1 vccd1 vccd1 _20896_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25422_ _23725_/X _27307_/Q _25426_/S vssd1 vssd1 vccd1 vccd1 _25423_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22634_ _24835_/A vssd1 vssd1 vccd1 vccd1 _22634_/X sky130_fd_sc_hd__buf_8
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25353_ _25353_/A vssd1 vssd1 vccd1 vccd1 _27276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22565_ _26302_/Q _22565_/B vssd1 vssd1 vccd1 vccd1 _22565_/Y sky130_fd_sc_hd__nand2_1
XFILLER_179_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24304_ _24312_/A _24309_/C vssd1 vssd1 vccd1 vccd1 _24304_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21516_ input55/X input90/X _21553_/S vssd1 vssd1 vccd1 vccd1 _21517_/A sky130_fd_sc_hd__mux2_8
XFILLER_182_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25284_ _25306_/A vssd1 vssd1 vccd1 vccd1 _25293_/S sky130_fd_sc_hd__buf_4
X_22496_ _22496_/A _22502_/B vssd1 vssd1 vccd1 vccd1 _22497_/A sky130_fd_sc_hd__and2_1
XFILLER_108_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27023_ _27058_/CLK _27023_/D vssd1 vssd1 vccd1 vccd1 _27023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24235_ _26968_/Q _24231_/B _24234_/Y vssd1 vssd1 vccd1 vccd1 _26968_/D sky130_fd_sc_hd__o21a_1
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21447_ _20664_/A _21415_/X _21350_/A _21446_/X vssd1 vssd1 vccd1 vccd1 _21447_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24166_ _26946_/Q _24169_/C _17414_/X vssd1 vssd1 vccd1 vccd1 _24166_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_135_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21378_ _21573_/A vssd1 vssd1 vccd1 vccd1 _21378_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_253_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23117_ _23590_/A vssd1 vssd1 vccd1 vccd1 _23117_/X sky130_fd_sc_hd__clkbuf_2
X_20329_ _19268_/A _18092_/A _19284_/X _20328_/X vssd1 vssd1 vccd1 vccd1 _20329_/Y
+ sky130_fd_sc_hd__a22oi_1
X_24097_ _24097_/A vssd1 vssd1 vccd1 vccd1 _26916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_268_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23048_ _26491_/Q _23047_/X _23051_/S vssd1 vssd1 vccd1 vccd1 _23049_/A sky130_fd_sc_hd__mux2_1
XTAP_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15870_ _17831_/A _16040_/B vssd1 vssd1 vccd1 vccd1 _16628_/B sky130_fd_sc_hd__nor2_2
XFILLER_88_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14821_ _16185_/A vssd1 vssd1 vccd1 vccd1 _16350_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_218_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26807_ _26900_/CLK _26807_/D vssd1 vssd1 vccd1 vccd1 _26807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24999_ _25142_/A vssd1 vssd1 vccd1 vccd1 _25159_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_218_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _15085_/A vssd1 vssd1 vccd1 vccd1 _14753_/A sky130_fd_sc_hd__clkbuf_2
X_17540_ _19636_/A vssd1 vssd1 vccd1 vccd1 _17540_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_217_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26738_ _27285_/CLK _26738_/D vssd1 vssd1 vccd1 vccd1 _26738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _13703_/A vssd1 vssd1 vccd1 vccd1 _14694_/A sky130_fd_sc_hd__buf_6
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17471_ _17471_/A _17701_/B _17694_/B _17470_/Y vssd1 vssd1 vccd1 vccd1 _21214_/A
+ sky130_fd_sc_hd__or4bb_1
XFILLER_189_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26669_ _26797_/CLK _26669_/D vssd1 vssd1 vccd1 vccd1 _26669_/Q sky130_fd_sc_hd__dfxtp_1
X_14683_ _14683_/A vssd1 vssd1 vccd1 vccd1 _14683_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_32_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19210_ _18666_/A _19208_/Y _17774_/X vssd1 vssd1 vccd1 vccd1 _19210_/X sky130_fd_sc_hd__o21a_1
X_13634_ _13010_/A _23539_/A _13633_/X _13028_/A vssd1 vssd1 vccd1 vccd1 _16846_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_32_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16422_ _26515_/Q _26387_/Q _16422_/S vssd1 vssd1 vccd1 vccd1 _16422_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16353_ _15085_/X _16351_/X _16352_/X _14802_/A vssd1 vssd1 vccd1 vccd1 _16353_/X
+ sky130_fd_sc_hd__a211o_1
X_19141_ _19141_/A _19472_/B vssd1 vssd1 vccd1 vccd1 _19141_/Y sky130_fd_sc_hd__nor2_1
X_13565_ input115/X input150/X _14033_/S vssd1 vssd1 vccd1 vccd1 _13565_/X sky130_fd_sc_hd__mux2_8
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15304_ _15110_/A _26706_/Q _26834_/Q _16086_/S _15210_/A vssd1 vssd1 vccd1 vccd1
+ _15304_/X sky130_fd_sc_hd__a221o_1
X_19072_ _18555_/X _19054_/X _19071_/X vssd1 vssd1 vccd1 vccd1 _19072_/X sky130_fd_sc_hd__a21o_4
XFILLER_158_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16284_ _25747_/Q _16283_/Y _16284_/S vssd1 vssd1 vccd1 vccd1 _16287_/B sky130_fd_sc_hd__mux2_2
X_13496_ _13485_/X _13487_/X _13495_/X _12755_/A vssd1 vssd1 vccd1 vccd1 _13497_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15235_ _14724_/X _15139_/Y _15234_/Y _14827_/X vssd1 vssd1 vccd1 vccd1 _19231_/A
+ sky130_fd_sc_hd__a211o_4
X_18023_ _18005_/X _18013_/X _18021_/X _18022_/X _14237_/B vssd1 vssd1 vccd1 vccd1
+ _18024_/B sky130_fd_sc_hd__a32o_1
XFILLER_145_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15166_ _26676_/Q _25716_/Q _16402_/S vssd1 vssd1 vccd1 vccd1 _15166_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14117_ _26913_/Q _14514_/S vssd1 vssd1 vccd1 vccd1 _14117_/X sky130_fd_sc_hd__or2_1
XFILLER_126_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19974_ _20006_/A _20006_/B vssd1 vssd1 vccd1 vccd1 _20080_/A sky130_fd_sc_hd__xnor2_1
X_15097_ _16341_/S vssd1 vssd1 vccd1 vccd1 _16428_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_259_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14048_ _13937_/A _26593_/Q _14369_/S _26333_/Q _14390_/S vssd1 vssd1 vccd1 vccd1
+ _14048_/X sky130_fd_sc_hd__o221a_1
X_18925_ _18705_/X _18912_/Y _18924_/X _18010_/C vssd1 vssd1 vccd1 vccd1 _18925_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18856_ _19354_/B _18905_/B _18855_/Y _18183_/X vssd1 vssd1 vccd1 vccd1 _18856_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_68_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17807_ _17807_/A vssd1 vssd1 vccd1 vccd1 _17807_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18787_ _19042_/A _18787_/B vssd1 vssd1 vccd1 vccd1 _18787_/Y sky130_fd_sc_hd__nand2_1
X_15999_ _15999_/A _15999_/B vssd1 vssd1 vccd1 vccd1 _15999_/X sky130_fd_sc_hd__or2_1
XFILLER_94_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17738_ _17738_/A _17738_/B vssd1 vssd1 vccd1 vccd1 _17739_/B sky130_fd_sc_hd__nand2_1
XFILLER_236_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_130 _16481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17669_ _17669_/A _17669_/B _17669_/C vssd1 vssd1 vccd1 vccd1 _17670_/C sky130_fd_sc_hd__or3_1
XFILLER_62_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_141 _16261_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_152 _23542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19408_ _19408_/A _19472_/B vssd1 vssd1 vccd1 vccd1 _19408_/Y sky130_fd_sc_hd__nor2_1
XFILLER_251_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_163 _13572_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20680_ _26282_/Q _20673_/X _20679_/X _20671_/X vssd1 vssd1 vccd1 vccd1 _25745_/D
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_174 _16419_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_185 _19800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_196 _14272_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19339_ _25528_/Q _18559_/X _19336_/X _19338_/X _18574_/X vssd1 vssd1 vccd1 vccd1
+ _19339_/X sky130_fd_sc_hd__o221a_1
XFILLER_176_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22350_ _17087_/A _26228_/Q _22350_/S vssd1 vssd1 vccd1 vccd1 _22350_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21301_ _21284_/X _18302_/X _21286_/X _25801_/Q _21641_/B vssd1 vssd1 vccd1 vccd1
+ _21301_/X sky130_fd_sc_hd__a221o_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22281_ _26206_/Q _22269_/X _22280_/X _22273_/X vssd1 vssd1 vccd1 vccd1 _26206_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24020_ _26882_/Q _23530_/X _24026_/S vssd1 vssd1 vccd1 vccd1 _24021_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21232_ _25866_/Q vssd1 vssd1 vccd1 vccd1 _21356_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21163_ _25926_/Q _21148_/X _21149_/X input26/X vssd1 vssd1 vccd1 vccd1 _21164_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20114_ _25740_/Q vssd1 vssd1 vccd1 vccd1 _20666_/A sky130_fd_sc_hd__buf_8
X_25971_ _27156_/CLK _25971_/D vssd1 vssd1 vccd1 vccd1 _25971_/Q sky130_fd_sc_hd__dfxtp_4
X_21094_ _21112_/A vssd1 vssd1 vccd1 vccd1 _21094_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24922_ _19790_/A _24913_/X _24920_/Y _24921_/X vssd1 vssd1 vccd1 vccd1 _27138_/D
+ sky130_fd_sc_hd__o211a_1
X_20045_ _27115_/Q _19877_/X _19967_/X _20044_/Y vssd1 vssd1 vccd1 vccd1 _20045_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_273_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24853_ _20670_/A _24848_/X _24719_/Y _24849_/X vssd1 vssd1 vccd1 vccd1 _24853_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23804_ _23706_/X _26786_/Q _23810_/S vssd1 vssd1 vccd1 vccd1 _23805_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24784_ _24780_/Y _24783_/X _22634_/X vssd1 vssd1 vccd1 vccd1 _27101_/D sky130_fd_sc_hd__a21oi_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21996_ _22018_/A vssd1 vssd1 vccd1 vccd1 _22005_/S sky130_fd_sc_hd__buf_4
XFILLER_226_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26523_ _26845_/CLK _26523_/D vssd1 vssd1 vccd1 vccd1 _26523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23735_ _23767_/A vssd1 vssd1 vccd1 vccd1 _23748_/S sky130_fd_sc_hd__buf_4
X_20947_ _20947_/A vssd1 vssd1 vccd1 vccd1 _25852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26454_ _27293_/CLK _26454_/D vssd1 vssd1 vccd1 vccd1 _26454_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23666_ _23666_/A vssd1 vssd1 vccd1 vccd1 _26739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20878_ _23693_/A vssd1 vssd1 vccd1 vccd1 _20878_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_197_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25405_ _25405_/A vssd1 vssd1 vccd1 vccd1 _27299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22617_ _22606_/X _22616_/Y _22614_/X vssd1 vssd1 vccd1 vccd1 _26321_/D sky130_fd_sc_hd__a21oi_1
X_26385_ _26580_/CLK _26385_/D vssd1 vssd1 vccd1 vccd1 _26385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23597_ _23597_/A vssd1 vssd1 vccd1 vccd1 _23597_/X sky130_fd_sc_hd__clkbuf_2
X_25336_ _25336_/A vssd1 vssd1 vccd1 vccd1 _27268_/D sky130_fd_sc_hd__clkbuf_1
X_13350_ _13488_/A vssd1 vssd1 vccd1 vccd1 _13351_/A sky130_fd_sc_hd__clkbuf_2
X_22548_ _22538_/X _22545_/Y _22547_/X vssd1 vssd1 vccd1 vccd1 _26295_/D sky130_fd_sc_hd__a21oi_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25267_ _23709_/X _27238_/Q _25271_/S vssd1 vssd1 vccd1 vccd1 _25268_/A sky130_fd_sc_hd__mux2_1
X_13281_ _13281_/A vssd1 vssd1 vccd1 vccd1 _15394_/A sky130_fd_sc_hd__buf_4
XFILLER_154_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22479_ _22479_/A vssd1 vssd1 vccd1 vccd1 _26265_/D sky130_fd_sc_hd__clkbuf_1
X_27006_ _27044_/CLK _27006_/D vssd1 vssd1 vccd1 vccd1 _27006_/Q sky130_fd_sc_hd__dfxtp_2
X_15020_ _15020_/A vssd1 vssd1 vccd1 vccd1 _15020_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24218_ _26963_/Q _24221_/C _24209_/X vssd1 vssd1 vccd1 vccd1 _24218_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25198_ _25198_/A vssd1 vssd1 vccd1 vccd1 _25198_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_146_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24149_ _17514_/C _24148_/X _22634_/X vssd1 vssd1 vccd1 vccd1 _26940_/D sky130_fd_sc_hd__a21oi_1
XFILLER_269_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16971_ _16971_/A vssd1 vssd1 vccd1 vccd1 _16971_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18710_ _18781_/B _18710_/B vssd1 vssd1 vccd1 vccd1 _18710_/Y sky130_fd_sc_hd__nand2_4
XFILLER_249_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15922_ _27308_/Q _26565_/Q _16110_/S vssd1 vssd1 vccd1 vccd1 _15922_/X sky130_fd_sc_hd__mux2_1
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19690_ _19687_/Y _27136_/Q _19820_/S vssd1 vssd1 vccd1 vccd1 _19690_/X sky130_fd_sc_hd__mux2_2
XFILLER_249_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18641_ _18547_/S _18363_/X _18640_/X vssd1 vssd1 vccd1 vccd1 _18641_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15853_ _13532_/X _15850_/X _15852_/X _15312_/A vssd1 vssd1 vccd1 vccd1 _15853_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14804_ _14804_/A vssd1 vssd1 vccd1 vccd1 _14804_/X sky130_fd_sc_hd__buf_2
X_18572_ _18572_/A vssd1 vssd1 vccd1 vccd1 _18572_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ _12996_/A vssd1 vssd1 vccd1 vccd1 _20868_/B sky130_fd_sc_hd__clkbuf_4
X_15784_ _13207_/A _23558_/A _15783_/Y vssd1 vssd1 vccd1 vccd1 _20055_/A sky130_fd_sc_hd__o21ai_4
XFILLER_92_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _24277_/A vssd1 vssd1 vccd1 vccd1 _24335_/A sky130_fd_sc_hd__buf_8
XFILLER_229_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14735_ _15209_/S vssd1 vssd1 vccd1 vccd1 _16422_/S sky130_fd_sc_hd__buf_2
XFILLER_33_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17454_ _17454_/A vssd1 vssd1 vccd1 vccd1 _17455_/A sky130_fd_sc_hd__buf_2
XFILLER_33_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14666_ _16134_/S vssd1 vssd1 vccd1 vccd1 _16387_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13617_ _14515_/S vssd1 vssd1 vccd1 vccd1 _14495_/A sky130_fd_sc_hd__buf_2
X_16405_ _16405_/A _16405_/B vssd1 vssd1 vccd1 vccd1 _16405_/Y sky130_fd_sc_hd__nand2_1
X_17385_ _17384_/X _17389_/C _17366_/X vssd1 vssd1 vccd1 vccd1 _17385_/Y sky130_fd_sc_hd__a21oi_1
X_14597_ _14597_/A vssd1 vssd1 vccd1 vccd1 _14597_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19124_ _19579_/C _19121_/Y _19328_/S vssd1 vssd1 vccd1 vccd1 _19124_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13548_ _13466_/X _23542_/A _13547_/X _15127_/A vssd1 vssd1 vccd1 vccd1 _19912_/A
+ sky130_fd_sc_hd__o211ai_4
X_16336_ _16336_/A vssd1 vssd1 vccd1 vccd1 _16336_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_9_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19055_ _19055_/A vssd1 vssd1 vccd1 vccd1 _19055_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16267_ _26675_/Q _25715_/Q _16267_/S vssd1 vssd1 vccd1 vccd1 _16267_/X sky130_fd_sc_hd__mux2_1
X_13479_ _13479_/A vssd1 vssd1 vccd1 vccd1 _14757_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15218_ _25821_/Q _27255_/Q _15221_/S vssd1 vssd1 vccd1 vccd1 _15218_/X sky130_fd_sc_hd__mux2_1
X_18006_ _25571_/Q _18006_/B _18006_/C vssd1 vssd1 vccd1 vccd1 _18010_/D sky130_fd_sc_hd__nor3_1
XFILLER_173_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput304 _27330_/X vssd1 vssd1 vccd1 vccd1 clk1 sky130_fd_sc_hd__clkbuf_1
X_16198_ _14751_/A _16196_/X _16197_/X _15333_/A vssd1 vssd1 vccd1 vccd1 _16198_/X
+ sky130_fd_sc_hd__a211o_1
Xoutput315 _16760_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[19] sky130_fd_sc_hd__buf_2
XFILLER_236_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput326 _16709_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[3] sky130_fd_sc_hd__buf_2
Xoutput337 _16871_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[12] sky130_fd_sc_hd__buf_2
XFILLER_273_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ _16154_/B vssd1 vssd1 vccd1 vccd1 _16388_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_99_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput348 _16931_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[22] sky130_fd_sc_hd__buf_2
Xoutput359 _16822_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[3] sky130_fd_sc_hd__buf_2
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19957_ _19957_/A _19957_/B vssd1 vssd1 vccd1 vccd1 _19957_/Y sky130_fd_sc_hd__nand2_1
X_18908_ _19049_/A _19582_/C _18907_/Y _18037_/X vssd1 vssd1 vccd1 vccd1 _18908_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_228_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19888_ _19918_/A _19918_/B vssd1 vssd1 vccd1 vccd1 _19980_/B sky130_fd_sc_hd__xnor2_1
XFILLER_110_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18839_ _19076_/A vssd1 vssd1 vccd1 vccd1 _18839_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21850_ _21850_/A vssd1 vssd1 vccd1 vccd1 _26053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_270_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20801_ _20801_/A vssd1 vssd1 vccd1 vccd1 _25796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21781_ _20601_/X _26023_/Q _21787_/S vssd1 vssd1 vccd1 vccd1 _21782_/A sky130_fd_sc_hd__mux2_1
XFILLER_282_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23520_ _23520_/A vssd1 vssd1 vccd1 vccd1 _23520_/X sky130_fd_sc_hd__clkbuf_4
X_20732_ _20732_/A vssd1 vssd1 vccd1 vccd1 _25763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23451_ _23451_/A vssd1 vssd1 vccd1 vccd1 _26657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20663_ _26275_/Q _20660_/X _20662_/X _20658_/X vssd1 vssd1 vccd1 vccd1 _25738_/D
+ sky130_fd_sc_hd__o211a_1
X_22402_ _22638_/B vssd1 vssd1 vccd1 vccd1 _22402_/X sky130_fd_sc_hd__buf_8
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26170_ _26238_/CLK _26170_/D vssd1 vssd1 vccd1 vccd1 _26170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23382_ _26627_/Q _23060_/X _23386_/S vssd1 vssd1 vccd1 vccd1 _23383_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20594_ _20594_/A vssd1 vssd1 vccd1 vccd1 _25716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25121_ _20679_/A _25113_/X _25120_/X vssd1 vssd1 vccd1 vccd1 _25121_/Y sky130_fd_sc_hd__o21ai_1
X_22333_ _26224_/Q _22269_/A _22332_/X _22330_/X vssd1 vssd1 vccd1 vccd1 _26224_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25052_ _25106_/A vssd1 vssd1 vccd1 vccd1 _25052_/X sky130_fd_sc_hd__clkbuf_2
X_22264_ _22310_/A vssd1 vssd1 vccd1 vccd1 _22264_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24003_ _24003_/A vssd1 vssd1 vccd1 vccd1 _26875_/D sky130_fd_sc_hd__clkbuf_1
X_21215_ _21221_/A _21221_/B vssd1 vssd1 vccd1 vccd1 _21277_/A sky130_fd_sc_hd__or2_1
XFILLER_104_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22195_ _22195_/A vssd1 vssd1 vccd1 vccd1 _22195_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21146_ _21154_/A _21146_/B vssd1 vssd1 vccd1 vccd1 _21147_/A sky130_fd_sc_hd__or2_1
XFILLER_116_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25954_ _25992_/CLK _25954_/D vssd1 vssd1 vccd1 vccd1 _25954_/Q sky130_fd_sc_hd__dfxtp_1
X_21077_ _21113_/A vssd1 vssd1 vccd1 vccd1 _21077_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_246_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24905_ _24548_/A _24978_/B _24314_/X vssd1 vssd1 vccd1 vccd1 _24905_/Y sky130_fd_sc_hd__a21oi_1
X_20028_ _19894_/X _20027_/X _19902_/X vssd1 vssd1 vccd1 vccd1 _20028_/X sky130_fd_sc_hd__a21o_1
XFILLER_74_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25885_ _26604_/CLK _25885_/D vssd1 vssd1 vccd1 vccd1 _25885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12850_ _25599_/Q _12873_/A vssd1 vssd1 vccd1 vccd1 _12850_/Y sky130_fd_sc_hd__nor2_1
XFILLER_274_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24836_ _24833_/Y _24834_/X _24835_/X vssd1 vssd1 vccd1 vccd1 _27114_/D sky130_fd_sc_hd__a21oi_1
XFILLER_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _25024_/A vssd1 vssd1 vccd1 vccd1 _12781_/X sky130_fd_sc_hd__buf_8
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_24767_ _24770_/A _24767_/B vssd1 vssd1 vccd1 vccd1 _27098_/D sky130_fd_sc_hd__nor2_1
X_21979_ _26103_/Q _20894_/X _21983_/S vssd1 vssd1 vccd1 vccd1 _21980_/A sky130_fd_sc_hd__mux2_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _26652_/Q _25692_/Q _14520_/S vssd1 vssd1 vccd1 vccd1 _14520_/X sky130_fd_sc_hd__mux2_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23718_ _23718_/A vssd1 vssd1 vccd1 vccd1 _23718_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_215_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26506_ _27313_/CLK _26506_/D vssd1 vssd1 vccd1 vccd1 _26506_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24698_ _27082_/Q _24680_/X _24696_/Y _24697_/X vssd1 vssd1 vccd1 vccd1 _24699_/B
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _13344_/A _14448_/X _14450_/X _16022_/A vssd1 vssd1 vccd1 vccd1 _14451_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_230_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26437_ _26468_/CLK _26437_/D vssd1 vssd1 vccd1 vccd1 _26437_/Q sky130_fd_sc_hd__dfxtp_4
X_23649_ _23649_/A vssd1 vssd1 vccd1 vccd1 _26731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13402_/A vssd1 vssd1 vccd1 vccd1 _14713_/B sky130_fd_sc_hd__buf_4
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17170_ _20646_/A vssd1 vssd1 vccd1 vccd1 _17170_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26368_ _27275_/CLK _26368_/D vssd1 vssd1 vccd1 vccd1 _26368_/Q sky130_fd_sc_hd__dfxtp_4
X_14382_ _14064_/X _14380_/X _14381_/X _14067_/X vssd1 vssd1 vccd1 vccd1 _14387_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16121_ _20168_/A vssd1 vssd1 vccd1 vccd1 _16121_/Y sky130_fd_sc_hd__clkinv_2
X_13333_ _15932_/A vssd1 vssd1 vccd1 vccd1 _13335_/A sky130_fd_sc_hd__clkbuf_4
X_25319_ _23785_/X _27262_/Q _25319_/S vssd1 vssd1 vccd1 vccd1 _25320_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26299_ _26327_/CLK _26299_/D vssd1 vssd1 vccd1 vccd1 _26299_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_183_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16052_ _15265_/X _16049_/X _16051_/X _15538_/X vssd1 vssd1 vccd1 vccd1 _16052_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_170_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13264_ _13255_/X _26695_/Q _26823_/Q _16341_/S _15424_/A vssd1 vssd1 vccd1 vccd1
+ _13264_/X sky130_fd_sc_hd__a221o_1
XFILLER_6_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15003_ _27291_/Q _26484_/Q _15003_/S vssd1 vssd1 vccd1 vccd1 _15003_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13195_ _13309_/A _14076_/A vssd1 vssd1 vccd1 vccd1 _13773_/A sky130_fd_sc_hd__nor2_4
XFILLER_29_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19811_ _19796_/X _19809_/Y _20208_/A vssd1 vssd1 vccd1 vccd1 _19811_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_124_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19742_ _25664_/Q _25663_/Q _25662_/Q vssd1 vssd1 vccd1 vccd1 _19762_/B sky130_fd_sc_hd__and3_1
XFILLER_111_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16954_ _16954_/A vssd1 vssd1 vccd1 vccd1 _16954_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15905_ _14153_/X _26601_/Q _14009_/S _26341_/Q _14264_/S vssd1 vssd1 vccd1 vccd1
+ _15905_/X sky130_fd_sc_hd__o221a_1
X_19673_ _19673_/A _19673_/B vssd1 vssd1 vccd1 vccd1 _19675_/B sky130_fd_sc_hd__xnor2_2
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16885_ _16893_/A _16885_/B vssd1 vssd1 vccd1 vccd1 _16886_/A sky130_fd_sc_hd__and2_1
XFILLER_265_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18624_ _18608_/X _18622_/X _18623_/X vssd1 vssd1 vccd1 vccd1 _18626_/B sky130_fd_sc_hd__a21oi_1
X_15836_ _15836_/A _15836_/B vssd1 vssd1 vccd1 vccd1 _15836_/X sky130_fd_sc_hd__or2_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18555_ _18555_/A vssd1 vssd1 vccd1 vccd1 _18555_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15767_ _26795_/Q _26439_/Q _15930_/S vssd1 vssd1 vccd1 vccd1 _15767_/X sky130_fd_sc_hd__mux2_1
X_12979_ _25609_/Q _12981_/A _12952_/Y _12978_/X vssd1 vssd1 vccd1 vccd1 _23546_/A
+ sky130_fd_sc_hd__o22a_4
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17506_ _17992_/B _17772_/B vssd1 vssd1 vccd1 vccd1 _17679_/B sky130_fd_sc_hd__and2_1
XFILLER_206_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14718_ _14718_/A vssd1 vssd1 vccd1 vccd1 _14718_/X sky130_fd_sc_hd__clkbuf_2
X_18486_ _18489_/S _18258_/X _18485_/X vssd1 vssd1 vccd1 vccd1 _18896_/B sky130_fd_sc_hd__o21ai_2
XFILLER_61_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15698_ _18946_/A vssd1 vssd1 vccd1 vccd1 _15698_/Y sky130_fd_sc_hd__inv_4
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17437_ _25563_/Q _17437_/B vssd1 vssd1 vccd1 vccd1 _17438_/B sky130_fd_sc_hd__and2_1
XFILLER_33_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14649_ _14649_/A vssd1 vssd1 vccd1 vccd1 _14650_/A sky130_fd_sc_hd__buf_2
XFILLER_268_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17368_ _17365_/X _17370_/C _17367_/Y vssd1 vssd1 vccd1 vccd1 _25541_/D sky130_fd_sc_hd__o21a_1
XFILLER_193_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19107_ _18682_/X _18685_/X _19106_/Y _19018_/A vssd1 vssd1 vccd1 vccd1 _19107_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_118_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16319_ _26121_/Q _26022_/Q _16319_/S vssd1 vssd1 vccd1 vccd1 _16319_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17299_ _25520_/Q vssd1 vssd1 vccd1 vccd1 _17299_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_284_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19038_ _25741_/Q _19037_/C _25742_/Q vssd1 vssd1 vccd1 vccd1 _19039_/B sky130_fd_sc_hd__a21oi_1
XFILLER_133_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21000_ _25871_/Q _20878_/X _21004_/S vssd1 vssd1 vccd1 vccd1 _21001_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22951_ _22951_/A vssd1 vssd1 vccd1 vccd1 _26450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_284_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21902_ _21959_/S vssd1 vssd1 vccd1 vccd1 _21911_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25670_ _25670_/CLK _25670_/D vssd1 vssd1 vccd1 vccd1 _25670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22882_ _26420_/Q _22733_/X _22884_/S vssd1 vssd1 vccd1 vccd1 _22883_/A sky130_fd_sc_hd__mux2_1
XFILLER_271_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24621_ _24621_/A _24621_/B vssd1 vssd1 vccd1 vccd1 _24621_/Y sky130_fd_sc_hd__nand2_1
XFILLER_243_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21833_ _21833_/A vssd1 vssd1 vccd1 vccd1 _26045_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_37_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26827_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24552_ _27038_/Q _24546_/X _24550_/Y _24551_/X vssd1 vssd1 vccd1 vccd1 _27038_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21764_ _21764_/A vssd1 vssd1 vccd1 vccd1 _26015_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23503_ _23503_/A vssd1 vssd1 vccd1 vccd1 _26681_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27271_ _27272_/CLK _27271_/D vssd1 vssd1 vccd1 vccd1 _27271_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20715_ _21887_/B vssd1 vssd1 vccd1 vccd1 _25249_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_197_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24483_ _24492_/A _24960_/A vssd1 vssd1 vccd1 vccd1 _24483_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21695_ _21695_/A vssd1 vssd1 vccd1 vccd1 _25986_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26222_ _26222_/CLK _26222_/D vssd1 vssd1 vccd1 vccd1 _26222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23434_ _26651_/Q _23136_/X _23434_/S vssd1 vssd1 vccd1 vccd1 _23435_/A sky130_fd_sc_hd__mux2_1
X_20646_ _20646_/A vssd1 vssd1 vccd1 vccd1 _20646_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26153_ _27252_/CLK _26153_/D vssd1 vssd1 vccd1 vccd1 _26153_/Q sky130_fd_sc_hd__dfxtp_1
X_23365_ _23421_/A vssd1 vssd1 vccd1 vccd1 _23434_/S sky130_fd_sc_hd__buf_6
XFILLER_192_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20577_ _20575_/X _25712_/Q _20593_/S vssd1 vssd1 vccd1 vccd1 _20578_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25104_ _24719_/Y _25097_/X _25103_/Y _25082_/X vssd1 vssd1 vccd1 vccd1 _25104_/X
+ sky130_fd_sc_hd__a31o_1
X_22316_ _22630_/B vssd1 vssd1 vccd1 vccd1 _22316_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26084_ _27315_/CLK _26084_/D vssd1 vssd1 vccd1 vccd1 _26084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23296_ _20496_/X _26589_/Q _23302_/S vssd1 vssd1 vccd1 vccd1 _23297_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25035_ _20637_/A _25031_/X _25034_/X vssd1 vssd1 vccd1 vccd1 _25035_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_279_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22247_ _26194_/Q _22222_/X _22238_/X _26295_/Q _22241_/X vssd1 vssd1 vccd1 vccd1
+ _22247_/X sky130_fd_sc_hd__a221o_1
XFILLER_106_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22178_ _26177_/Q _22169_/X _22177_/X _22164_/X vssd1 vssd1 vccd1 vccd1 _26177_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21129_ _21129_/A vssd1 vssd1 vccd1 vccd1 _25916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26986_ _26987_/CLK _26986_/D vssd1 vssd1 vccd1 vccd1 _26986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13951_ _26526_/Q _26134_/Q _13951_/S vssd1 vssd1 vccd1 vccd1 _13951_/X sky130_fd_sc_hd__mux2_1
X_25937_ _27154_/CLK _25937_/D vssd1 vssd1 vccd1 vccd1 _25937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12902_ _12902_/A vssd1 vssd1 vccd1 vccd1 _12902_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13882_ _14269_/S vssd1 vssd1 vccd1 vccd1 _15890_/S sky130_fd_sc_hd__clkbuf_4
X_16670_ _21235_/A _21198_/A vssd1 vssd1 vccd1 vccd1 _21603_/A sky130_fd_sc_hd__or2_4
X_25868_ _27293_/CLK _25868_/D vssd1 vssd1 vccd1 vccd1 _25868_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_235_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15621_ _25614_/Q _14596_/A _15620_/X _14617_/A vssd1 vssd1 vccd1 vccd1 _23562_/A
+ sky130_fd_sc_hd__o22a_4
X_12833_ _13916_/A vssd1 vssd1 vccd1 vccd1 _14025_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24819_ _20648_/A _24810_/X _24682_/Y _24811_/X vssd1 vssd1 vccd1 vccd1 _24819_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_27_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25799_ _26520_/CLK _25799_/D vssd1 vssd1 vccd1 vccd1 _25799_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _18340_/A vssd1 vssd1 vccd1 vccd1 _19256_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _25585_/Q vssd1 vssd1 vccd1 vccd1 _13582_/A sky130_fd_sc_hd__inv_2
X_15552_ _15538_/X _15546_/X _15551_/X _14677_/A vssd1 vssd1 vccd1 vccd1 _15552_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _13890_/X _26588_/Q _15989_/S _26328_/Q _13862_/A vssd1 vssd1 vccd1 vccd1
+ _14503_/X sky130_fd_sc_hd__o221a_1
XFILLER_188_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18271_ _18598_/S _18271_/B vssd1 vssd1 vccd1 vccd1 _18271_/X sky130_fd_sc_hd__or2_2
X_15483_ _15441_/X _15526_/S _15244_/A _15482_/Y vssd1 vssd1 vccd1 vccd1 _17840_/A
+ sky130_fd_sc_hd__o22a_4
X_12695_ _25588_/Q vssd1 vssd1 vccd1 vccd1 _13105_/B sky130_fd_sc_hd__buf_8
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17222_ _17222_/A _17222_/B vssd1 vssd1 vccd1 vccd1 _17223_/A sky130_fd_sc_hd__and2_1
X_14434_ _14153_/A _25830_/Q _26030_/Q _14520_/S _14352_/S vssd1 vssd1 vccd1 vccd1
+ _14434_/X sky130_fd_sc_hd__a221o_1
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 core_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14365_ _27265_/Q _26458_/Q _14365_/S vssd1 vssd1 vccd1 vccd1 _14365_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17153_ _17200_/A _17153_/B vssd1 vssd1 vccd1 vccd1 _17154_/A sky130_fd_sc_hd__and2_1
Xinput25 core_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_1
Xinput36 core_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 dout0[13] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13316_ _26791_/Q _26435_/Q _16277_/S vssd1 vssd1 vccd1 vccd1 _13316_/X sky130_fd_sc_hd__mux2_1
X_16104_ _16104_/A _16104_/B vssd1 vssd1 vccd1 vccd1 _16104_/X sky130_fd_sc_hd__or2_1
Xinput58 dout0[23] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_2
X_17084_ _26234_/Q vssd1 vssd1 vccd1 vccd1 _17085_/A sky130_fd_sc_hd__buf_2
XFILLER_6_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput69 dout0[33] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_1
X_14296_ _26523_/Q _26131_/Q _14296_/S vssd1 vssd1 vccd1 vccd1 _14296_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13247_ _15300_/A vssd1 vssd1 vccd1 vccd1 _16261_/S sky130_fd_sc_hd__buf_6
X_16035_ _17828_/A _16035_/B vssd1 vssd1 vccd1 vccd1 _18735_/S sky130_fd_sc_hd__nand2_1
XFILLER_115_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13178_ _17971_/B _18006_/C vssd1 vssd1 vccd1 vccd1 _13179_/A sky130_fd_sc_hd__nor2_2
XFILLER_69_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17986_ _17986_/A _18271_/B vssd1 vssd1 vccd1 vccd1 _18364_/A sky130_fd_sc_hd__or2_1
XFILLER_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19725_ _19766_/A vssd1 vssd1 vccd1 vccd1 _19725_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_266_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16937_ _15192_/B _16952_/A _16812_/A vssd1 vssd1 vccd1 vccd1 _16942_/A sky130_fd_sc_hd__o21a_1
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19656_ _24706_/A vssd1 vssd1 vccd1 vccd1 _19905_/A sky130_fd_sc_hd__clkbuf_2
X_16868_ _16868_/A _16868_/B vssd1 vssd1 vccd1 vccd1 _16868_/X sky130_fd_sc_hd__or2_1
XFILLER_265_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18607_ _18596_/Y _18606_/X _18003_/A vssd1 vssd1 vccd1 vccd1 _18607_/X sky130_fd_sc_hd__a21o_1
X_15819_ _15815_/X _15818_/X _15819_/S vssd1 vssd1 vccd1 vccd1 _15819_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19587_ _19583_/Y _19586_/X _17512_/X vssd1 vssd1 vccd1 vccd1 _19670_/A sky130_fd_sc_hd__a21oi_4
XFILLER_281_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16799_ _19639_/A vssd1 vssd1 vccd1 vccd1 _16838_/A sky130_fd_sc_hd__buf_4
XFILLER_280_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18538_ _18942_/B vssd1 vssd1 vccd1 vccd1 _19235_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18469_ _18469_/A vssd1 vssd1 vccd1 vccd1 _18469_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_221_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20500_ _23693_/A vssd1 vssd1 vccd1 vccd1 _20500_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21480_ _21544_/A vssd1 vssd1 vccd1 vccd1 _21480_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20431_ _27162_/Q vssd1 vssd1 vccd1 vccd1 _20434_/A sky130_fd_sc_hd__buf_2
XFILLER_193_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_155_wb_clk_i clkbuf_opt_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27188_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_147_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23150_ _26524_/Q _23050_/X _23150_/S vssd1 vssd1 vccd1 vccd1 _23151_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20362_ _20362_/A _20362_/B vssd1 vssd1 vccd1 vccd1 _20362_/X sky130_fd_sc_hd__and2_1
XFILLER_174_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22101_ _26158_/Q _20967_/X _22103_/S vssd1 vssd1 vccd1 vccd1 _22102_/A sky130_fd_sc_hd__mux2_1
X_23081_ _23081_/A vssd1 vssd1 vccd1 vccd1 _26501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20293_ _20268_/X _20271_/Y _20291_/Y _20292_/X vssd1 vssd1 vccd1 vccd1 _20293_/Y
+ sky130_fd_sc_hd__o211ai_2
X_22032_ _22032_/A vssd1 vssd1 vccd1 vccd1 _26127_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26840_ _26904_/CLK _26840_/D vssd1 vssd1 vccd1 vccd1 _26840_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26771_ _26931_/CLK _26771_/D vssd1 vssd1 vccd1 vccd1 _26771_/Q sky130_fd_sc_hd__dfxtp_1
X_23983_ _26866_/Q _23581_/X _23987_/S vssd1 vssd1 vccd1 vccd1 _23984_/A sky130_fd_sc_hd__mux2_1
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22934_ _26443_/Q _22704_/X _22934_/S vssd1 vssd1 vccd1 vccd1 _22935_/A sky130_fd_sc_hd__mux2_1
X_25722_ _27293_/CLK _25722_/D vssd1 vssd1 vccd1 vccd1 _25722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25653_ _25660_/CLK _25653_/D vssd1 vssd1 vccd1 vccd1 _25653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22865_ _26412_/Q _22707_/X _22873_/S vssd1 vssd1 vccd1 vccd1 _22866_/A sky130_fd_sc_hd__mux2_1
XFILLER_272_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21816_ _26038_/Q _20900_/X _21816_/S vssd1 vssd1 vccd1 vccd1 _21817_/A sky130_fd_sc_hd__mux2_1
X_24604_ _27057_/Q _24602_/X _24603_/Y _24593_/X vssd1 vssd1 vccd1 vccd1 _27057_/D
+ sky130_fd_sc_hd__o211a_1
X_25584_ _26684_/CLK _25584_/D vssd1 vssd1 vccd1 vccd1 _25584_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_19_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22796_ _26382_/Q _22714_/X _22800_/S vssd1 vssd1 vccd1 vccd1 _22797_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24535_ _26324_/Q _24473_/X _24474_/X input239/X _21885_/A vssd1 vssd1 vccd1 vccd1
+ _24535_/X sky130_fd_sc_hd__a221o_1
X_27323_ _27324_/CLK _27323_/D vssd1 vssd1 vccd1 vccd1 _27323_/Q sky130_fd_sc_hd__dfxtp_1
X_21747_ _21747_/A vssd1 vssd1 vccd1 vccd1 _26007_/D sky130_fd_sc_hd__clkbuf_1
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24466_ _24494_/A vssd1 vssd1 vccd1 vccd1 _24492_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27254_ _27319_/CLK _27254_/D vssd1 vssd1 vccd1 vccd1 _27254_/Q sky130_fd_sc_hd__dfxtp_1
X_21678_ _21678_/A vssd1 vssd1 vccd1 vccd1 _25978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26205_ _26257_/CLK _26205_/D vssd1 vssd1 vccd1 vccd1 _26205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23417_ _26643_/Q _23111_/X _23419_/S vssd1 vssd1 vccd1 vccd1 _23418_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20629_ _26263_/Q _17190_/X _20628_/X _19965_/X vssd1 vssd1 vccd1 vccd1 _25726_/D
+ sky130_fd_sc_hd__o211a_1
X_27185_ _27188_/CLK _27185_/D vssd1 vssd1 vccd1 vccd1 _27185_/Q sky130_fd_sc_hd__dfxtp_1
X_24397_ _24392_/X _25603_/Q _24396_/X vssd1 vssd1 vccd1 vccd1 _24920_/A sky130_fd_sc_hd__o21ai_4
XFILLER_149_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26136_ _26601_/CLK _26136_/D vssd1 vssd1 vccd1 vccd1 _26136_/Q sky130_fd_sc_hd__dfxtp_4
X_14150_ _14148_/X _14149_/X _14272_/S vssd1 vssd1 vccd1 vccd1 _14150_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23348_ _23348_/A vssd1 vssd1 vccd1 vccd1 _23357_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_192_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13101_ _15806_/S vssd1 vssd1 vccd1 vccd1 _13402_/A sky130_fd_sc_hd__clkbuf_4
X_26067_ _26593_/CLK _26067_/D vssd1 vssd1 vccd1 vccd1 _26067_/Q sky130_fd_sc_hd__dfxtp_1
X_14081_ _14560_/S _19769_/A _14080_/X vssd1 vssd1 vccd1 vccd1 _17801_/B sky130_fd_sc_hd__a21boi_4
XFILLER_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23279_ _26582_/Q _23133_/X _23281_/S vssd1 vssd1 vccd1 vccd1 _23280_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13032_ _13993_/A vssd1 vssd1 vccd1 vccd1 _14176_/S sky130_fd_sc_hd__buf_2
X_25018_ _24649_/Y _25014_/X _25017_/Y _24773_/X vssd1 vssd1 vccd1 vccd1 _25018_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_279_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17840_ _17840_/A _15528_/B vssd1 vssd1 vccd1 vccd1 _17840_/X sky130_fd_sc_hd__or2b_1
XFILLER_120_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17771_ _18383_/A vssd1 vssd1 vccd1 vccd1 _18474_/A sky130_fd_sc_hd__clkbuf_2
X_26969_ _27001_/CLK _26969_/D vssd1 vssd1 vccd1 vccd1 _26969_/Q sky130_fd_sc_hd__dfxtp_1
X_14983_ _14733_/A _14981_/X _14982_/X _14760_/A vssd1 vssd1 vccd1 vccd1 _14987_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19510_ _25639_/Q _19510_/B vssd1 vssd1 vccd1 vccd1 _19510_/X sky130_fd_sc_hd__or2_1
X_16722_ _25667_/Q vssd1 vssd1 vccd1 vccd1 _22485_/A sky130_fd_sc_hd__buf_4
XFILLER_47_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13934_ _25636_/Q _15443_/B _13578_/A _25604_/Q vssd1 vssd1 vccd1 vccd1 _13934_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_219_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19441_ _18742_/X _19431_/X _19440_/X vssd1 vssd1 vccd1 vccd1 _19441_/X sky130_fd_sc_hd__a21o_4
XFILLER_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16653_ _25683_/Q _25682_/Q _25681_/Q _25680_/Q vssd1 vssd1 vccd1 vccd1 _16654_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_62_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13865_ _14263_/S vssd1 vssd1 vccd1 vccd1 _14245_/S sky130_fd_sc_hd__buf_2
XFILLER_74_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_504 _25925_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_515 _17067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15604_ _15924_/A _15604_/B vssd1 vssd1 vccd1 vccd1 _15604_/X sky130_fd_sc_hd__or2_1
XINSDIODE2_526 _17040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19372_ _17327_/X _18444_/A _19369_/X _19371_/X _18469_/A vssd1 vssd1 vccd1 vccd1
+ _19372_/X sky130_fd_sc_hd__o221a_1
X_12816_ _25500_/Q vssd1 vssd1 vccd1 vccd1 _12822_/A sky130_fd_sc_hd__dlymetal6s2s_1
XINSDIODE2_537 _17011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16584_ _19571_/B vssd1 vssd1 vccd1 vccd1 _16853_/A sky130_fd_sc_hd__buf_2
XINSDIODE2_548 _14559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13796_ _13274_/X _13778_/X _13787_/X _13795_/X _14722_/A vssd1 vssd1 vccd1 vccd1
+ _13796_/X sky130_fd_sc_hd__a221o_2
XFILLER_215_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18323_ _18904_/A vssd1 vssd1 vccd1 vccd1 _18942_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_203_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15535_ _27312_/Q _26569_/Q _16305_/A vssd1 vssd1 vccd1 vccd1 _15535_/X sky130_fd_sc_hd__mux2_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _16071_/S vssd1 vssd1 vccd1 vccd1 _15376_/S sky130_fd_sc_hd__buf_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18254_ _18254_/A vssd1 vssd1 vccd1 vccd1 _18262_/S sky130_fd_sc_hd__clkbuf_4
X_15466_ _16059_/S _15463_/X _15465_/X _15538_/A vssd1 vssd1 vccd1 vccd1 _15466_/X
+ sky130_fd_sc_hd__a211o_1
X_12678_ _25571_/Q vssd1 vssd1 vccd1 vccd1 _17504_/A sky130_fd_sc_hd__clkinv_2
XFILLER_230_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17205_ _17205_/A vssd1 vssd1 vccd1 vccd1 _25494_/D sky130_fd_sc_hd__clkbuf_1
X_14417_ _26065_/Q _14713_/D _14416_/X _15990_/S vssd1 vssd1 vccd1 vccd1 _14421_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_156_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18185_ _18251_/C _18185_/B vssd1 vssd1 vccd1 vccd1 _19571_/C sky130_fd_sc_hd__and2_1
X_15397_ _15321_/X _26896_/Q _26768_/Q _15209_/S _14791_/A vssd1 vssd1 vccd1 vccd1
+ _15397_/X sky130_fd_sc_hd__a221o_1
XFILLER_184_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17136_ _25475_/Q _17105_/X _17107_/X _25572_/Q vssd1 vssd1 vccd1 vccd1 _17137_/B
+ sky130_fd_sc_hd__a22o_1
X_14348_ _25831_/Q _26031_/Q _14348_/S vssd1 vssd1 vccd1 vccd1 _14348_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14279_ _14523_/A _14251_/X _14261_/X _14278_/X vssd1 vssd1 vccd1 vccd1 _14279_/X
+ sky130_fd_sc_hd__o31a_2
X_17067_ _25975_/Q _17061_/X _16995_/X _17063_/X vssd1 vssd1 vccd1 vccd1 _17067_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_144_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16018_ _13813_/X _26108_/Q _26009_/Q _13534_/S _13814_/X vssd1 vssd1 vccd1 vccd1
+ _16018_/X sky130_fd_sc_hd__a221o_1
XFILLER_171_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ _25571_/Q _17971_/A _18006_/B vssd1 vssd1 vccd1 vccd1 _17978_/C sky130_fd_sc_hd__or3_1
XFILLER_214_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19708_ _19708_/A vssd1 vssd1 vccd1 vccd1 _20091_/A sky130_fd_sc_hd__buf_2
XFILLER_84_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20980_ _26584_/Q _20986_/B _25867_/D vssd1 vssd1 vccd1 vccd1 _20981_/A sky130_fd_sc_hd__and3_1
XFILLER_226_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19639_ _19639_/A _19639_/B _25119_/A vssd1 vssd1 vccd1 vccd1 _25114_/A sky130_fd_sc_hd__nor3_4
XFILLER_53_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22650_ _23693_/A vssd1 vssd1 vccd1 vccd1 _22650_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_207_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21601_ _21599_/X _21600_/X _21589_/X vssd1 vssd1 vccd1 vccd1 _21601_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22581_ _22607_/A vssd1 vssd1 vccd1 vccd1 _22591_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_240_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24320_ _26998_/Q _24320_/B vssd1 vssd1 vccd1 vccd1 _24326_/C sky130_fd_sc_hd__and2_1
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21532_ _25957_/Q _21506_/X _21530_/Y _21531_/X vssd1 vssd1 vccd1 vccd1 _25957_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_221_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24251_ _24285_/A _24251_/B _24252_/B vssd1 vssd1 vccd1 vccd1 _26973_/D sky130_fd_sc_hd__nor3_1
X_21463_ input50/X input85/X _21489_/S vssd1 vssd1 vccd1 vccd1 _21464_/A sky130_fd_sc_hd__mux2_8
XFILLER_239_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23202_ _23202_/A vssd1 vssd1 vccd1 vccd1 _26547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20414_ _20389_/A _20391_/B _20389_/B vssd1 vssd1 vccd1 vccd1 _20415_/B sky130_fd_sc_hd__a21boi_2
X_24182_ _26951_/Q _24184_/C _17137_/A vssd1 vssd1 vccd1 vccd1 _24183_/B sky130_fd_sc_hd__o21ai_1
XFILLER_119_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21394_ _21342_/X _21393_/X _21336_/X vssd1 vssd1 vccd1 vccd1 _21394_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_146_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23133_ _23606_/A vssd1 vssd1 vccd1 vccd1 _23133_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20345_ _20179_/X _20344_/X _20186_/X vssd1 vssd1 vccd1 vccd1 _20345_/X sky130_fd_sc_hd__a21o_1
XFILLER_49_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23064_ _26496_/Q _23063_/X _23067_/S vssd1 vssd1 vccd1 vccd1 _23065_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20276_ _20276_/A vssd1 vssd1 vccd1 vccd1 _20276_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22015_ _22015_/A vssd1 vssd1 vccd1 vccd1 _26119_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput204 localMemory_wb_adr_i[22] vssd1 vssd1 vccd1 vccd1 _17456_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_216_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput215 localMemory_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input215/X sky130_fd_sc_hd__buf_6
XFILLER_76_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput226 localMemory_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input226/X sky130_fd_sc_hd__clkbuf_8
XTAP_5448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26823_ _26823_/CLK _26823_/D vssd1 vssd1 vccd1 vccd1 _26823_/Q sky130_fd_sc_hd__dfxtp_2
Xinput237 localMemory_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input237/X sky130_fd_sc_hd__buf_4
XTAP_5459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26856_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput248 localMemory_wb_sel_i[1] vssd1 vssd1 vccd1 vccd1 input248/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput259 manufacturerID[5] vssd1 vssd1 vccd1 vccd1 input259/X sky130_fd_sc_hd__clkbuf_2
XFILLER_276_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26754_ _27301_/CLK _26754_/D vssd1 vssd1 vccd1 vccd1 _26754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23966_ _23966_/A vssd1 vssd1 vccd1 vccd1 _26858_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25705_ _27276_/CLK _25705_/D vssd1 vssd1 vccd1 vccd1 _25705_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_216_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22917_ _26435_/Q _22679_/X _22923_/S vssd1 vssd1 vccd1 vccd1 _22918_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26685_ _26877_/CLK _26685_/D vssd1 vssd1 vccd1 vccd1 _26685_/Q sky130_fd_sc_hd__dfxtp_1
X_23897_ _23897_/A vssd1 vssd1 vccd1 vccd1 _26827_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22848_ _22848_/A vssd1 vssd1 vccd1 vccd1 _26404_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25636_ _26297_/CLK _25636_/D vssd1 vssd1 vccd1 vccd1 _25636_/Q sky130_fd_sc_hd__dfxtp_1
X_13650_ _13832_/A _13647_/X _13649_/X _15769_/A vssd1 vssd1 vccd1 vccd1 _13650_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_32_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13581_ _26497_/Q _26369_/Q _13589_/S vssd1 vssd1 vccd1 vccd1 _13581_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22779_ _22779_/A vssd1 vssd1 vccd1 vccd1 _26374_/D sky130_fd_sc_hd__clkbuf_1
X_25567_ _25596_/CLK _25567_/D vssd1 vssd1 vccd1 vccd1 _25567_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27306_ _27306_/CLK _27306_/D vssd1 vssd1 vccd1 vccd1 _27306_/Q sky130_fd_sc_hd__dfxtp_1
X_15320_ _27317_/Q _26574_/Q _16433_/S vssd1 vssd1 vccd1 vccd1 _15320_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24518_ _24518_/A _24621_/A vssd1 vssd1 vccd1 vccd1 _24518_/Y sky130_fd_sc_hd__nand2_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25498_ _26683_/CLK _25498_/D vssd1 vssd1 vccd1 vccd1 _25498_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27237_ _27238_/CLK _27237_/D vssd1 vssd1 vccd1 vccd1 _27237_/Q sky130_fd_sc_hd__dfxtp_1
X_15251_ _27317_/Q _26574_/Q _16377_/S vssd1 vssd1 vccd1 vccd1 _15251_/X sky130_fd_sc_hd__mux2_1
X_24449_ _26308_/Q _21881_/X _21883_/X input221/X _24404_/X vssd1 vssd1 vccd1 vccd1
+ _24449_/X sky130_fd_sc_hd__a221o_1
XFILLER_32_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14202_ _15588_/A _26688_/Q _26816_/Q _13675_/S _12738_/C vssd1 vssd1 vccd1 vccd1
+ _14202_/X sky130_fd_sc_hd__a221o_1
X_15182_ _15180_/X _15181_/X _16397_/S vssd1 vssd1 vccd1 vccd1 _15182_/X sky130_fd_sc_hd__mux2_1
X_27168_ _27173_/CLK _27168_/D vssd1 vssd1 vccd1 vccd1 _27168_/Q sky130_fd_sc_hd__dfxtp_1
X_14133_ _14133_/A _14133_/B vssd1 vssd1 vccd1 vccd1 _14133_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26119_ _27329_/A _26119_/D vssd1 vssd1 vccd1 vccd1 _26119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19990_ _24749_/A vssd1 vssd1 vccd1 vccd1 _24768_/A sky130_fd_sc_hd__buf_4
X_27099_ _27198_/CLK _27099_/D vssd1 vssd1 vccd1 vccd1 _27099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14064_ _14468_/A vssd1 vssd1 vccd1 vccd1 _14064_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_140_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18941_ _18941_/A _18941_/B vssd1 vssd1 vccd1 vccd1 _18941_/Y sky130_fd_sc_hd__xnor2_2
X_13015_ _13015_/A vssd1 vssd1 vccd1 vccd1 _14355_/A sky130_fd_sc_hd__buf_2
XFILLER_239_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18872_ _27051_/Q _18747_/X _18869_/X _18871_/X _18761_/X vssd1 vssd1 vccd1 vccd1
+ _18872_/X sky130_fd_sc_hd__o221a_2
XFILLER_39_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17823_ _13554_/A _17820_/Y _17822_/Y vssd1 vssd1 vccd1 vccd1 _17823_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_39_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__buf_2
XFILLER_48_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17754_ _18391_/A vssd1 vssd1 vccd1 vccd1 _18815_/A sky130_fd_sc_hd__buf_2
XFILLER_48_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14966_ _14693_/S _14963_/X _14965_/X _14662_/A vssd1 vssd1 vccd1 vccd1 _14966_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_270_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16705_ _16770_/A vssd1 vssd1 vccd1 vccd1 _16705_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13917_ _14323_/B vssd1 vssd1 vccd1 vccd1 _14485_/B sky130_fd_sc_hd__clkbuf_2
X_17685_ _17685_/A vssd1 vssd1 vccd1 vccd1 _21283_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_263_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14897_ _16359_/S vssd1 vssd1 vccd1 vccd1 _16354_/S sky130_fd_sc_hd__buf_2
XINSDIODE2_301 _26464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_312 _19620_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19424_ _16557_/A _19389_/C _17849_/Y vssd1 vssd1 vccd1 vccd1 _19424_/X sky130_fd_sc_hd__o21a_1
XFILLER_223_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_323 _19616_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16636_ _16751_/A _16748_/A _16636_/C _16636_/D vssd1 vssd1 vccd1 vccd1 _16637_/D
+ sky130_fd_sc_hd__or4_1
X_13848_ _13346_/A _13846_/X _13847_/X _14228_/A vssd1 vssd1 vccd1 vccd1 _13848_/X
+ sky130_fd_sc_hd__a31o_1
XINSDIODE2_334 _19609_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_345 _19617_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_356 _19612_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_367 _20487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19355_ _19355_/A _19355_/B _19355_/C vssd1 vssd1 vccd1 vccd1 _19356_/B sky130_fd_sc_hd__and3_1
XFILLER_62_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16567_ _19325_/A _16567_/B vssd1 vssd1 vccd1 vccd1 _19318_/B sky130_fd_sc_hd__xnor2_4
XINSDIODE2_378 _16998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13779_ _13779_/A vssd1 vssd1 vccd1 vccd1 _14727_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_389 _17027_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18306_ _18805_/A _18306_/B _18306_/C vssd1 vssd1 vccd1 vccd1 _18306_/X sky130_fd_sc_hd__or3_2
X_15518_ _15488_/A _26926_/Q _26410_/Q _15596_/S _15760_/A vssd1 vssd1 vccd1 vccd1
+ _15518_/X sky130_fd_sc_hd__a221o_1
XFILLER_149_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19286_ _19042_/A _19256_/B _19218_/X _19774_/A _19253_/X vssd1 vssd1 vccd1 vccd1
+ _19286_/X sky130_fd_sc_hd__a221o_2
XFILLER_203_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16498_ _26519_/Q _26391_/Q _16498_/S vssd1 vssd1 vccd1 vccd1 _16498_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18237_ _27104_/Q _19056_/A _18235_/X _18236_/X vssd1 vssd1 vccd1 vccd1 _18237_/X
+ sky130_fd_sc_hd__o22a_2
X_15449_ _26638_/Q _26734_/Q _15471_/S vssd1 vssd1 vccd1 vccd1 _15449_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18168_ _18458_/A vssd1 vssd1 vccd1 vccd1 _18825_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_175_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17119_ _24630_/A vssd1 vssd1 vccd1 vccd1 _22377_/A sky130_fd_sc_hd__buf_4
X_18099_ _18440_/A vssd1 vssd1 vccd1 vccd1 _18557_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_209_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20130_ _27118_/Q _20079_/X _20112_/X _20129_/X vssd1 vssd1 vccd1 vccd1 _20130_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20061_ _20061_/A _20061_/B vssd1 vssd1 vccd1 vccd1 _20061_/X sky130_fd_sc_hd__and2_1
XFILLER_258_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_16 _18888_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_27 _19172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_38 _19441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23820_ _23820_/A vssd1 vssd1 vccd1 vccd1 _26793_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_49 _20628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23751_ _23767_/A vssd1 vssd1 vccd1 vccd1 _23764_/S sky130_fd_sc_hd__buf_4
X_20963_ _20963_/A vssd1 vssd1 vccd1 vccd1 _25857_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22702_ _26346_/Q _22701_/X _22705_/S vssd1 vssd1 vccd1 vccd1 _22703_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26470_ _27277_/CLK _26470_/D vssd1 vssd1 vccd1 vccd1 _26470_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_246_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23682_ _26747_/Q _23609_/X _23682_/S vssd1 vssd1 vccd1 vccd1 _23683_/A sky130_fd_sc_hd__mux2_1
X_20894_ _23709_/A vssd1 vssd1 vccd1 vccd1 _20894_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22633_ _22633_/A _22638_/C vssd1 vssd1 vccd1 vccd1 _22633_/X sky130_fd_sc_hd__or2_1
XFILLER_242_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25421_ _25421_/A vssd1 vssd1 vccd1 vccd1 _27306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_170_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25670_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_41_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25352_ _27276_/Q _23728_/A _25354_/S vssd1 vssd1 vccd1 vccd1 _25353_/A sky130_fd_sc_hd__mux2_1
X_22564_ _22553_/X _22563_/Y _22561_/X vssd1 vssd1 vccd1 vccd1 _26301_/D sky130_fd_sc_hd__a21oi_1
XFILLER_210_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24303_ _26992_/Q _24303_/B vssd1 vssd1 vccd1 vccd1 _24309_/C sky130_fd_sc_hd__and2_1
X_21515_ _21480_/X _21514_/X _21473_/X vssd1 vssd1 vccd1 vccd1 _21515_/Y sky130_fd_sc_hd__o21ai_1
X_25283_ _25283_/A vssd1 vssd1 vccd1 vccd1 _27245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22495_ _22495_/A vssd1 vssd1 vccd1 vccd1 _26272_/D sky130_fd_sc_hd__clkbuf_1
X_24234_ _24237_/A _24240_/C vssd1 vssd1 vccd1 vccd1 _24234_/Y sky130_fd_sc_hd__nor2_1
X_27022_ _27022_/CLK _27022_/D vssd1 vssd1 vccd1 vccd1 _27022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21446_ _21444_/X _21445_/X _21433_/X vssd1 vssd1 vccd1 vccd1 _21446_/X sky130_fd_sc_hd__a21o_1
XFILLER_163_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24165_ _26945_/Q _24163_/B _24164_/Y vssd1 vssd1 vccd1 vccd1 _26945_/D sky130_fd_sc_hd__o21a_1
X_21377_ _25945_/Q _21310_/X _21376_/Y _21330_/X vssd1 vssd1 vccd1 vccd1 _25945_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_107_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23116_ _23116_/A vssd1 vssd1 vccd1 vccd1 _26512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20328_ _20376_/A vssd1 vssd1 vccd1 vccd1 _20328_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_24096_ _26916_/Q _23536_/X _24098_/S vssd1 vssd1 vccd1 vccd1 _24097_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23047_ _23520_/A vssd1 vssd1 vccd1 vccd1 _23047_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20259_ _20379_/A _20259_/B vssd1 vssd1 vccd1 vccd1 _20305_/B sky130_fd_sc_hd__and2_1
XFILLER_62_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26806_ _27322_/CLK _26806_/D vssd1 vssd1 vccd1 vccd1 _26806_/Q sky130_fd_sc_hd__dfxtp_1
X_14820_ _14820_/A vssd1 vssd1 vccd1 vccd1 _16185_/A sky130_fd_sc_hd__clkbuf_4
XTAP_5289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24998_ _25124_/A vssd1 vssd1 vccd1 vccd1 _25142_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _14751_/A vssd1 vssd1 vccd1 vccd1 _15085_/A sky130_fd_sc_hd__buf_2
X_26737_ _27252_/CLK _26737_/D vssd1 vssd1 vccd1 vccd1 _26737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_251_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23949_ _23949_/A vssd1 vssd1 vccd1 vccd1 _26850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _15141_/A _13700_/X _13701_/X _12702_/A vssd1 vssd1 vccd1 vccd1 _13702_/X
+ sky130_fd_sc_hd__o211a_1
X_17470_ _17470_/A _17706_/B vssd1 vssd1 vccd1 vccd1 _17470_/Y sky130_fd_sc_hd__nor2_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _14682_/A vssd1 vssd1 vccd1 vccd1 _14683_/A sky130_fd_sc_hd__buf_2
XFILLER_72_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26668_ _26671_/CLK _26668_/D vssd1 vssd1 vccd1 vccd1 _26668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16421_ _15095_/S _16418_/X _16420_/X _14802_/A vssd1 vssd1 vccd1 vccd1 _16421_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_72_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13633_ _13717_/A _13607_/X _13632_/X _13174_/A vssd1 vssd1 vccd1 vccd1 _13633_/X
+ sky130_fd_sc_hd__a211o_4
X_25619_ _27327_/CLK _25619_/D vssd1 vssd1 vccd1 vccd1 _25619_/Q sky130_fd_sc_hd__dfxtp_2
X_26599_ _26599_/CLK _26599_/D vssd1 vssd1 vccd1 vccd1 _26599_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19140_ _19140_/A vssd1 vssd1 vccd1 vccd1 _19472_/B sky130_fd_sc_hd__clkbuf_2
X_16352_ _15111_/X _25783_/Q _15119_/S _26869_/Q _16442_/S vssd1 vssd1 vccd1 vccd1
+ _16352_/X sky130_fd_sc_hd__o221a_1
XFILLER_197_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13564_ _15791_/A _14604_/B _16292_/A vssd1 vssd1 vccd1 vccd1 _13564_/Y sky130_fd_sc_hd__nor3_1
XFILLER_12_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15303_ _16087_/S vssd1 vssd1 vccd1 vccd1 _16086_/S sky130_fd_sc_hd__clkbuf_4
X_19071_ _17299_/X _18559_/X _19067_/X _19070_/X _18574_/X vssd1 vssd1 vccd1 vccd1
+ _19071_/X sky130_fd_sc_hd__o221a_1
X_13495_ _15109_/A _26694_/Q _26822_/Q _13492_/X _13494_/X vssd1 vssd1 vccd1 vccd1
+ _13495_/X sky130_fd_sc_hd__a221o_1
XFILLER_157_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16283_ _20280_/A vssd1 vssd1 vccd1 vccd1 _16283_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18022_ _19253_/A vssd1 vssd1 vccd1 vccd1 _18022_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15234_ _15217_/X _15233_/X _14724_/A vssd1 vssd1 vccd1 vccd1 _15234_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_172_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15165_ _15376_/S vssd1 vssd1 vccd1 vccd1 _15165_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14116_ _27300_/Q _26557_/Q _14176_/S vssd1 vssd1 vccd1 vccd1 _14116_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19973_ _20654_/A _19727_/X _19972_/X _18016_/A vssd1 vssd1 vccd1 vccd1 _20006_/B
+ sky130_fd_sc_hd__a2bb2oi_1
X_15096_ _25823_/Q _27257_/Q _16422_/S vssd1 vssd1 vccd1 vccd1 _15096_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18924_ _18435_/A _18923_/X _18912_/B vssd1 vssd1 vccd1 vccd1 _18924_/X sky130_fd_sc_hd__a21o_1
X_14047_ _14047_/A vssd1 vssd1 vccd1 vccd1 _14390_/S sky130_fd_sc_hd__buf_2
XFILLER_262_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18855_ _18855_/A _18855_/B _18855_/C vssd1 vssd1 vccd1 vccd1 _18855_/Y sky130_fd_sc_hd__nand3_2
XFILLER_268_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17806_ _17941_/A _14562_/B vssd1 vssd1 vccd1 vccd1 _18251_/B sky130_fd_sc_hd__or2b_1
XFILLER_283_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18786_ _19449_/A vssd1 vssd1 vccd1 vccd1 _19042_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_283_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15998_ _26632_/Q _26728_/Q _16020_/S vssd1 vssd1 vccd1 vccd1 _15999_/B sky130_fd_sc_hd__mux2_1
XFILLER_36_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17737_ _17762_/A _17762_/B _17747_/C vssd1 vssd1 vccd1 vccd1 _18119_/A sky130_fd_sc_hd__or3_1
XFILLER_76_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14949_ _14944_/X _14948_/X _16221_/S vssd1 vssd1 vccd1 vccd1 _14949_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17668_ _18138_/A vssd1 vssd1 vccd1 vccd1 _17769_/A sky130_fd_sc_hd__inv_2
XINSDIODE2_120 _23047_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_131 _17992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_142 _14228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19407_ _18742_/X _19397_/X _19406_/X vssd1 vssd1 vccd1 vccd1 _19407_/X sky130_fd_sc_hd__a21o_4
XINSDIODE2_153 _23542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16619_ _16625_/A _16626_/B _18938_/S vssd1 vssd1 vccd1 vccd1 _18975_/A sky130_fd_sc_hd__o21ai_4
XFILLER_62_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_164 _13585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17599_ _14773_/X _17551_/X _17553_/X _17598_/X vssd1 vssd1 vccd1 vccd1 _17600_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_126_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_175 _16419_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_186 _19800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19338_ _25560_/Q _18568_/X _19337_/X _19069_/X _18572_/X vssd1 vssd1 vccd1 vccd1
+ _19338_/X sky130_fd_sc_hd__a221o_1
XFILLER_206_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_197 _19700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19269_ _18435_/X _19267_/X _19268_/Y vssd1 vssd1 vccd1 vccd1 _19271_/B sky130_fd_sc_hd__a21oi_1
XFILLER_164_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21300_ _21300_/A _21332_/B vssd1 vssd1 vccd1 vccd1 _21300_/X sky130_fd_sc_hd__or2_1
XFILLER_276_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22280_ _26205_/Q _22279_/X _22270_/X _26306_/Q _22271_/X vssd1 vssd1 vccd1 vccd1
+ _22280_/X sky130_fd_sc_hd__a221o_1
XFILLER_163_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21231_ _21271_/A vssd1 vssd1 vccd1 vccd1 _21231_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_3_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_145_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21162_ _21162_/A vssd1 vssd1 vccd1 vccd1 _25925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_278_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20113_ _22507_/A _20151_/C vssd1 vssd1 vccd1 vccd1 _20113_/X sky130_fd_sc_hd__xor2_1
XFILLER_131_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25970_ _27156_/CLK _25970_/D vssd1 vssd1 vccd1 vccd1 _25970_/Q sky130_fd_sc_hd__dfxtp_1
X_21093_ _21093_/A vssd1 vssd1 vccd1 vccd1 _25906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24921_ _25221_/A vssd1 vssd1 vccd1 vccd1 _24921_/X sky130_fd_sc_hd__clkbuf_2
X_20044_ _20098_/C _20031_/Y _19941_/X _20043_/X vssd1 vssd1 vccd1 vccd1 _20044_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_131_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24852_ _27119_/Q _24856_/B vssd1 vssd1 vccd1 vccd1 _24852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23803_ _23803_/A vssd1 vssd1 vccd1 vccd1 _26785_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ _21995_/A vssd1 vssd1 vccd1 vccd1 _26110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24783_ _20624_/A _19642_/X _24781_/Y _24782_/X vssd1 vssd1 vccd1 vccd1 _24783_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26522_ _27297_/CLK _26522_/D vssd1 vssd1 vccd1 vccd1 _26522_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23734_ _23734_/A vssd1 vssd1 vccd1 vccd1 _23734_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_198_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20946_ _25852_/Q _20945_/X _20949_/S vssd1 vssd1 vccd1 vccd1 _20947_/A sky130_fd_sc_hd__mux2_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26453_ _26453_/CLK _26453_/D vssd1 vssd1 vccd1 vccd1 _26453_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20877_ _20877_/A vssd1 vssd1 vccd1 vccd1 _25830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23665_ _26739_/Q _23584_/X _23667_/S vssd1 vssd1 vccd1 vccd1 _23666_/A sky130_fd_sc_hd__mux2_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25404_ _23699_/X _27299_/Q _25404_/S vssd1 vssd1 vccd1 vccd1 _25405_/A sky130_fd_sc_hd__mux2_1
X_22616_ _26321_/Q _22618_/B vssd1 vssd1 vccd1 vccd1 _22616_/Y sky130_fd_sc_hd__nand2_1
X_23596_ _23596_/A vssd1 vssd1 vccd1 vccd1 _26710_/D sky130_fd_sc_hd__clkbuf_1
X_26384_ _27287_/CLK _26384_/D vssd1 vssd1 vccd1 vccd1 _26384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25335_ _27268_/Q _23702_/A _25343_/S vssd1 vssd1 vccd1 vccd1 _25336_/A sky130_fd_sc_hd__mux2_1
X_22547_ _22600_/A vssd1 vssd1 vccd1 vccd1 _22547_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_220_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13280_ _15576_/A vssd1 vssd1 vccd1 vccd1 _13281_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_212_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25266_ _25266_/A vssd1 vssd1 vccd1 vccd1 _27237_/D sky130_fd_sc_hd__clkbuf_1
X_22478_ _22478_/A _22480_/B vssd1 vssd1 vccd1 vccd1 _22479_/A sky130_fd_sc_hd__and2_1
XFILLER_154_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27005_ _27137_/CLK _27005_/D vssd1 vssd1 vccd1 vccd1 _27005_/Q sky130_fd_sc_hd__dfxtp_1
X_24217_ _26962_/Q _24215_/B _24216_/Y vssd1 vssd1 vccd1 vccd1 _26962_/D sky130_fd_sc_hd__o21a_1
X_21429_ _21429_/A _21495_/B vssd1 vssd1 vccd1 vccd1 _21429_/X sky130_fd_sc_hd__or2_1
X_25197_ _24686_/B _25189_/X _25196_/X _27209_/Q _25191_/X vssd1 vssd1 vccd1 vccd1
+ _27209_/D sky130_fd_sc_hd__o221a_1
XFILLER_5_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24148_ _27327_/Q _17224_/A _18028_/A _20707_/C _20487_/A vssd1 vssd1 vccd1 vccd1
+ _24148_/X sky130_fd_sc_hd__a41o_1
XFILLER_269_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24079_ _26908_/Q _23508_/X _24087_/S vssd1 vssd1 vccd1 vccd1 _24080_/A sky130_fd_sc_hd__mux2_1
X_16970_ _16980_/A _16970_/B _16970_/C vssd1 vssd1 vccd1 vccd1 _16971_/A sky130_fd_sc_hd__and3_2
XFILLER_122_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15921_ _15921_/A _15921_/B vssd1 vssd1 vccd1 vccd1 _15921_/Y sky130_fd_sc_hd__nor2_2
XFILLER_49_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18640_ _17920_/X _18210_/X _18639_/X vssd1 vssd1 vccd1 vccd1 _18640_/X sky130_fd_sc_hd__a21o_1
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15852_ _15852_/A _15852_/B vssd1 vssd1 vccd1 vccd1 _15852_/X sky130_fd_sc_hd__or2_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _14803_/A vssd1 vssd1 vccd1 vccd1 _14804_/A sky130_fd_sc_hd__clkbuf_4
X_18571_ _26949_/Q _18569_/X _18570_/X _26981_/Q vssd1 vssd1 vccd1 vccd1 _18571_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _13466_/A _15766_/Y _15782_/Y _14827_/A vssd1 vssd1 vccd1 vccd1 _15783_/Y
+ sky130_fd_sc_hd__a31oi_4
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12995_ _20488_/A _14518_/S _13139_/A _13197_/A _12994_/X vssd1 vssd1 vccd1 vccd1
+ _13005_/A sky130_fd_sc_hd__a221o_1
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _25176_/A vssd1 vssd1 vccd1 vccd1 _24277_/A sky130_fd_sc_hd__clkbuf_16
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14734_ _16189_/S vssd1 vssd1 vccd1 vccd1 _15209_/S sky130_fd_sc_hd__clkbuf_4
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17453_ _17453_/A vssd1 vssd1 vccd1 vccd1 _17454_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_189_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14665_ _16163_/S vssd1 vssd1 vccd1 vccd1 _16134_/S sky130_fd_sc_hd__buf_2
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16404_ _15044_/X _16402_/X _16403_/X vssd1 vssd1 vccd1 vccd1 _16405_/B sky130_fd_sc_hd__o21ai_1
X_13616_ _26529_/Q _26137_/Q _13616_/S vssd1 vssd1 vccd1 vccd1 _13616_/X sky130_fd_sc_hd__mux2_1
X_17384_ _25547_/Q vssd1 vssd1 vccd1 vccd1 _17384_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_220_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14596_ _14596_/A vssd1 vssd1 vccd1 vccd1 _14597_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19123_ _19123_/A _19123_/B vssd1 vssd1 vccd1 vccd1 _19579_/C sky130_fd_sc_hd__xnor2_2
X_16335_ _25749_/Q vssd1 vssd1 vccd1 vccd1 _20690_/A sky130_fd_sc_hd__clkinv_4
X_13547_ _14786_/A _13497_/X _13506_/X _14722_/A _13546_/X vssd1 vssd1 vccd1 vccd1
+ _13547_/X sky130_fd_sc_hd__a311o_4
XFILLER_200_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19054_ _17299_/X _18556_/X _18557_/X _25552_/Q vssd1 vssd1 vccd1 vccd1 _19054_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16266_ _14807_/A _16254_/X _16258_/X _16265_/X vssd1 vssd1 vccd1 vccd1 _16266_/X
+ sky130_fd_sc_hd__a31o_1
X_13478_ _13939_/A vssd1 vssd1 vccd1 vccd1 _13479_/A sky130_fd_sc_hd__clkbuf_4
X_18005_ _18005_/A _19003_/A _18005_/C _18004_/X vssd1 vssd1 vccd1 vccd1 _18005_/X
+ sky130_fd_sc_hd__or4b_1
X_15217_ _16350_/A _15217_/B vssd1 vssd1 vccd1 vccd1 _15217_/X sky130_fd_sc_hd__or2_1
Xoutput305 _16689_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[0] sky130_fd_sc_hd__buf_2
X_16197_ _15110_/A _26609_/Q _15299_/S _26349_/Q _15606_/X vssd1 vssd1 vccd1 vccd1
+ _16197_/X sky130_fd_sc_hd__o221a_1
XFILLER_154_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput316 _16691_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[1] sky130_fd_sc_hd__buf_2
XFILLER_154_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput327 _16715_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[4] sky130_fd_sc_hd__buf_2
XFILLER_154_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput338 _16876_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[13] sky130_fd_sc_hd__buf_2
X_15148_ _16073_/B vssd1 vssd1 vccd1 vccd1 _16154_/B sky130_fd_sc_hd__buf_2
Xoutput349 _16936_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[23] sky130_fd_sc_hd__buf_2
XFILLER_273_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_9_0_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_9_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15079_ _15079_/A _15079_/B _15079_/C vssd1 vssd1 vccd1 vccd1 _15079_/X sky130_fd_sc_hd__or3_4
X_19956_ _19957_/A _19957_/B vssd1 vssd1 vccd1 vccd1 _19956_/X sky130_fd_sc_hd__or2_1
XFILLER_45_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18907_ _18932_/B _19049_/A vssd1 vssd1 vccd1 vccd1 _18907_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19887_ _19887_/A _19887_/B vssd1 vssd1 vccd1 vccd1 _19918_/B sky130_fd_sc_hd__nor2_1
XFILLER_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18838_ _18838_/A _18838_/B vssd1 vssd1 vccd1 vccd1 _18848_/B sky130_fd_sc_hd__xnor2_4
Xclkbuf_leaf_109_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25545_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_95_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18769_ _25545_/Q _18763_/X _18766_/X _18767_/X _18768_/X vssd1 vssd1 vccd1 vccd1
+ _18769_/X sky130_fd_sc_hd__a221o_1
XFILLER_215_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20800_ _22368_/A _20800_/B vssd1 vssd1 vccd1 vccd1 _20801_/A sky130_fd_sc_hd__and2_1
XFILLER_35_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21780_ _21780_/A vssd1 vssd1 vccd1 vccd1 _26022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20731_ _20512_/X _25763_/Q _20739_/S vssd1 vssd1 vccd1 vccd1 _20732_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23450_ _26657_/Q _23053_/X _23458_/S vssd1 vssd1 vccd1 vccd1 _23451_/A sky130_fd_sc_hd__mux2_1
X_20662_ _20662_/A _20670_/B vssd1 vssd1 vccd1 vccd1 _20662_/X sky130_fd_sc_hd__or2_1
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22401_ _22361_/B _22395_/B _22379_/A vssd1 vssd1 vccd1 vccd1 _22401_/X sky130_fd_sc_hd__a21bo_1
XFILLER_52_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23381_ _23381_/A vssd1 vssd1 vccd1 vccd1 _26626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20593_ _20592_/X _25716_/Q _20593_/S vssd1 vssd1 vccd1 vccd1 _20594_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22332_ _26223_/Q _22154_/A _22270_/A _26324_/Q _22271_/A vssd1 vssd1 vccd1 vccd1
+ _22332_/X sky130_fd_sc_hd__a221o_1
X_25120_ _22516_/A _25119_/X _25114_/X _16638_/B _25106_/X vssd1 vssd1 vccd1 vccd1
+ _25120_/X sky130_fd_sc_hd__a221o_1
XFILLER_149_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25051_ _27175_/Q _25030_/X _25050_/X vssd1 vssd1 vccd1 vccd1 _27175_/D sky130_fd_sc_hd__o21ba_1
X_22263_ _26200_/Q _22254_/X _22262_/X _22258_/X vssd1 vssd1 vccd1 vccd1 _26200_/D
+ sky130_fd_sc_hd__o211a_1
X_24002_ _26875_/Q _23609_/X _24002_/S vssd1 vssd1 vccd1 vccd1 _24003_/A sky130_fd_sc_hd__mux2_1
X_21214_ _21214_/A _21214_/B vssd1 vssd1 vccd1 vccd1 _21221_/B sky130_fd_sc_hd__or2_1
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22194_ _26182_/Q _22186_/X _22179_/A input266/X _22187_/X vssd1 vssd1 vccd1 vccd1
+ _22194_/X sky130_fd_sc_hd__a221o_1
XFILLER_279_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21145_ _25921_/Q _21130_/X _21131_/X input20/X vssd1 vssd1 vccd1 vccd1 _21146_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_105_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25953_ _25992_/CLK _25953_/D vssd1 vssd1 vccd1 vccd1 _25953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21076_ _21167_/A vssd1 vssd1 vccd1 vccd1 _21113_/A sky130_fd_sc_hd__buf_4
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24904_ _24954_/A vssd1 vssd1 vccd1 vccd1 _24978_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_19_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20027_ _19649_/A _20024_/Y _20025_/X _20026_/X vssd1 vssd1 vccd1 vccd1 _20027_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_219_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25884_ _27281_/CLK _25884_/D vssd1 vssd1 vccd1 vccd1 _25884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24835_ _24835_/A vssd1 vssd1 vccd1 vccd1 _24835_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _25106_/A vssd1 vssd1 vccd1 vccd1 _25024_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24766_ _20478_/A _24636_/A _25159_/A _24660_/X vssd1 vssd1 vccd1 vccd1 _24767_/B
+ sky130_fd_sc_hd__o22a_1
X_21978_ _21978_/A vssd1 vssd1 vccd1 vccd1 _26102_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26505_ _27280_/CLK _26505_/D vssd1 vssd1 vccd1 vccd1 _26505_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23717_ _23717_/A vssd1 vssd1 vccd1 vccd1 _26757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20929_ _23744_/A vssd1 vssd1 vccd1 vccd1 _20929_/X sky130_fd_sc_hd__clkbuf_2
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24697_ _24720_/A vssd1 vssd1 vccd1 vccd1 _24697_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26436_ _26468_/CLK _26436_/D vssd1 vssd1 vccd1 vccd1 _26436_/Q sky130_fd_sc_hd__dfxtp_2
X_14450_ _26065_/Q _14307_/S _14449_/X _14043_/X vssd1 vssd1 vccd1 vccd1 _14450_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_214_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23648_ _26731_/Q _23558_/X _23656_/S vssd1 vssd1 vccd1 vccd1 _23649_/A sky130_fd_sc_hd__mux2_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13401_ _25608_/Q _12981_/A _13398_/Y _13400_/X vssd1 vssd1 vccd1 vccd1 _23542_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_168_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26367_ _26433_/CLK _26367_/D vssd1 vssd1 vccd1 vccd1 _26367_/Q sky130_fd_sc_hd__dfxtp_1
X_14381_ _13520_/A _26686_/Q _26814_/Q _14391_/S _12731_/A vssd1 vssd1 vccd1 vccd1
+ _14381_/X sky130_fd_sc_hd__a221o_1
XFILLER_183_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23579_ _26705_/Q _23578_/X _23588_/S vssd1 vssd1 vccd1 vccd1 _23580_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16120_ _14789_/A _23571_/A _16119_/Y _15127_/A vssd1 vssd1 vccd1 vccd1 _20168_/A
+ sky130_fd_sc_hd__o211ai_4
X_13332_ _13821_/A vssd1 vssd1 vccd1 vccd1 _15932_/A sky130_fd_sc_hd__buf_2
X_25318_ _25318_/A vssd1 vssd1 vccd1 vccd1 _27261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_259_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26298_ _26327_/CLK _26298_/D vssd1 vssd1 vccd1 vccd1 _26298_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16051_ _15167_/A _26411_/Q _15141_/A _16050_/X vssd1 vssd1 vccd1 vccd1 _16051_/X
+ sky130_fd_sc_hd__o211a_1
X_13263_ _15322_/A vssd1 vssd1 vccd1 vccd1 _16341_/S sky130_fd_sc_hd__buf_4
X_25249_ _25249_/A _25249_/B _25249_/C vssd1 vssd1 vccd1 vccd1 _25306_/A sky130_fd_sc_hd__or3_4
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15002_ _26092_/Q _25897_/Q _15003_/S vssd1 vssd1 vccd1 vccd1 _15002_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13194_ _14458_/S vssd1 vssd1 vccd1 vccd1 _13244_/A sky130_fd_sc_hd__buf_4
XFILLER_29_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19810_ _19926_/A vssd1 vssd1 vccd1 vccd1 _20208_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_7_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26929_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_285_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19741_ _25663_/Q _25662_/Q _25664_/Q vssd1 vssd1 vccd1 vccd1 _19741_/Y sky130_fd_sc_hd__a21oi_1
X_16953_ _15079_/X _16952_/X _16834_/A vssd1 vssd1 vccd1 vccd1 _16959_/B sky130_fd_sc_hd__o21ai_2
XFILLER_110_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15904_ _26501_/Q _26373_/Q _15904_/S vssd1 vssd1 vccd1 vccd1 _15904_/X sky130_fd_sc_hd__mux2_1
XFILLER_277_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19672_ _12722_/B _19589_/A _20092_/B _25574_/Q vssd1 vssd1 vccd1 vccd1 _19673_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_238_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16884_ _16855_/A _16882_/X _16883_/X _16842_/A vssd1 vssd1 vccd1 vccd1 _16885_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_264_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18623_ _19140_/A _19882_/A vssd1 vssd1 vccd1 vccd1 _18623_/X sky130_fd_sc_hd__and2b_1
X_15835_ _26634_/Q _26730_/Q _15857_/S vssd1 vssd1 vccd1 vccd1 _15836_/B sky130_fd_sc_hd__mux2_1
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18554_ _18554_/A vssd1 vssd1 vccd1 vccd1 _18554_/X sky130_fd_sc_hd__clkbuf_2
X_15766_ _15754_/X _15757_/X _15765_/X vssd1 vssd1 vccd1 vccd1 _15766_/Y sky130_fd_sc_hd__o21ai_2
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12978_ _25641_/Q _16212_/B _14401_/B _25609_/Q _14616_/A vssd1 vssd1 vccd1 vccd1
+ _12978_/X sky130_fd_sc_hd__a221o_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _17662_/A _17662_/B vssd1 vssd1 vccd1 vccd1 _19603_/A sky130_fd_sc_hd__nor2_1
XFILLER_233_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14717_ _25596_/Q _16170_/A _14833_/A vssd1 vssd1 vccd1 vccd1 _14718_/A sky130_fd_sc_hd__a21oi_1
X_18485_ _18485_/A _18345_/S vssd1 vssd1 vccd1 vccd1 _18485_/X sky130_fd_sc_hd__or2b_1
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15697_ _14789_/A _23562_/A _15696_/Y _15127_/A vssd1 vssd1 vccd1 vccd1 _18946_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17436_ _25562_/Q _17430_/B _17435_/Y vssd1 vssd1 vccd1 vccd1 _25562_/D sky130_fd_sc_hd__o21a_1
XFILLER_21_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14648_ _15019_/A vssd1 vssd1 vccd1 vccd1 _14649_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17367_ _17365_/X _17370_/C _17366_/X vssd1 vssd1 vccd1 vccd1 _17367_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_220_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14579_ _18686_/A _14579_/B vssd1 vssd1 vccd1 vccd1 _18678_/A sky130_fd_sc_hd__xor2_4
XFILLER_174_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19106_ _18861_/X _19105_/X _15439_/B vssd1 vssd1 vccd1 vccd1 _19106_/Y sky130_fd_sc_hd__a21oi_2
X_16318_ _26545_/Q _26153_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _16318_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17298_ _25519_/Q _17296_/B _17297_/Y vssd1 vssd1 vccd1 vccd1 _25519_/D sky130_fd_sc_hd__o21a_1
XFILLER_284_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19037_ _25742_/Q _25741_/Q _19037_/C vssd1 vssd1 vccd1 vccd1 _19081_/B sky130_fd_sc_hd__and3_1
XFILLER_118_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16249_ _16463_/A _23584_/A _16248_/X _15388_/X vssd1 vssd1 vccd1 vccd1 _16932_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_173_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19939_ _25671_/Q _19985_/C vssd1 vssd1 vccd1 vccd1 _20017_/C sky130_fd_sc_hd__and2_1
XFILLER_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22950_ _26450_/Q _22727_/X _22956_/S vssd1 vssd1 vccd1 vccd1 _22951_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21901_ _21901_/A vssd1 vssd1 vccd1 vccd1 _26068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_255_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22881_ _22881_/A vssd1 vssd1 vccd1 vccd1 _26419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24620_ _27063_/Q _24615_/X _24618_/Y _24619_/X vssd1 vssd1 vccd1 vccd1 _27063_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21832_ _26045_/Q _20923_/X _21838_/S vssd1 vssd1 vccd1 vccd1 _21833_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24551_ _24551_/A vssd1 vssd1 vccd1 vccd1 _24551_/X sky130_fd_sc_hd__clkbuf_2
X_21763_ _20567_/X _26015_/Q _21765_/S vssd1 vssd1 vccd1 vccd1 _21764_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23502_ _26681_/Q _23130_/X _23502_/S vssd1 vssd1 vccd1 vccd1 _23503_/A sky130_fd_sc_hd__mux2_1
X_20714_ _20709_/Y _20712_/X _24770_/A vssd1 vssd1 vccd1 vccd1 _25757_/D sky130_fd_sc_hd__a21oi_1
X_27270_ _27272_/CLK _27270_/D vssd1 vssd1 vccd1 vccd1 _27270_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_77_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26593_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21694_ _25986_/Q input198/X _21696_/S vssd1 vssd1 vccd1 vccd1 _21695_/A sky130_fd_sc_hd__mux2_1
X_24482_ _24454_/X _25618_/Q _24481_/X vssd1 vssd1 vccd1 vccd1 _24960_/A sky130_fd_sc_hd__o21ai_4
XFILLER_169_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26221_ _26222_/CLK _26221_/D vssd1 vssd1 vccd1 vccd1 _26221_/Q sky130_fd_sc_hd__dfxtp_1
X_20645_ _26269_/Q _20633_/X _20643_/X _20644_/X vssd1 vssd1 vccd1 vccd1 _25732_/D
+ sky130_fd_sc_hd__o211a_1
X_23433_ _23433_/A vssd1 vssd1 vccd1 vccd1 _26650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26152_ _27329_/A _26152_/D vssd1 vssd1 vccd1 vccd1 _26152_/Q sky130_fd_sc_hd__dfxtp_1
X_23364_ _25393_/A _23860_/B vssd1 vssd1 vccd1 vccd1 _23421_/A sky130_fd_sc_hd__nor2_4
XFILLER_164_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20576_ _20597_/A vssd1 vssd1 vccd1 vccd1 _20593_/S sky130_fd_sc_hd__buf_4
XFILLER_176_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25103_ _20670_/A _25086_/X _25102_/X vssd1 vssd1 vccd1 vccd1 _25103_/Y sky130_fd_sc_hd__o21ai_1
X_22315_ _22315_/A vssd1 vssd1 vccd1 vccd1 _22315_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23295_ _23295_/A vssd1 vssd1 vccd1 vccd1 _26588_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26083_ _27282_/CLK _26083_/D vssd1 vssd1 vccd1 vccd1 _26083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22246_ _26194_/Q _22235_/X _22245_/X _22243_/X vssd1 vssd1 vccd1 vccd1 _26194_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_219_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25034_ _25665_/Q _25015_/X _25033_/X _18357_/A _25024_/X vssd1 vssd1 vccd1 vccd1
+ _25034_/X sky130_fd_sc_hd__a221o_1
XFILLER_152_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22177_ _26176_/Q _22171_/X _22160_/X input275/X _22172_/X vssd1 vssd1 vccd1 vccd1
+ _22177_/X sky130_fd_sc_hd__a221o_1
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21128_ _21136_/A _21128_/B vssd1 vssd1 vccd1 vccd1 _21129_/A sky130_fd_sc_hd__or2_1
XFILLER_78_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26985_ _26987_/CLK _26985_/D vssd1 vssd1 vccd1 vccd1 _26985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13950_ _13484_/A _13948_/X _13949_/X _13945_/X vssd1 vssd1 vccd1 vccd1 _13954_/B
+ sky130_fd_sc_hd__o211a_1
X_25936_ _27156_/CLK _25936_/D vssd1 vssd1 vccd1 vccd1 _25936_/Q sky130_fd_sc_hd__dfxtp_1
X_21059_ _25898_/Q _20964_/X _21059_/S vssd1 vssd1 vccd1 vccd1 _21060_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12901_ _12915_/A vssd1 vssd1 vccd1 vccd1 _12902_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13881_ _26627_/Q _26723_/Q _14008_/S vssd1 vssd1 vccd1 vccd1 _13881_/X sky130_fd_sc_hd__mux2_1
X_25867_ _25867_/CLK _25867_/D vssd1 vssd1 vccd1 vccd1 _25867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15620_ _14600_/A _15618_/Y _15619_/X _15135_/A vssd1 vssd1 vccd1 vccd1 _15620_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12832_ _12862_/A _12873_/A vssd1 vssd1 vccd1 vccd1 _13916_/A sky130_fd_sc_hd__nor2_2
X_24818_ _27110_/Q _24818_/B vssd1 vssd1 vccd1 vccd1 _24818_/Y sky130_fd_sc_hd__nand2_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25798_ _26520_/CLK _25798_/D vssd1 vssd1 vccd1 vccd1 _25798_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15551_ _16079_/S _15548_/X _15550_/X _15039_/A vssd1 vssd1 vccd1 vccd1 _15551_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12763_ _17444_/C _12778_/B vssd1 vssd1 vccd1 vccd1 _12763_/Y sky130_fd_sc_hd__nor2_8
X_24749_ _24749_/A vssd1 vssd1 vccd1 vccd1 _24781_/A sky130_fd_sc_hd__buf_4
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _15979_/S _14496_/X _14498_/X _14501_/X _14440_/S vssd1 vssd1 vccd1 vccd1
+ _14502_/X sky130_fd_sc_hd__o311a_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18270_ _18348_/S _17894_/X _17981_/Y vssd1 vssd1 vccd1 vccd1 _18270_/X sky130_fd_sc_hd__o21a_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _15482_/A _16901_/A vssd1 vssd1 vccd1 vccd1 _15482_/Y sky130_fd_sc_hd__nor2_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _25575_/Q _25574_/Q _25573_/Q _25572_/Q vssd1 vssd1 vccd1 vccd1 _17669_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_230_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _25499_/Q _17529_/A _17146_/A _20249_/A vssd1 vssd1 vccd1 vccd1 _17222_/B
+ sky130_fd_sc_hd__a22o_1
X_14433_ _26781_/Q _26425_/Q _14433_/S vssd1 vssd1 vccd1 vccd1 _14433_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26419_ _26903_/CLK _26419_/D vssd1 vssd1 vccd1 vccd1 _26419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17152_ _22817_/B _17151_/X _17146_/X _25575_/Q vssd1 vssd1 vccd1 vccd1 _17153_/B
+ sky130_fd_sc_hd__a22o_1
X_14364_ _14562_/A vssd1 vssd1 vccd1 vccd1 _17941_/A sky130_fd_sc_hd__buf_2
Xinput15 core_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_1
Xinput26 core_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput37 core_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_1
Xinput48 dout0[14] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_2
X_16103_ _26539_/Q _26147_/Q _16176_/S vssd1 vssd1 vccd1 vccd1 _16104_/B sky130_fd_sc_hd__mux2_1
XFILLER_171_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13315_ _13292_/X _13306_/X _13314_/X vssd1 vssd1 vccd1 vccd1 _13315_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_155_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput59 dout0[24] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_2
X_17083_ _17087_/A _17091_/C _17087_/C _17085_/C vssd1 vssd1 vccd1 vccd1 _22239_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_156_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14295_ _13484_/A _14293_/X _14294_/X _13945_/X vssd1 vssd1 vccd1 vccd1 _14299_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16034_ _18686_/A _14579_/B _13381_/Y vssd1 vssd1 vccd1 vccd1 _18726_/B sky130_fd_sc_hd__o21ba_4
XFILLER_115_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13246_ _13779_/A vssd1 vssd1 vccd1 vccd1 _15300_/A sky130_fd_sc_hd__buf_4
XFILLER_6_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13177_ _25568_/Q _25567_/Q _18028_/B vssd1 vssd1 vccd1 vccd1 _18006_/C sky130_fd_sc_hd__nand3b_4
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17985_ _18492_/A _18487_/B _17984_/Y vssd1 vssd1 vccd1 vccd1 _18898_/B sky130_fd_sc_hd__a21oi_2
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19724_ _24749_/A vssd1 vssd1 vccd1 vccd1 _19724_/X sky130_fd_sc_hd__clkbuf_2
X_16936_ _16936_/A vssd1 vssd1 vccd1 vccd1 _16936_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_270_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16867_ _16463_/X _23549_/A _15994_/Y _16860_/B vssd1 vssd1 vccd1 vccd1 _16867_/X
+ sky130_fd_sc_hd__o211a_4
X_19655_ _24641_/A vssd1 vssd1 vccd1 vccd1 _24706_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15818_ _15816_/X _15817_/X _15818_/S vssd1 vssd1 vccd1 vccd1 _15818_/X sky130_fd_sc_hd__mux2_1
X_18606_ _18597_/X _18600_/X _18601_/Y _18602_/X _18605_/X vssd1 vssd1 vccd1 vccd1
+ _18606_/X sky130_fd_sc_hd__o221a_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19586_ _17956_/S _19583_/B _19584_/X _19585_/X vssd1 vssd1 vccd1 vccd1 _19586_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16798_ _16938_/B vssd1 vssd1 vccd1 vccd1 _16842_/A sky130_fd_sc_hd__buf_2
XFILLER_34_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18537_ _18537_/A vssd1 vssd1 vccd1 vccd1 _25605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15749_ _13641_/B _16581_/A _15243_/A _15748_/X vssd1 vssd1 vccd1 vccd1 _17826_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_252_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18468_ _18468_/A vssd1 vssd1 vccd1 vccd1 _18469_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17419_ _17428_/A _17419_/B _17420_/B vssd1 vssd1 vccd1 vccd1 _25557_/D sky130_fd_sc_hd__nor3_1
XFILLER_194_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18399_ _18823_/A vssd1 vssd1 vccd1 vccd1 _18519_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_165_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20430_ _27130_/Q _19691_/X _19905_/A vssd1 vssd1 vccd1 vccd1 _20430_/X sky130_fd_sc_hd__o21a_1
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20361_ _20398_/A _20352_/Y _20354_/X _19833_/A vssd1 vssd1 vccd1 vccd1 _20362_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_146_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22100_ _22100_/A vssd1 vssd1 vccd1 vccd1 _26157_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23080_ _26501_/Q _23079_/X _23083_/S vssd1 vssd1 vccd1 vccd1 _23081_/A sky130_fd_sc_hd__mux2_1
X_20292_ _27156_/Q _27090_/Q vssd1 vssd1 vccd1 vccd1 _20292_/X sky130_fd_sc_hd__or2_1
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_195_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26932_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22031_ _26127_/Q _20970_/X _22031_/S vssd1 vssd1 vccd1 vccd1 _22032_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_124_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27049_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26770_ _26932_/CLK _26770_/D vssd1 vssd1 vccd1 vccd1 _26770_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23982_ _23982_/A vssd1 vssd1 vccd1 vccd1 _26865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_263_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25721_ _27291_/CLK _25721_/D vssd1 vssd1 vccd1 vccd1 _25721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22933_ _22933_/A vssd1 vssd1 vccd1 vccd1 _26442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25652_ _25660_/CLK _25652_/D vssd1 vssd1 vccd1 vccd1 _25652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22864_ _22875_/A vssd1 vssd1 vccd1 vccd1 _22873_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_44_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24603_ _24960_/A _24608_/B vssd1 vssd1 vccd1 vccd1 _24603_/Y sky130_fd_sc_hd__nand2_1
X_21815_ _21815_/A vssd1 vssd1 vccd1 vccd1 _26037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_251_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25583_ _26843_/CLK _25583_/D vssd1 vssd1 vccd1 vccd1 _25583_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22795_ _22795_/A vssd1 vssd1 vccd1 vccd1 _26381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27322_ _27322_/CLK _27322_/D vssd1 vssd1 vccd1 vccd1 _27322_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24534_ _27035_/Q _24372_/A _24533_/Y _24523_/X vssd1 vssd1 vccd1 vccd1 _27035_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21746_ _20533_/X _26007_/Q _21754_/S vssd1 vssd1 vccd1 vccd1 _21747_/A sky130_fd_sc_hd__mux2_1
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27253_ _27253_/CLK _27253_/D vssd1 vssd1 vccd1 vccd1 _27253_/Q sky130_fd_sc_hd__dfxtp_1
X_24465_ _27022_/Q _24448_/X _24464_/Y _24442_/X vssd1 vssd1 vccd1 vccd1 _27022_/D
+ sky130_fd_sc_hd__o211a_1
X_21677_ _25978_/Q input213/X _21685_/S vssd1 vssd1 vccd1 vccd1 _21678_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26204_ _26307_/CLK _26204_/D vssd1 vssd1 vccd1 vccd1 _26204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23416_ _23416_/A vssd1 vssd1 vccd1 vccd1 _26642_/D sky130_fd_sc_hd__clkbuf_1
X_20628_ _20628_/A _20630_/B vssd1 vssd1 vccd1 vccd1 _20628_/X sky130_fd_sc_hd__or2_1
X_27184_ _27188_/CLK _27184_/D vssd1 vssd1 vccd1 vccd1 _27184_/Q sky130_fd_sc_hd__dfxtp_1
X_24396_ _26298_/Q _24393_/X _24394_/X input242/X _24395_/X vssd1 vssd1 vccd1 vccd1
+ _24396_/X sky130_fd_sc_hd__a221o_1
XFILLER_138_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26135_ _26462_/CLK _26135_/D vssd1 vssd1 vccd1 vccd1 _26135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20559_ _23738_/A vssd1 vssd1 vccd1 vccd1 _20559_/X sky130_fd_sc_hd__clkbuf_2
X_23347_ _23347_/A vssd1 vssd1 vccd1 vccd1 _26612_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13100_ _14010_/S vssd1 vssd1 vccd1 vccd1 _15806_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26066_ _26909_/CLK _26066_/D vssd1 vssd1 vccd1 vccd1 _26066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14080_ _25729_/Q _14481_/B vssd1 vssd1 vccd1 vccd1 _14080_/X sky130_fd_sc_hd__or2_1
X_23278_ _23278_/A vssd1 vssd1 vccd1 vccd1 _26581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13031_ _13031_/A vssd1 vssd1 vccd1 vccd1 _15187_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_140_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25017_ _20628_/A _25003_/X _25016_/X vssd1 vssd1 vccd1 vccd1 _25017_/Y sky130_fd_sc_hd__o21ai_1
X_22229_ _26230_/Q vssd1 vssd1 vccd1 vccd1 _22337_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17770_ _18945_/A vssd1 vssd1 vccd1 vccd1 _18383_/A sky130_fd_sc_hd__clkbuf_2
X_26968_ _27000_/CLK _26968_/D vssd1 vssd1 vccd1 vccd1 _26968_/Q sky130_fd_sc_hd__dfxtp_1
X_14982_ _14890_/X _25857_/Q _26057_/Q _14984_/S _14754_/A vssd1 vssd1 vccd1 vccd1
+ _14982_/X sky130_fd_sc_hd__a221o_1
XFILLER_94_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16721_ _22483_/A _16703_/X _16705_/X _18424_/A vssd1 vssd1 vccd1 vccd1 _16721_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_247_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13933_ _13933_/A vssd1 vssd1 vccd1 vccd1 _15443_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25919_ _27087_/CLK _25919_/D vssd1 vssd1 vccd1 vccd1 _25919_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_275_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26899_ _26931_/CLK _26899_/D vssd1 vssd1 vccd1 vccd1 _26899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19440_ _25531_/Q _18746_/X _19437_/X _19439_/X _18770_/X vssd1 vssd1 vccd1 vccd1
+ _19440_/X sky130_fd_sc_hd__o221a_1
XFILLER_207_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16652_ _25679_/Q _25678_/Q _25677_/Q _25676_/Q vssd1 vssd1 vccd1 vccd1 _16654_/C
+ sky130_fd_sc_hd__or4_1
X_13864_ _13431_/X _13859_/X _13861_/X _13863_/X vssd1 vssd1 vccd1 vccd1 _13864_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_505 _21235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_516 _16997_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15603_ _25814_/Q _27248_/Q _15923_/S vssd1 vssd1 vccd1 vccd1 _15604_/B sky130_fd_sc_hd__mux2_1
X_19371_ _25561_/Q _18459_/A _19370_/X _18829_/X _18466_/A vssd1 vssd1 vccd1 vccd1
+ _19371_/X sky130_fd_sc_hd__a221o_1
XINSDIODE2_527 _17040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12815_ _15482_/A vssd1 vssd1 vccd1 vccd1 _15659_/A sky130_fd_sc_hd__clkbuf_2
X_16583_ _17998_/A _16800_/B vssd1 vssd1 vccd1 vccd1 _19571_/B sky130_fd_sc_hd__nor2_4
XFILLER_262_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13795_ _14777_/A _13790_/X _13794_/X _13367_/X vssd1 vssd1 vccd1 vccd1 _13795_/X
+ sky130_fd_sc_hd__o31a_1
XINSDIODE2_538 _17018_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_549 _25816_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18322_ _18324_/B _18309_/X _18312_/Y _18936_/A _18321_/Y vssd1 vssd1 vccd1 vccd1
+ _18322_/X sky130_fd_sc_hd__o221a_1
X_15534_ _25615_/Q _14595_/A _15533_/X _14616_/A vssd1 vssd1 vccd1 vccd1 _23565_/A
+ sky130_fd_sc_hd__o22a_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12746_ _15559_/S vssd1 vssd1 vccd1 vccd1 _16071_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_188_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18253_ _19571_/D _18230_/B _19157_/S vssd1 vssd1 vccd1 vccd1 _18253_/X sky130_fd_sc_hd__mux2_1
X_15465_ _12771_/A _26410_/Q _15460_/S _15464_/X vssd1 vssd1 vccd1 vccd1 _15465_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12677_ _25595_/Q vssd1 vssd1 vccd1 vccd1 _19916_/A sky130_fd_sc_hd__buf_6
X_17204_ _17222_/A _17204_/B vssd1 vssd1 vccd1 vccd1 _17205_/A sky130_fd_sc_hd__and2_1
X_14416_ _25870_/Q _13706_/A _14331_/X _14415_/X vssd1 vssd1 vccd1 vccd1 _14416_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_175_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18184_ _18184_/A _18184_/B _18184_/C vssd1 vssd1 vccd1 vccd1 _18185_/B sky130_fd_sc_hd__nand3_1
XFILLER_191_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15396_ _15321_/X _26704_/Q _26832_/Q _15209_/S _14801_/A vssd1 vssd1 vccd1 vccd1
+ _15396_/X sky130_fd_sc_hd__a221o_1
XFILLER_200_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17135_ _21320_/A _17114_/X _17133_/X _17134_/X vssd1 vssd1 vccd1 vccd1 _25474_/D
+ sky130_fd_sc_hd__o211a_1
X_14347_ _26782_/Q _26426_/Q _14351_/S vssd1 vssd1 vccd1 vccd1 _14347_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17066_ _25974_/Q _17061_/X _16994_/X _17063_/X vssd1 vssd1 vccd1 vccd1 _17066_/X
+ sky130_fd_sc_hd__a22o_4
X_14278_ _15885_/A _14268_/X _14277_/X _14421_/A vssd1 vssd1 vccd1 vccd1 _14278_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16017_ _13835_/X _25841_/Q _26041_/Q _13534_/S _15999_/A vssd1 vssd1 vccd1 vccd1
+ _16017_/X sky130_fd_sc_hd__a221o_1
X_13229_ _26663_/Q _25703_/Q _15422_/S vssd1 vssd1 vccd1 vccd1 _13229_/X sky130_fd_sc_hd__mux2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17968_ _17219_/A _18036_/A _18597_/A vssd1 vssd1 vccd1 vccd1 _17978_/B sky130_fd_sc_hd__and3b_1
XFILLER_97_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19707_ _19881_/A vssd1 vssd1 vccd1 vccd1 _20115_/A sky130_fd_sc_hd__buf_2
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16919_ _16924_/A _16919_/B vssd1 vssd1 vccd1 vccd1 _16920_/A sky130_fd_sc_hd__and2_1
X_17899_ _17842_/B _16035_/B _17933_/S vssd1 vssd1 vccd1 vccd1 _17899_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19638_ _20225_/A vssd1 vssd1 vccd1 vccd1 _19638_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_253_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19569_ _19512_/A _19471_/X _19568_/X _19566_/X vssd1 vssd1 vccd1 vccd1 _25661_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21600_ _21586_/X _19340_/X _21587_/X _25824_/Q _21547_/X vssd1 vssd1 vccd1 vccd1
+ _21600_/X sky130_fd_sc_hd__a221o_1
X_22580_ _22606_/A vssd1 vssd1 vccd1 vccd1 _22580_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_240_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21531_ _21597_/A vssd1 vssd1 vccd1 vccd1 _21531_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_194_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24250_ _26973_/Q _26972_/Q _24250_/C vssd1 vssd1 vccd1 vccd1 _24252_/B sky130_fd_sc_hd__and3_1
X_21462_ _25864_/Q vssd1 vssd1 vccd1 vccd1 _21462_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_193_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23201_ _26547_/Q _23124_/X _23205_/S vssd1 vssd1 vccd1 vccd1 _23202_/A sky130_fd_sc_hd__mux2_1
X_20413_ _20413_/A _20412_/Y vssd1 vssd1 vccd1 vccd1 _20415_/A sky130_fd_sc_hd__or2b_1
X_24181_ _26951_/Q _24184_/C vssd1 vssd1 vccd1 vccd1 _24183_/A sky130_fd_sc_hd__and2_1
XFILLER_193_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21393_ _20652_/A _21343_/X _21350_/X _21392_/X vssd1 vssd1 vccd1 vccd1 _21393_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23132_ _23132_/A vssd1 vssd1 vccd1 vccd1 _26517_/D sky130_fd_sc_hd__clkbuf_1
X_20344_ _27158_/Q _20343_/Y _20371_/S vssd1 vssd1 vccd1 vccd1 _20344_/X sky130_fd_sc_hd__mux2_2
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23063_ _23536_/A vssd1 vssd1 vccd1 vccd1 _23063_/X sky130_fd_sc_hd__clkbuf_2
X_20275_ _22518_/A _20225_/X _20267_/X _20274_/Y _20223_/X vssd1 vssd1 vccd1 vccd1
+ _25682_/D sky130_fd_sc_hd__o221a_1
XFILLER_255_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22014_ _26119_/Q _20945_/X _22016_/S vssd1 vssd1 vccd1 vccd1 _22015_/A sky130_fd_sc_hd__mux2_1
XFILLER_276_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput205 localMemory_wb_adr_i[23] vssd1 vssd1 vccd1 vccd1 _21235_/A sky130_fd_sc_hd__buf_4
XTAP_5416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput216 localMemory_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input216/X sky130_fd_sc_hd__buf_6
XFILLER_89_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput227 localMemory_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 input227/X sky130_fd_sc_hd__buf_6
X_26822_ _26856_/CLK _26822_/D vssd1 vssd1 vccd1 vccd1 _26822_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_124_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput238 localMemory_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 input238/X sky130_fd_sc_hd__buf_8
XTAP_5449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput249 localMemory_wb_sel_i[2] vssd1 vssd1 vccd1 vccd1 input249/X sky130_fd_sc_hd__clkbuf_1
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26753_ _26880_/CLK _26753_/D vssd1 vssd1 vccd1 vccd1 _26753_/Q sky130_fd_sc_hd__dfxtp_2
X_23965_ _26858_/Q _23555_/X _23965_/S vssd1 vssd1 vccd1 vccd1 _23966_/A sky130_fd_sc_hd__mux2_1
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25704_ _27307_/CLK _25704_/D vssd1 vssd1 vccd1 vccd1 _25704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22916_ _22916_/A vssd1 vssd1 vccd1 vccd1 _26434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_92_wb_clk_i _25501_/CLK vssd1 vssd1 vccd1 vccd1 _26248_/CLK sky130_fd_sc_hd__clkbuf_16
X_26684_ _26684_/CLK _26684_/D vssd1 vssd1 vccd1 vccd1 _26684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23896_ _23734_/X _26827_/Q _23904_/S vssd1 vssd1 vccd1 vccd1 _23897_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25635_ _26297_/CLK _25635_/D vssd1 vssd1 vccd1 vccd1 _25635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22847_ _26404_/Q _22682_/X _22851_/S vssd1 vssd1 vccd1 vccd1 _22848_/A sky130_fd_sc_hd__mux2_1
XFILLER_271_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27288_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_17_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _16639_/A _13576_/X _13579_/X vssd1 vssd1 vccd1 vccd1 _23539_/A sky130_fd_sc_hd__a21o_4
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25566_ _25590_/CLK _25566_/D vssd1 vssd1 vccd1 vccd1 _25566_/Q sky130_fd_sc_hd__dfxtp_1
X_22778_ _26374_/Q _22688_/X _22778_/S vssd1 vssd1 vccd1 vccd1 _22779_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27305_ _27305_/CLK _27305_/D vssd1 vssd1 vccd1 vccd1 _27305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24517_ _24758_/B vssd1 vssd1 vccd1 vccd1 _24621_/A sky130_fd_sc_hd__inv_2
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21729_ _21729_/A vssd1 vssd1 vccd1 vccd1 _25999_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25497_ _26940_/CLK _25497_/D vssd1 vssd1 vccd1 vccd1 _25497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27236_ _27301_/CLK _27236_/D vssd1 vssd1 vccd1 vccd1 _27236_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15250_ _23581_/A vssd1 vssd1 vccd1 vccd1 _15250_/Y sky130_fd_sc_hd__inv_2
X_24448_ _24506_/A vssd1 vssd1 vccd1 vccd1 _24448_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14201_ _26624_/Q _26720_/Q _15292_/A vssd1 vssd1 vccd1 vccd1 _14201_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15181_ _25853_/Q _26053_/Q _16400_/S vssd1 vssd1 vccd1 vccd1 _15181_/X sky130_fd_sc_hd__mux2_1
X_27167_ _27173_/CLK _27167_/D vssd1 vssd1 vccd1 vccd1 _27167_/Q sky130_fd_sc_hd__dfxtp_2
X_24379_ _24415_/A vssd1 vssd1 vccd1 vccd1 _24379_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_193_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14132_ input119/X input154/X _14132_/S vssd1 vssd1 vccd1 vccd1 _14133_/B sky130_fd_sc_hd__mux2_8
XFILLER_165_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26118_ _26611_/CLK _26118_/D vssd1 vssd1 vccd1 vccd1 _26118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27098_ _27228_/CLK _27098_/D vssd1 vssd1 vccd1 vccd1 _27098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14063_ _14473_/S _14061_/X _14062_/X _13477_/A vssd1 vssd1 vccd1 vccd1 _14069_/B
+ sky130_fd_sc_hd__o211a_1
X_18940_ _18940_/A _18940_/B vssd1 vssd1 vccd1 vccd1 _18940_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26049_ _27283_/CLK _26049_/D vssd1 vssd1 vccd1 vccd1 _26049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13014_ _14272_/S vssd1 vssd1 vccd1 vccd1 _13431_/A sky130_fd_sc_hd__buf_2
X_18871_ _27019_/Q _18756_/X _18870_/X _18821_/X vssd1 vssd1 vccd1 vccd1 _18871_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_267_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17822_ _18676_/B vssd1 vssd1 vccd1 vccd1 _17822_/Y sky130_fd_sc_hd__inv_2
XFILLER_227_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14965_ _25825_/Q _14692_/S _14952_/S _14964_/X vssd1 vssd1 vccd1 vccd1 _14965_/X
+ sky130_fd_sc_hd__o211a_1
X_17753_ _17753_/A _18108_/B vssd1 vssd1 vccd1 vccd1 _18391_/A sky130_fd_sc_hd__and2_1
XFILLER_207_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13916_ _13916_/A _13916_/B _13916_/C _13916_/D vssd1 vssd1 vccd1 vccd1 _14323_/B
+ sky130_fd_sc_hd__and4_1
X_16704_ _16951_/A vssd1 vssd1 vccd1 vccd1 _16770_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17684_ _21214_/B _17684_/B vssd1 vssd1 vccd1 vccd1 _17685_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14896_ _16262_/S vssd1 vssd1 vccd1 vccd1 _16359_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_262_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_302 _26368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19423_ _25161_/A _19423_/B vssd1 vssd1 vccd1 vccd1 _19423_/X sky130_fd_sc_hd__or2_1
X_16635_ _16635_/A _16697_/D _16635_/C _16635_/D vssd1 vssd1 vccd1 vccd1 _16636_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13847_ _13813_/X _26103_/Q _26004_/Q _15485_/S _16015_/A vssd1 vssd1 vccd1 vccd1
+ _13847_/X sky130_fd_sc_hd__a221o_1
XINSDIODE2_313 _19620_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_324 _19616_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_335 _19609_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_346 _19617_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_357 _19612_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19354_ _19385_/B _19354_/B vssd1 vssd1 vccd1 vccd1 _19354_/Y sky130_fd_sc_hd__nor2_1
X_16566_ _16566_/A vssd1 vssd1 vccd1 vccd1 _16575_/B sky130_fd_sc_hd__clkinv_2
XFILLER_250_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13778_ _14816_/A _13761_/X _13765_/X _13777_/X vssd1 vssd1 vccd1 vccd1 _13778_/X
+ sky130_fd_sc_hd__a31o_1
XINSDIODE2_368 _20487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_379 _16998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15517_ _15852_/A _15514_/X _15516_/X _13241_/A vssd1 vssd1 vccd1 vccd1 _15521_/A
+ sky130_fd_sc_hd__o211a_1
X_18305_ _18910_/A _18303_/X _18998_/A vssd1 vssd1 vccd1 vccd1 _18306_/C sky130_fd_sc_hd__o21a_1
X_12729_ _25581_/Q vssd1 vssd1 vccd1 vccd1 _14384_/A sky130_fd_sc_hd__clkinv_2
X_19285_ _18976_/X _19280_/X _19284_/X _19003_/X vssd1 vssd1 vccd1 vccd1 _19285_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_203_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16497_ _26359_/Q _26619_/Q _16500_/S vssd1 vssd1 vccd1 vccd1 _16497_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18236_ _27072_/Q _19058_/A _19059_/A _27170_/Q _19060_/A vssd1 vssd1 vccd1 vccd1
+ _18236_/X sky130_fd_sc_hd__a221o_1
X_15448_ _15446_/X _15447_/X _15473_/S vssd1 vssd1 vccd1 vccd1 _15448_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18167_ _27165_/Q _18121_/A _18121_/B _18166_/X vssd1 vssd1 vccd1 vccd1 _18167_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_8_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15379_ _26672_/Q _16240_/S _15378_/X _15169_/X vssd1 vssd1 vccd1 vccd1 _15379_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17118_ _20978_/A vssd1 vssd1 vccd1 vccd1 _24630_/A sky130_fd_sc_hd__buf_8
X_18098_ _18438_/A vssd1 vssd1 vccd1 vccd1 _18556_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_183_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17049_ _17042_/X _16986_/B _17039_/X input239/X vssd1 vssd1 vccd1 vccd1 _17049_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_143_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20060_ _20084_/A _20084_/B vssd1 vssd1 vccd1 vccd1 _20082_/B sky130_fd_sc_hd__xnor2_2
XFILLER_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_17 _18916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_28 _19207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_39 _19441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23750_ _23750_/A vssd1 vssd1 vccd1 vccd1 _23750_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20962_ _25857_/Q _20961_/X _20965_/S vssd1 vssd1 vccd1 vccd1 _20963_/A sky130_fd_sc_hd__mux2_1
XFILLER_260_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22701_ _23744_/A vssd1 vssd1 vccd1 vccd1 _22701_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23681_ _23681_/A vssd1 vssd1 vccd1 vccd1 _26746_/D sky130_fd_sc_hd__clkbuf_1
X_20893_ _20893_/A vssd1 vssd1 vccd1 vccd1 _25835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25420_ _23722_/X _27306_/Q _25426_/S vssd1 vssd1 vccd1 vccd1 _25421_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22632_ _22638_/A _22632_/B _22632_/C vssd1 vssd1 vccd1 vccd1 _22632_/X sky130_fd_sc_hd__or3_1
XFILLER_242_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25351_ _25351_/A vssd1 vssd1 vccd1 vccd1 _27275_/D sky130_fd_sc_hd__clkbuf_1
X_22563_ _26301_/Q _22565_/B vssd1 vssd1 vccd1 vccd1 _22563_/Y sky130_fd_sc_hd__nand2_1
XFILLER_139_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24302_ _24327_/A _24302_/B _24303_/B vssd1 vssd1 vccd1 vccd1 _26991_/D sky130_fd_sc_hd__nor3_1
XFILLER_210_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21514_ _20677_/A _21481_/X _21459_/X _21513_/X vssd1 vssd1 vccd1 vccd1 _21514_/X
+ sky130_fd_sc_hd__o211a_1
X_25282_ _23731_/X _27245_/Q _25282_/S vssd1 vssd1 vccd1 vccd1 _25283_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22494_ _22494_/A _22502_/B vssd1 vssd1 vccd1 vccd1 _22495_/A sky130_fd_sc_hd__and2_1
X_27021_ _27058_/CLK _27021_/D vssd1 vssd1 vccd1 vccd1 _27021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24233_ _26968_/Q _26967_/Q _24233_/C vssd1 vssd1 vccd1 vccd1 _24240_/C sky130_fd_sc_hd__and3_1
X_21445_ _21430_/X _18923_/X _21431_/X _25812_/Q _21403_/X vssd1 vssd1 vccd1 vccd1
+ _21445_/X sky130_fd_sc_hd__a221o_1
XFILLER_175_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24164_ _24164_/A _24169_/C vssd1 vssd1 vccd1 vccd1 _24164_/Y sky130_fd_sc_hd__nor2_1
XFILLER_207_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21376_ _21370_/Y _21375_/X _21359_/X vssd1 vssd1 vccd1 vccd1 _21376_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23115_ _26512_/Q _23114_/X _23115_/S vssd1 vssd1 vccd1 vccd1 _23116_/A sky130_fd_sc_hd__mux2_1
X_20327_ _20470_/A _20353_/A _20313_/A vssd1 vssd1 vccd1 vccd1 _20332_/A sky130_fd_sc_hd__a21o_1
X_24095_ _24095_/A vssd1 vssd1 vccd1 vccd1 _26915_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_268_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23046_ _23046_/A vssd1 vssd1 vccd1 vccd1 _26490_/D sky130_fd_sc_hd__clkbuf_1
X_20258_ _20470_/A _20259_/B vssd1 vssd1 vccd1 vccd1 _20261_/A sky130_fd_sc_hd__nor2_1
XTAP_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20189_ _20189_/A _20189_/B vssd1 vssd1 vccd1 vccd1 _20190_/A sky130_fd_sc_hd__and2_1
XFILLER_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26805_ _27288_/CLK _26805_/D vssd1 vssd1 vccd1 vccd1 _26805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_276_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24997_ _24341_/A _24900_/C _24776_/C _24777_/A vssd1 vssd1 vccd1 vccd1 _25124_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_57_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26736_ _27315_/CLK _26736_/D vssd1 vssd1 vccd1 vccd1 _26736_/Q sky130_fd_sc_hd__dfxtp_1
X_14750_ _14813_/S vssd1 vssd1 vccd1 vccd1 _14767_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_218_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23948_ _26850_/Q _23530_/X _23954_/S vssd1 vssd1 vccd1 vccd1 _23949_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _15063_/A _26104_/Q _26005_/Q _16050_/B _14713_/B vssd1 vssd1 vccd1 vccd1
+ _13701_/X sky130_fd_sc_hd__a221o_1
XFILLER_72_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26667_ _27249_/CLK _26667_/D vssd1 vssd1 vccd1 vccd1 _26667_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _14681_/A vssd1 vssd1 vccd1 vccd1 _14682_/A sky130_fd_sc_hd__clkbuf_4
X_23879_ _23879_/A vssd1 vssd1 vccd1 vccd1 _26819_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16420_ _26091_/Q _15221_/S _16419_/X _14753_/A vssd1 vssd1 vccd1 vccd1 _16420_/X
+ sky130_fd_sc_hd__o211a_1
X_13632_ _13608_/X _13615_/X _13620_/X _13631_/X _13168_/A vssd1 vssd1 vccd1 vccd1
+ _13632_/X sky130_fd_sc_hd__o311a_1
XFILLER_71_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25618_ _26940_/CLK _25618_/D vssd1 vssd1 vccd1 vccd1 _25618_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_189_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26598_ _27277_/CLK _26598_/D vssd1 vssd1 vccd1 vccd1 _26598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16351_ _25822_/Q _27256_/Q _16354_/S vssd1 vssd1 vccd1 vccd1 _16351_/X sky130_fd_sc_hd__mux2_1
X_25549_ _27000_/CLK _25549_/D vssd1 vssd1 vccd1 vccd1 _25549_/Q sky130_fd_sc_hd__dfxtp_1
X_13563_ _14237_/A _15708_/B _13562_/X _12944_/X vssd1 vssd1 vccd1 vccd1 _16292_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15302_ _26642_/Q _26738_/Q _15414_/A vssd1 vssd1 vccd1 vccd1 _15302_/X sky130_fd_sc_hd__mux2_1
X_19070_ _25552_/Q _18568_/X _19068_/X _19069_/X _18572_/X vssd1 vssd1 vccd1 vccd1
+ _19070_/X sky130_fd_sc_hd__a221o_1
XFILLER_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16282_ _16282_/A _16282_/B vssd1 vssd1 vccd1 vccd1 _20280_/A sky130_fd_sc_hd__nand2_8
XFILLER_201_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13494_ _14768_/A vssd1 vssd1 vccd1 vccd1 _13494_/X sky130_fd_sc_hd__buf_2
XFILLER_145_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18021_ _18721_/A _18976_/A _18019_/X _20624_/A vssd1 vssd1 vccd1 vccd1 _18021_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_157_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27219_ _27221_/CLK _27219_/D vssd1 vssd1 vccd1 vccd1 _27219_/Q sky130_fd_sc_hd__dfxtp_1
X_15233_ _14808_/A _15220_/X _15224_/X _15232_/X _16280_/S vssd1 vssd1 vccd1 vccd1
+ _15233_/X sky130_fd_sc_hd__a311o_1
XFILLER_200_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15164_ _14623_/A _15145_/X _15152_/X _15163_/X _14683_/A vssd1 vssd1 vccd1 vccd1
+ _15164_/X sky130_fd_sc_hd__a311o_1
XFILLER_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14115_ _14113_/X _14114_/X _14115_/S vssd1 vssd1 vccd1 vccd1 _14115_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19972_ _20194_/B _18781_/X _19911_/X _19971_/Y vssd1 vssd1 vccd1 vccd1 _19972_/X
+ sky130_fd_sc_hd__a31o_1
X_15095_ _15093_/X _15094_/X _15095_/S vssd1 vssd1 vccd1 vccd1 _15095_/X sky130_fd_sc_hd__mux2_1
XFILLER_268_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14046_ _26493_/Q _26365_/Q _14307_/S vssd1 vssd1 vccd1 vccd1 _14046_/X sky130_fd_sc_hd__mux2_1
X_18923_ _18555_/A _18913_/X _18922_/X vssd1 vssd1 vccd1 vccd1 _18923_/X sky130_fd_sc_hd__a21o_4
XFILLER_141_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18854_ _18855_/B _18855_/C _18855_/A vssd1 vssd1 vccd1 vccd1 _18905_/B sky130_fd_sc_hd__a21o_1
XFILLER_268_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17805_ _18317_/S _17805_/B vssd1 vssd1 vccd1 vccd1 _18325_/A sky130_fd_sc_hd__nor2_1
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15997_ _26664_/Q _25704_/Q _16013_/S vssd1 vssd1 vccd1 vccd1 _15997_/X sky130_fd_sc_hd__mux2_1
X_18785_ _18785_/A vssd1 vssd1 vccd1 vccd1 _19449_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_283_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17736_ _17736_/A _17736_/B _17736_/C _17736_/D vssd1 vssd1 vccd1 vccd1 _17747_/C
+ sky130_fd_sc_hd__or4_1
X_14948_ _14946_/X _14947_/X _14948_/S vssd1 vssd1 vccd1 vccd1 _14948_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_110 _21878_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14879_ _12775_/A _26713_/Q _26841_/Q _14846_/B _14688_/A vssd1 vssd1 vccd1 vccd1
+ _14879_/X sky130_fd_sc_hd__a221o_1
X_17667_ _18377_/A vssd1 vssd1 vccd1 vccd1 _19003_/A sky130_fd_sc_hd__buf_2
XFILLER_250_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_121 _23067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19406_ _25530_/Q _18746_/X _19403_/X _19405_/X _18770_/X vssd1 vssd1 vccd1 vccd1
+ _19406_/X sky130_fd_sc_hd__o221a_1
XFILLER_224_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_132 _12738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_143 _14228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16618_ _19011_/A _19034_/B vssd1 vssd1 vccd1 vccd1 _16637_/B sky130_fd_sc_hd__xnor2_4
XFILLER_250_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_154 _23542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17598_ _25918_/Q _17597_/X _13742_/Y _17518_/X vssd1 vssd1 vccd1 vccd1 _17598_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_165 _15808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_176 _16419_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19337_ _26968_/Q _18569_/X _18570_/X _27000_/Q vssd1 vssd1 vccd1 vccd1 _19337_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_250_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16549_ _16550_/A _17927_/A vssd1 vssd1 vccd1 vccd1 _17857_/A sky130_fd_sc_hd__and2_1
XINSDIODE2_187 _16830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_198 _19700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19268_ _19268_/A _19268_/B vssd1 vssd1 vccd1 vccd1 _19268_/Y sky130_fd_sc_hd__nor2_1
X_18219_ _18183_/X _18187_/X _18193_/Y _18218_/X vssd1 vssd1 vccd1 vccd1 _18219_/Y
+ sky130_fd_sc_hd__o22ai_4
X_19199_ _27092_/Q _19058_/X _19059_/X _27190_/Q _19060_/X vssd1 vssd1 vccd1 vccd1
+ _19199_/X sky130_fd_sc_hd__a221o_1
XFILLER_102_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21230_ _21552_/A _25862_/Q vssd1 vssd1 vccd1 vccd1 _21271_/A sky130_fd_sc_hd__nand2_2
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21161_ _21172_/A _21161_/B vssd1 vssd1 vccd1 vccd1 _21162_/A sky130_fd_sc_hd__or2_1
XFILLER_144_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20112_ _20276_/A vssd1 vssd1 vccd1 vccd1 _20112_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21092_ _21100_/A _21092_/B vssd1 vssd1 vccd1 vccd1 _21093_/A sky130_fd_sc_hd__or2_1
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24920_ _24920_/A _24923_/B vssd1 vssd1 vccd1 vccd1 _24920_/Y sky130_fd_sc_hd__nand2_1
X_20043_ _19796_/X _20042_/Y _20208_/A vssd1 vssd1 vccd1 vccd1 _20043_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24851_ _24847_/Y _24850_/X _24835_/X vssd1 vssd1 vccd1 vccd1 _27118_/D sky130_fd_sc_hd__a21oi_1
XFILLER_74_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23802_ _23702_/X _26785_/Q _23810_/S vssd1 vssd1 vccd1 vccd1 _23803_/A sky130_fd_sc_hd__mux2_1
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24782_ _24801_/A vssd1 vssd1 vccd1 vccd1 _24782_/X sky130_fd_sc_hd__buf_2
X_21994_ _26110_/Q _20916_/X _21994_/S vssd1 vssd1 vccd1 vccd1 _21995_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26521_ _27297_/CLK _26521_/D vssd1 vssd1 vccd1 vccd1 _26521_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23733_ _23733_/A vssd1 vssd1 vccd1 vccd1 _26762_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20945_ _23760_/A vssd1 vssd1 vccd1 vccd1 _20945_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26452_ _26453_/CLK _26452_/D vssd1 vssd1 vccd1 vccd1 _26452_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23664_ _23664_/A vssd1 vssd1 vccd1 vccd1 _26738_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20876_ _25830_/Q _20875_/X _20885_/S vssd1 vssd1 vccd1 vccd1 _20877_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25403_ _25403_/A vssd1 vssd1 vccd1 vccd1 _27298_/D sky130_fd_sc_hd__clkbuf_1
X_22615_ _22606_/X _22612_/Y _22614_/X vssd1 vssd1 vccd1 vccd1 _26320_/D sky130_fd_sc_hd__a21oi_1
XFILLER_186_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26383_ _27287_/CLK _26383_/D vssd1 vssd1 vccd1 vccd1 _26383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23595_ _26710_/Q _23594_/X _23604_/S vssd1 vssd1 vccd1 vccd1 _23596_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25334_ _25391_/S vssd1 vssd1 vccd1 vccd1 _25343_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22546_ _24277_/A vssd1 vssd1 vccd1 vccd1 _22600_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25265_ _23706_/X _27237_/Q _25271_/S vssd1 vssd1 vccd1 vccd1 _25266_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22477_ _22477_/A vssd1 vssd1 vccd1 vccd1 _26264_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27004_ _27004_/CLK _27004_/D vssd1 vssd1 vccd1 vccd1 _27004_/Q sky130_fd_sc_hd__dfxtp_1
X_24216_ _24216_/A _24221_/C vssd1 vssd1 vccd1 vccd1 _24216_/Y sky130_fd_sc_hd__nor2_1
XFILLER_154_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21428_ _21559_/B vssd1 vssd1 vccd1 vccd1 _21495_/B sky130_fd_sc_hd__clkbuf_1
X_25196_ _25225_/A vssd1 vssd1 vccd1 vccd1 _25196_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24147_ _24147_/A vssd1 vssd1 vccd1 vccd1 _26939_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_269_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21359_ _21556_/A vssd1 vssd1 vccd1 vccd1 _21359_/X sky130_fd_sc_hd__buf_4
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24078_ _24146_/S vssd1 vssd1 vccd1 vccd1 _24087_/S sky130_fd_sc_hd__buf_6
XFILLER_122_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15920_ _15606_/X _15918_/X _15919_/X _13545_/A vssd1 vssd1 vccd1 vccd1 _15921_/B
+ sky130_fd_sc_hd__a31o_1
X_23029_ _23029_/A vssd1 vssd1 vccd1 vccd1 _26485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_265_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15851_ _26534_/Q _26142_/Q _15857_/S vssd1 vssd1 vccd1 vccd1 _15852_/B sky130_fd_sc_hd__mux2_1
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _14802_/A vssd1 vssd1 vccd1 vccd1 _14803_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18570_ _18570_/A vssd1 vssd1 vccd1 vccd1 _18570_/X sky130_fd_sc_hd__clkbuf_2
X_15782_ _15770_/X _15773_/X _15781_/Y vssd1 vssd1 vccd1 vccd1 _15782_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_252_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ _20868_/A _13590_/A _13012_/A _22641_/B vssd1 vssd1 vccd1 vccd1 _12994_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14733_ _14733_/A vssd1 vssd1 vccd1 vccd1 _16524_/A sky130_fd_sc_hd__clkbuf_2
X_17521_ _22535_/B _17521_/B vssd1 vssd1 vccd1 vccd1 _25565_/D sky130_fd_sc_hd__nor2_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26719_ _26880_/CLK _26719_/D vssd1 vssd1 vccd1 vccd1 _26719_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17452_ _17458_/B vssd1 vssd1 vccd1 vccd1 _17453_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14664_ _16050_/B vssd1 vssd1 vccd1 vccd1 _16163_/S sky130_fd_sc_hd__buf_4
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ _12774_/A _26711_/Q _26839_/Q _16242_/S _15048_/X vssd1 vssd1 vccd1 vccd1
+ _16403_/X sky130_fd_sc_hd__a221o_1
X_13615_ _12745_/A _13609_/X _13612_/X _15819_/S vssd1 vssd1 vccd1 vccd1 _13615_/X
+ sky130_fd_sc_hd__o211a_1
X_17383_ _25546_/Q _17381_/B _17382_/Y vssd1 vssd1 vccd1 vccd1 _25546_/D sky130_fd_sc_hd__o21a_1
XFILLER_158_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14595_ _14595_/A vssd1 vssd1 vccd1 vccd1 _14596_/A sky130_fd_sc_hd__buf_2
XFILLER_158_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19122_ _19122_/A _19122_/B vssd1 vssd1 vccd1 vccd1 _19123_/B sky130_fd_sc_hd__nand2_1
XFILLER_41_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16334_ _25590_/Q _16284_/S _16333_/Y vssd1 vssd1 vccd1 vccd1 _17784_/A sky130_fd_sc_hd__o21ai_4
X_13546_ _13531_/X _13544_/X _14820_/A vssd1 vssd1 vccd1 vccd1 _13546_/X sky130_fd_sc_hd__o21a_1
XFILLER_201_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19053_ _18636_/X _19046_/Y _19049_/X _19052_/X vssd1 vssd1 vccd1 vccd1 _19053_/X
+ sky130_fd_sc_hd__a31o_1
X_16265_ _14801_/A _16261_/X _16264_/X _13314_/A vssd1 vssd1 vccd1 vccd1 _16265_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13477_ _13477_/A vssd1 vssd1 vccd1 vccd1 _13939_/A sky130_fd_sc_hd__buf_2
XFILLER_187_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15216_ _15201_/X _15208_/X _15212_/X _15215_/X _14759_/A _14779_/A vssd1 vssd1 vccd1
+ vccd1 _15217_/B sky130_fd_sc_hd__mux4_2
X_18004_ _17856_/X _17859_/X _18000_/X _18003_/X vssd1 vssd1 vccd1 vccd1 _18004_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_173_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16196_ _26509_/Q _26381_/Q _16260_/S vssd1 vssd1 vccd1 vccd1 _16196_/X sky130_fd_sc_hd__mux2_1
Xoutput306 _16736_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[10] sky130_fd_sc_hd__buf_2
Xoutput317 _16763_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[20] sky130_fd_sc_hd__buf_2
XFILLER_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput328 _16718_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[5] sky130_fd_sc_hd__buf_2
XFILLER_127_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15147_ _16061_/B vssd1 vssd1 vccd1 vccd1 _16073_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_236_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput339 _16881_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[14] sky130_fd_sc_hd__buf_2
XFILLER_236_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19955_ _27112_/Q _19691_/X _19905_/A vssd1 vssd1 vccd1 vccd1 _19955_/X sky130_fd_sc_hd__o21a_1
X_15078_ _16463_/A _23594_/A vssd1 vssd1 vccd1 vccd1 _15079_/C sky130_fd_sc_hd__nor2_1
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14029_ _25915_/Q _14029_/B vssd1 vssd1 vccd1 vccd1 _15874_/B sky130_fd_sc_hd__or2_1
X_18906_ _18906_/A _18906_/B vssd1 vssd1 vccd1 vccd1 _19582_/C sky130_fd_sc_hd__xor2_2
XFILLER_45_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19886_ _19920_/A _19883_/X _19885_/Y vssd1 vssd1 vccd1 vccd1 _19918_/A sky130_fd_sc_hd__o21ai_1
XFILLER_267_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18837_ _18775_/X _18835_/Y _18382_/A vssd1 vssd1 vccd1 vccd1 _18837_/X sky130_fd_sc_hd__o21ba_1
XFILLER_95_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18768_ _18830_/A vssd1 vssd1 vccd1 vccd1 _18768_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_209_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17719_ _17738_/A _21208_/B _17697_/Y vssd1 vssd1 vccd1 vccd1 _18161_/A sky130_fd_sc_hd__o21a_1
XFILLER_208_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18699_ _26952_/Q _18461_/X _18463_/X _26984_/Q vssd1 vssd1 vccd1 vccd1 _18699_/X
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_149_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27230_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20730_ _20787_/S vssd1 vssd1 vccd1 vccd1 _20739_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_251_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20661_ _20674_/A vssd1 vssd1 vccd1 vccd1 _20670_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_11_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22400_ _22400_/A _22400_/B vssd1 vssd1 vccd1 vccd1 _22400_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23380_ _26626_/Q _23057_/X _23386_/S vssd1 vssd1 vccd1 vccd1 _23381_/A sky130_fd_sc_hd__mux2_1
X_20592_ _23763_/A vssd1 vssd1 vccd1 vccd1 _20592_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22331_ _26223_/Q _22269_/A _22329_/X _22330_/X vssd1 vssd1 vccd1 vccd1 _26223_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25050_ _24674_/Y _25043_/X _25049_/Y _25027_/X vssd1 vssd1 vccd1 vccd1 _25050_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_118_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22262_ _26199_/Q _22249_/X _22255_/X _26300_/Q _22256_/X vssd1 vssd1 vccd1 vccd1
+ _22262_/X sky130_fd_sc_hd__a221o_1
XFILLER_118_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24001_ _24001_/A vssd1 vssd1 vccd1 vccd1 _26874_/D sky130_fd_sc_hd__clkbuf_1
X_21213_ _21866_/C _21211_/X _21562_/D vssd1 vssd1 vccd1 vccd1 _21244_/B sky130_fd_sc_hd__a21oi_1
XFILLER_151_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22193_ _26182_/Q _22185_/X _22192_/X _22181_/X vssd1 vssd1 vccd1 vccd1 _26182_/D
+ sky130_fd_sc_hd__o211a_1
X_21144_ _21144_/A vssd1 vssd1 vccd1 vccd1 _25920_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25952_ _25992_/CLK _25952_/D vssd1 vssd1 vccd1 vccd1 _25952_/Q sky130_fd_sc_hd__dfxtp_1
X_21075_ _21075_/A _21075_/B vssd1 vssd1 vccd1 vccd1 _21167_/A sky130_fd_sc_hd__or2_4
XFILLER_265_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24903_ _24941_/A vssd1 vssd1 vccd1 vccd1 _24954_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_20026_ _27146_/Q _20295_/B vssd1 vssd1 vccd1 vccd1 _20026_/X sky130_fd_sc_hd__and2_1
XFILLER_86_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25883_ _26599_/CLK _25883_/D vssd1 vssd1 vccd1 vccd1 _25883_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_247_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24834_ _20656_/A _24829_/X _24696_/Y _24830_/X vssd1 vssd1 vccd1 vccd1 _24834_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24765_ _24765_/A _24765_/B vssd1 vssd1 vccd1 vccd1 _25159_/A sky130_fd_sc_hd__nand2_4
XFILLER_61_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21977_ _26102_/Q _20891_/X _21983_/S vssd1 vssd1 vccd1 vccd1 _21978_/A sky130_fd_sc_hd__mux2_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26504_ _26604_/CLK _26504_/D vssd1 vssd1 vccd1 vccd1 _26504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23716_ _23715_/X _26757_/Q _23716_/S vssd1 vssd1 vccd1 vccd1 _23717_/A sky130_fd_sc_hd__mux2_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20928_ _20928_/A vssd1 vssd1 vccd1 vccd1 _25846_/D sky130_fd_sc_hd__clkbuf_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24696_ _24703_/A _24696_/B vssd1 vssd1 vccd1 vccd1 _24696_/Y sky130_fd_sc_hd__nand2_1
XFILLER_199_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26435_ _26467_/CLK _26435_/D vssd1 vssd1 vccd1 vccd1 _26435_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23647_ _23669_/A vssd1 vssd1 vccd1 vccd1 _23656_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_230_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20859_ _20859_/A vssd1 vssd1 vccd1 vccd1 _25825_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13400_ _25640_/Q _16130_/B _14401_/B _25608_/Q _12977_/A vssd1 vssd1 vccd1 vccd1
+ _13400_/X sky130_fd_sc_hd__a221o_1
XFILLER_168_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26366_ _26462_/CLK _26366_/D vssd1 vssd1 vccd1 vccd1 _26366_/Q sky130_fd_sc_hd__dfxtp_1
X_14380_ _26622_/Q _26718_/Q _14553_/S vssd1 vssd1 vccd1 vccd1 _14380_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23578_ _23578_/A vssd1 vssd1 vccd1 vccd1 _23578_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13331_ _27306_/Q _26563_/Q _16193_/S vssd1 vssd1 vccd1 vccd1 _13331_/X sky130_fd_sc_hd__mux2_1
X_25317_ _23782_/X _27261_/Q _25319_/S vssd1 vssd1 vccd1 vccd1 _25318_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22529_ _22529_/A vssd1 vssd1 vccd1 vccd1 _26288_/D sky130_fd_sc_hd__clkbuf_1
X_26297_ _26297_/CLK _26297_/D vssd1 vssd1 vccd1 vccd1 _26297_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16050_ _26927_/Q _16050_/B vssd1 vssd1 vccd1 vccd1 _16050_/X sky130_fd_sc_hd__or2_1
X_13262_ _13262_/A vssd1 vssd1 vccd1 vccd1 _15322_/A sky130_fd_sc_hd__clkbuf_4
X_25248_ _27230_/Q _25217_/A _25228_/X _24772_/B _25247_/X vssd1 vssd1 vccd1 vccd1
+ _27230_/D sky130_fd_sc_hd__o221a_1
XFILLER_183_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15001_ _14794_/X _14997_/X _15000_/X _17181_/A vssd1 vssd1 vccd1 vccd1 _15001_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13193_ _14047_/A vssd1 vssd1 vccd1 vccd1 _14458_/S sky130_fd_sc_hd__buf_2
XFILLER_151_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25179_ _25179_/A vssd1 vssd1 vccd1 vccd1 _25179_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19740_ _19833_/A vssd1 vssd1 vccd1 vccd1 _19740_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16952_ _16952_/A vssd1 vssd1 vccd1 vccd1 _16952_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_284_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15903_ _15901_/X _15902_/X _15903_/S vssd1 vssd1 vccd1 vccd1 _15903_/X sky130_fd_sc_hd__mux2_1
X_19671_ _19671_/A vssd1 vssd1 vccd1 vccd1 _20092_/B sky130_fd_sc_hd__clkbuf_4
X_16883_ _16906_/A _16883_/B vssd1 vssd1 vccd1 vccd1 _16883_/X sky130_fd_sc_hd__or2_1
XFILLER_65_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18622_ _18437_/A _18609_/X _18621_/X vssd1 vssd1 vccd1 vccd1 _18622_/X sky130_fd_sc_hd__a21o_4
XFILLER_37_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15834_ _26666_/Q _25706_/Q _15834_/S vssd1 vssd1 vccd1 vccd1 _15834_/X sky130_fd_sc_hd__mux2_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ _18542_/X _18544_/Y _18551_/Y _18552_/X vssd1 vssd1 vccd1 vccd1 _18553_/X
+ sky130_fd_sc_hd__o31a_1
X_15765_ _15761_/X _15764_/X _13313_/A vssd1 vssd1 vccd1 vccd1 _15765_/X sky130_fd_sc_hd__o21a_1
X_12977_ _12977_/A vssd1 vssd1 vccd1 vccd1 _14616_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _17504_/A _17504_/B _17504_/C vssd1 vssd1 vccd1 vccd1 _17662_/A sky130_fd_sc_hd__or3_4
X_14716_ _14593_/X _14620_/Y _14712_/Y _15079_/A vssd1 vssd1 vccd1 vccd1 _14716_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_206_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18484_ _19046_/B _19573_/A _18483_/X _18359_/X vssd1 vssd1 vccd1 vccd1 _18484_/X
+ sky130_fd_sc_hd__o211a_1
X_15696_ _15668_/Y _15679_/Y _15695_/Y _13314_/X _13466_/X vssd1 vssd1 vccd1 vccd1
+ _15696_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_75_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17435_ _24164_/A _17437_/B vssd1 vssd1 vccd1 vccd1 _17435_/Y sky130_fd_sc_hd__nor2_1
X_14647_ _14647_/A vssd1 vssd1 vccd1 vccd1 _15019_/A sky130_fd_sc_hd__buf_4
XFILLER_162_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17366_ _17414_/A vssd1 vssd1 vccd1 vccd1 _17366_/X sky130_fd_sc_hd__clkbuf_2
X_14578_ _16735_/A _16735_/B _18645_/S vssd1 vssd1 vccd1 vccd1 _14579_/B sky130_fd_sc_hd__a21oi_4
XFILLER_220_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19105_ _18371_/A _18686_/B _19105_/S vssd1 vssd1 vccd1 vccd1 _19105_/X sky130_fd_sc_hd__mux2_1
X_13529_ _13529_/A vssd1 vssd1 vccd1 vccd1 _14806_/A sky130_fd_sc_hd__buf_6
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16317_ _15165_/X _16315_/X _16316_/X vssd1 vssd1 vccd1 vccd1 _16317_/X sky130_fd_sc_hd__o21a_1
X_17297_ _17334_/A _17303_/C vssd1 vssd1 vccd1 vccd1 _17297_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16248_ _16230_/X _16247_/X _15071_/X vssd1 vssd1 vccd1 vccd1 _16248_/X sky130_fd_sc_hd__a21o_4
X_19036_ _18552_/X _19019_/Y _19035_/X _18779_/X vssd1 vssd1 vccd1 vccd1 _19036_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_161_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16179_ _13255_/A _26705_/Q _26833_/Q _15322_/A _15210_/A vssd1 vssd1 vccd1 vccd1
+ _16179_/X sky130_fd_sc_hd__a221o_1
XFILLER_102_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19938_ _22491_/A _19638_/X _19937_/X _19566_/X vssd1 vssd1 vccd1 vccd1 _25670_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19869_ _19864_/X _19865_/Y _19867_/Y _19868_/Y _19820_/S vssd1 vssd1 vccd1 vccd1
+ _19869_/X sky130_fd_sc_hd__a311o_1
XFILLER_110_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21900_ _20508_/X _26068_/Q _21900_/S vssd1 vssd1 vccd1 vccd1 _21901_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22880_ _26419_/Q _22730_/X _22884_/S vssd1 vssd1 vccd1 vccd1 _22881_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21831_ _21831_/A vssd1 vssd1 vccd1 vccd1 _26044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24550_ _24550_/A _24553_/B vssd1 vssd1 vccd1 vccd1 _24550_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21762_ _21762_/A vssd1 vssd1 vccd1 vccd1 _26014_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23501_ _23501_/A vssd1 vssd1 vccd1 vccd1 _26680_/D sky130_fd_sc_hd__clkbuf_1
X_20713_ _25466_/A vssd1 vssd1 vccd1 vccd1 _24770_/A sky130_fd_sc_hd__buf_8
X_24481_ _26313_/Q _24455_/X _24456_/X input227/X _24457_/X vssd1 vssd1 vccd1 vccd1
+ _24481_/X sky130_fd_sc_hd__a221o_1
X_21693_ _21693_/A vssd1 vssd1 vccd1 vccd1 _25985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26220_ _26222_/CLK _26220_/D vssd1 vssd1 vccd1 vccd1 _26220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23432_ _26650_/Q _23133_/X _23434_/S vssd1 vssd1 vccd1 vccd1 _23433_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20644_ _20644_/A vssd1 vssd1 vccd1 vccd1 _20644_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26151_ _27329_/A _26151_/D vssd1 vssd1 vccd1 vccd1 _26151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_258_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23363_ _23363_/A _23363_/B _25479_/Q vssd1 vssd1 vccd1 vccd1 _23860_/B sky130_fd_sc_hd__or3b_4
X_20575_ _23750_/A vssd1 vssd1 vccd1 vccd1 _20575_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_178_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25102_ _22509_/A _25092_/X _25087_/X _16637_/B _25079_/X vssd1 vssd1 vccd1 vccd1
+ _25102_/X sky130_fd_sc_hd__a221o_1
X_22314_ _26217_/Q _22299_/X _22313_/X _22304_/X vssd1 vssd1 vccd1 vccd1 _26217_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26082_ _27281_/CLK _26082_/D vssd1 vssd1 vccd1 vccd1 _26082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23294_ _20484_/X _26588_/Q _23302_/S vssd1 vssd1 vccd1 vccd1 _23295_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_46_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26823_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25033_ _25139_/A vssd1 vssd1 vccd1 vccd1 _25033_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22245_ _26193_/Q _22222_/X _22238_/X _26294_/Q _22241_/X vssd1 vssd1 vccd1 vccd1
+ _22245_/X sky130_fd_sc_hd__a221o_1
XFILLER_180_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22176_ _26176_/Q _22169_/X _22175_/X _22164_/X vssd1 vssd1 vccd1 vccd1 _26176_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_274_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21127_ _25916_/Q _21112_/X _21113_/X input15/X vssd1 vssd1 vccd1 vccd1 _21128_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_121_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26984_ _26987_/CLK _26984_/D vssd1 vssd1 vccd1 vccd1 _26984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_266_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21058_ _21058_/A vssd1 vssd1 vccd1 vccd1 _25897_/D sky130_fd_sc_hd__clkbuf_1
X_25935_ _26278_/CLK _25935_/D vssd1 vssd1 vccd1 vccd1 _25935_/Q sky130_fd_sc_hd__dfxtp_1
X_12900_ _13737_/A vssd1 vssd1 vccd1 vccd1 _12915_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20009_ _19824_/B _18845_/X _19663_/X _20008_/X vssd1 vssd1 vccd1 vccd1 _20009_/X
+ sky130_fd_sc_hd__o31a_1
X_13880_ _13878_/X _13879_/X _14010_/S vssd1 vssd1 vccd1 vccd1 _13880_/X sky130_fd_sc_hd__mux2_1
X_25866_ _26881_/CLK _25866_/D vssd1 vssd1 vccd1 vccd1 _25866_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12831_ _25598_/Q vssd1 vssd1 vccd1 vccd1 _12873_/A sky130_fd_sc_hd__inv_2
XFILLER_62_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24817_ _24814_/Y _24815_/X _24816_/X vssd1 vssd1 vccd1 vccd1 _27109_/D sky130_fd_sc_hd__a21oi_1
XFILLER_62_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25797_ _26297_/CLK _25797_/D vssd1 vssd1 vccd1 vccd1 _25797_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_62_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15550_ _26081_/Q _16078_/S _13723_/A _15549_/X vssd1 vssd1 vccd1 vccd1 _15550_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _19570_/A _19570_/B _12762_/C _12790_/C vssd1 vssd1 vccd1 vccd1 _12778_/B
+ sky130_fd_sc_hd__or4_4
X_24748_ _24764_/A _24748_/B vssd1 vssd1 vccd1 vccd1 _27093_/D sky130_fd_sc_hd__nor2_1
XFILLER_203_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14111_/X _14499_/X _14500_/X _13409_/A vssd1 vssd1 vccd1 vccd1 _14501_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _13011_/A _23568_/A _15480_/X _13028_/A vssd1 vssd1 vccd1 vccd1 _16901_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24679_ _24723_/A vssd1 vssd1 vccd1 vccd1 _24699_/A sky130_fd_sc_hd__clkbuf_2
X_12693_ _20249_/A _19916_/A _18138_/A vssd1 vssd1 vccd1 vccd1 _19570_/A sky130_fd_sc_hd__or3_2
XFILLER_230_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _13049_/A _14428_/X _14431_/X vssd1 vssd1 vccd1 vccd1 _14432_/X sky130_fd_sc_hd__a21o_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _25498_/Q _17131_/B _17219_/Y _17188_/X vssd1 vssd1 vccd1 vccd1 _25498_/D
+ sky130_fd_sc_hd__o211a_1
X_26418_ _26483_/CLK _26418_/D vssd1 vssd1 vccd1 vccd1 _26418_/Q sky130_fd_sc_hd__dfxtp_1
X_17151_ _17210_/A vssd1 vssd1 vccd1 vccd1 _17151_/X sky130_fd_sc_hd__buf_2
X_26349_ _26609_/CLK _26349_/D vssd1 vssd1 vccd1 vccd1 _26349_/Q sky130_fd_sc_hd__dfxtp_1
X_14363_ _14361_/X _14362_/Y _13179_/A vssd1 vssd1 vccd1 vccd1 _14562_/A sky130_fd_sc_hd__a21oi_2
Xinput16 core_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput27 core_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16102_ _26799_/Q _26443_/Q _16256_/B vssd1 vssd1 vccd1 vccd1 _16102_/X sky130_fd_sc_hd__mux2_1
X_13314_ _13314_/A vssd1 vssd1 vccd1 vccd1 _13314_/X sky130_fd_sc_hd__buf_6
Xinput38 core_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
X_17082_ _26232_/Q vssd1 vssd1 vccd1 vccd1 _17085_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_7_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput49 dout0[15] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14294_ _13664_/A _26879_/Q _26751_/Q _15775_/S _13943_/A vssd1 vssd1 vccd1 vccd1
+ _14294_/X sky130_fd_sc_hd__a221o_1
XFILLER_171_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16033_ _17828_/A _16035_/B vssd1 vssd1 vccd1 vccd1 _16633_/B sky130_fd_sc_hd__nor2_4
X_13245_ _14223_/S vssd1 vssd1 vccd1 vccd1 _13779_/A sky130_fd_sc_hd__buf_2
XFILLER_155_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13176_ _23546_/A _15073_/A _15388_/A _13175_/X vssd1 vssd1 vccd1 vccd1 _16860_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17984_ _18598_/S _18271_/B vssd1 vssd1 vccd1 vccd1 _17984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19723_ _24641_/A vssd1 vssd1 vccd1 vccd1 _24749_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16935_ _16986_/A _16935_/B vssd1 vssd1 vccd1 vccd1 _16936_/A sky130_fd_sc_hd__and2_1
XFILLER_238_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19654_ _19941_/A vssd1 vssd1 vccd1 vccd1 _20079_/A sky130_fd_sc_hd__buf_2
XFILLER_266_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16866_ _16895_/A vssd1 vssd1 vccd1 vccd1 _16893_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_237_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18605_ _13689_/A _17819_/B _18548_/A _18604_/X vssd1 vssd1 vccd1 vccd1 _18605_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_15817_ _12769_/A _26698_/Q _26826_/Q _13043_/A vssd1 vssd1 vccd1 vccd1 _15817_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19585_ _18597_/A _18078_/A _19585_/S vssd1 vssd1 vccd1 vccd1 _19585_/X sky130_fd_sc_hd__mux2_1
XFILLER_252_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16797_ _16932_/B vssd1 vssd1 vccd1 vccd1 _16952_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_280_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18536_ _18630_/A _18536_/B vssd1 vssd1 vccd1 vccd1 _18537_/A sky130_fd_sc_hd__and2_1
XFILLER_93_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15748_ _13010_/A _15750_/A _15747_/X _13027_/A _13756_/B vssd1 vssd1 vccd1 vccd1
+ _15748_/X sky130_fd_sc_hd__o2111a_2
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18467_ _25539_/Q _18459_/X _18464_/X _18154_/A _18466_/X vssd1 vssd1 vccd1 vccd1
+ _18467_/X sky130_fd_sc_hd__a221o_1
XFILLER_34_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15679_ _15673_/X _15678_/X _14817_/A vssd1 vssd1 vccd1 vccd1 _15679_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17418_ _17418_/A _25557_/Q _17418_/C vssd1 vssd1 vccd1 vccd1 _17420_/B sky130_fd_sc_hd__and3_1
XFILLER_194_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18398_ _27010_/Q _19063_/A _18397_/X _18565_/A vssd1 vssd1 vccd1 vccd1 _18398_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17349_ _17347_/X _17351_/C _17348_/Y vssd1 vssd1 vccd1 vccd1 _25535_/D sky130_fd_sc_hd__o21a_1
XFILLER_193_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20360_ _20352_/Y _20354_/X _20398_/A vssd1 vssd1 vccd1 vccd1 _20362_/A sky130_fd_sc_hd__o21ai_1
XFILLER_228_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19019_ _18792_/X _19013_/X _19018_/X vssd1 vssd1 vccd1 vccd1 _19019_/Y sky130_fd_sc_hd__o21ai_1
X_20291_ _27156_/Q _27090_/Q vssd1 vssd1 vccd1 vccd1 _20291_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22030_ _22030_/A vssd1 vssd1 vccd1 vccd1 _26126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23981_ _26865_/Q _23578_/X _23987_/S vssd1 vssd1 vccd1 vccd1 _23982_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_164_wb_clk_i clkbuf_opt_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26278_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25720_ _26904_/CLK _25720_/D vssd1 vssd1 vccd1 vccd1 _25720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22932_ _26442_/Q _22701_/X _22934_/S vssd1 vssd1 vccd1 vccd1 _22933_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25651_ _25661_/CLK _25651_/D vssd1 vssd1 vccd1 vccd1 _25651_/Q sky130_fd_sc_hd__dfxtp_1
X_22863_ _22863_/A vssd1 vssd1 vccd1 vccd1 _26411_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_249_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24602_ _24615_/A vssd1 vssd1 vccd1 vccd1 _24602_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21814_ _26037_/Q _20897_/X _21816_/S vssd1 vssd1 vccd1 vccd1 _21815_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25582_ _26684_/CLK _25582_/D vssd1 vssd1 vccd1 vccd1 _25582_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_58_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22794_ _26381_/Q _22711_/X _22800_/S vssd1 vssd1 vccd1 vccd1 _22795_/A sky130_fd_sc_hd__mux2_1
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27321_ _27321_/CLK _27321_/D vssd1 vssd1 vccd1 vccd1 _27321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_252_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24533_ _24538_/A _24627_/A vssd1 vssd1 vccd1 vccd1 _24533_/Y sky130_fd_sc_hd__nand2_1
XFILLER_169_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21745_ _21791_/S vssd1 vssd1 vccd1 vccd1 _21754_/S sky130_fd_sc_hd__buf_2
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27252_ _27252_/CLK _27252_/D vssd1 vssd1 vccd1 vccd1 _27252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24464_ _24464_/A hold3/A vssd1 vssd1 vccd1 vccd1 _24464_/Y sky130_fd_sc_hd__nand2_1
XFILLER_237_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21676_ _21698_/A vssd1 vssd1 vccd1 vccd1 _21685_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_212_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26203_ _26307_/CLK _26203_/D vssd1 vssd1 vccd1 vccd1 _26203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23415_ _26642_/Q _23108_/X _23419_/S vssd1 vssd1 vccd1 vccd1 _23416_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20627_ _26262_/Q _17190_/X _20626_/X _19965_/X vssd1 vssd1 vccd1 vccd1 _25725_/D
+ sky130_fd_sc_hd__o211a_1
X_27183_ _27188_/CLK _27183_/D vssd1 vssd1 vccd1 vccd1 _27183_/Q sky130_fd_sc_hd__dfxtp_2
X_24395_ _24457_/A vssd1 vssd1 vccd1 vccd1 _24395_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26134_ _26462_/CLK _26134_/D vssd1 vssd1 vccd1 vccd1 _26134_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_165_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23346_ _20592_/X _26612_/Q _23346_/S vssd1 vssd1 vccd1 vccd1 _23347_/A sky130_fd_sc_hd__mux2_1
X_20558_ _23562_/A vssd1 vssd1 vccd1 vccd1 _23738_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26065_ _26909_/CLK _26065_/D vssd1 vssd1 vccd1 vccd1 _26065_/Q sky130_fd_sc_hd__dfxtp_1
X_23277_ _26581_/Q _23130_/X _23277_/S vssd1 vssd1 vccd1 vccd1 _23278_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20489_ _20868_/B _21793_/B vssd1 vssd1 vccd1 vccd1 _25249_/C sky130_fd_sc_hd__nand2_4
XFILLER_180_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13030_ _15885_/A vssd1 vssd1 vccd1 vccd1 _13031_/A sky130_fd_sc_hd__clkbuf_4
X_25016_ _22474_/A _25015_/X _25004_/X _18151_/B _25005_/X vssd1 vssd1 vccd1 vccd1
+ _25016_/X sky130_fd_sc_hd__a221o_1
XFILLER_279_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22228_ _26191_/Q _22152_/A _22227_/X _22217_/X vssd1 vssd1 vccd1 vccd1 _26191_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22159_ _26171_/Q _22152_/X _22158_/X _22148_/X vssd1 vssd1 vccd1 vccd1 _26171_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_160_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26967_ _27000_/CLK _26967_/D vssd1 vssd1 vccd1 vccd1 _26967_/Q sky130_fd_sc_hd__dfxtp_1
X_14981_ _26808_/Q _26452_/Q _14981_/S vssd1 vssd1 vccd1 vccd1 _14981_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16720_ _17813_/B _16720_/B vssd1 vssd1 vccd1 vccd1 _18424_/A sky130_fd_sc_hd__xnor2_4
XFILLER_248_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13932_ _13915_/X _13930_/X _14602_/A vssd1 vssd1 vccd1 vccd1 _13932_/X sky130_fd_sc_hd__mux2_1
X_25918_ _27087_/CLK _25918_/D vssd1 vssd1 vccd1 vccd1 _25918_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_247_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26898_ _27285_/CLK _26898_/D vssd1 vssd1 vccd1 vccd1 _26898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_275_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13863_ _13863_/A vssd1 vssd1 vccd1 vccd1 _13863_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_219_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16651_ _25675_/Q _25674_/Q _25673_/Q _25672_/Q vssd1 vssd1 vccd1 vccd1 _16654_/B
+ sky130_fd_sc_hd__or4_1
X_25849_ _27283_/CLK _25849_/D vssd1 vssd1 vccd1 vccd1 _25849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_506 input253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15602_ _27312_/Q _26569_/Q _16110_/S vssd1 vssd1 vccd1 vccd1 _15602_/X sky130_fd_sc_hd__mux2_1
X_12814_ _13636_/B vssd1 vssd1 vccd1 vccd1 _15482_/A sky130_fd_sc_hd__dlymetal6s2s_1
XINSDIODE2_517 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19370_ _26969_/Q _18461_/A _18463_/A _27001_/Q vssd1 vssd1 vccd1 vccd1 _19370_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_222_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13794_ _16336_/A _13792_/X _13793_/X _14757_/A vssd1 vssd1 vccd1 vccd1 _13794_/X
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_528 _17007_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16582_ _17871_/A _17807_/A vssd1 vssd1 vccd1 vccd1 _16800_/B sky130_fd_sc_hd__nor2_2
XFILLER_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_539 _17019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18321_ _18321_/A _18321_/B vssd1 vssd1 vccd1 vccd1 _18321_/Y sky130_fd_sc_hd__nand2_1
X_12745_ _12745_/A vssd1 vssd1 vccd1 vccd1 _15559_/S sky130_fd_sc_hd__buf_2
X_15533_ _14599_/A _15531_/Y _15532_/X _14612_/A vssd1 vssd1 vccd1 vccd1 _15533_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15464_ _26926_/Q _15464_/B vssd1 vssd1 vccd1 vccd1 _15464_/X sky130_fd_sc_hd__or2_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ _18325_/B _18252_/B vssd1 vssd1 vccd1 vccd1 _19571_/D sky130_fd_sc_hd__nor2_1
XFILLER_176_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _20189_/A vssd1 vssd1 vccd1 vccd1 _20249_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_179_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14415_ _12673_/A _26489_/Q _26361_/Q _14173_/B _13022_/A vssd1 vssd1 vccd1 vccd1
+ _14415_/X sky130_fd_sc_hd__o221a_1
X_17203_ _25494_/Q _17151_/X _17146_/X _12721_/A vssd1 vssd1 vccd1 vccd1 _17204_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_169_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18183_ _18792_/A vssd1 vssd1 vccd1 vccd1 _18183_/X sky130_fd_sc_hd__buf_2
X_15395_ _14792_/A _15392_/X _15394_/X _15313_/X vssd1 vssd1 vccd1 vccd1 _15399_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14346_ _14342_/X _14343_/X _14344_/X _14345_/X _14431_/A _13121_/B vssd1 vssd1 vccd1
+ vccd1 _14346_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17134_ _22377_/A vssd1 vssd1 vccd1 vccd1 _17134_/X sky130_fd_sc_hd__buf_2
XFILLER_265_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17065_ _25973_/Q _17061_/X _16993_/X _17063_/X vssd1 vssd1 vccd1 vccd1 _17065_/X
+ sky130_fd_sc_hd__a22o_4
X_14277_ _14165_/A _14272_/X _14276_/X _12700_/A vssd1 vssd1 vccd1 vccd1 _14277_/X
+ sky130_fd_sc_hd__o211a_1
X_16016_ _13806_/X _16013_/X _16015_/X _13339_/A vssd1 vssd1 vccd1 vccd1 _16016_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13228_ _15662_/S vssd1 vssd1 vccd1 vccd1 _15422_/S sky130_fd_sc_hd__buf_4
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _13159_/A vssd1 vssd1 vccd1 vccd1 _15039_/A sky130_fd_sc_hd__buf_4
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _18799_/A vssd1 vssd1 vccd1 vccd1 _17967_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19706_ _19943_/B vssd1 vssd1 vccd1 vccd1 _19881_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16918_ _16907_/X _16968_/C _16917_/X vssd1 vssd1 vccd1 vccd1 _16919_/B sky130_fd_sc_hd__o21a_2
XFILLER_266_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17898_ _15528_/B _16038_/B _17933_/S vssd1 vssd1 vccd1 vccd1 _17898_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_19637_ _20052_/A vssd1 vssd1 vccd1 vccd1 _20225_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_265_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16849_ _16836_/X _16847_/Y _16946_/A _16842_/X vssd1 vssd1 vccd1 vccd1 _16850_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19568_ _25661_/Q _19568_/B vssd1 vssd1 vccd1 vccd1 _19568_/X sky130_fd_sc_hd__or2_1
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18519_ _18519_/A vssd1 vssd1 vccd1 vccd1 _18519_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_222_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19499_ _19512_/A vssd1 vssd1 vccd1 vccd1 _19499_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21530_ _21526_/Y _21529_/X _21492_/X vssd1 vssd1 vccd1 vccd1 _21530_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_22_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21461_ _21414_/X _21460_/X _21407_/X vssd1 vssd1 vccd1 vccd1 _21461_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_159_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23200_ _23200_/A vssd1 vssd1 vccd1 vccd1 _26546_/D sky130_fd_sc_hd__clkbuf_1
X_20412_ _27161_/Q _27095_/Q vssd1 vssd1 vccd1 vccd1 _20412_/Y sky130_fd_sc_hd__nand2_1
X_24180_ _26950_/Q _24176_/B _24179_/Y vssd1 vssd1 vccd1 vccd1 _26950_/D sky130_fd_sc_hd__o21a_1
X_21392_ _21390_/X _21391_/X _21367_/X vssd1 vssd1 vccd1 vccd1 _21392_/X sky130_fd_sc_hd__a21o_1
XFILLER_135_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23131_ _26517_/Q _23130_/X _23131_/S vssd1 vssd1 vccd1 vccd1 _23132_/A sky130_fd_sc_hd__mux2_1
X_20343_ _20343_/A _20343_/B vssd1 vssd1 vccd1 vccd1 _20343_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_108_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23062_ _23062_/A vssd1 vssd1 vccd1 vccd1 _26495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20274_ _19905_/X _20273_/X _20052_/X vssd1 vssd1 vccd1 vccd1 _20274_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_255_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22013_ _22013_/A vssd1 vssd1 vccd1 vccd1 _26118_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput206 localMemory_wb_adr_i[2] vssd1 vssd1 vccd1 vccd1 input206/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput217 localMemory_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input217/X sky130_fd_sc_hd__buf_6
X_26821_ _27301_/CLK _26821_/D vssd1 vssd1 vccd1 vccd1 _26821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_276_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput228 localMemory_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 input228/X sky130_fd_sc_hd__buf_6
XFILLER_248_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput239 localMemory_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 input239/X sky130_fd_sc_hd__buf_8
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26752_ _27301_/CLK _26752_/D vssd1 vssd1 vccd1 vccd1 _26752_/Q sky130_fd_sc_hd__dfxtp_1
X_23964_ _23964_/A vssd1 vssd1 vccd1 vccd1 _26857_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_271_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22915_ _26434_/Q _22675_/X _22923_/S vssd1 vssd1 vccd1 vccd1 _22916_/A sky130_fd_sc_hd__mux2_1
XFILLER_272_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25703_ _27277_/CLK _25703_/D vssd1 vssd1 vccd1 vccd1 _25703_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_244_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26683_ _26683_/CLK _26683_/D vssd1 vssd1 vccd1 vccd1 _26683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23895_ _23917_/A vssd1 vssd1 vccd1 vccd1 _23904_/S sky130_fd_sc_hd__buf_4
XFILLER_217_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22846_ _22846_/A vssd1 vssd1 vccd1 vccd1 _26403_/D sky130_fd_sc_hd__clkbuf_1
X_25634_ _26813_/CLK _25634_/D vssd1 vssd1 vccd1 vccd1 _25634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25565_ _25590_/CLK _25565_/D vssd1 vssd1 vccd1 vccd1 _25565_/Q sky130_fd_sc_hd__dfxtp_1
X_22777_ _22777_/A vssd1 vssd1 vccd1 vccd1 _26373_/D sky130_fd_sc_hd__clkbuf_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27304_ _27304_/CLK _27304_/D vssd1 vssd1 vccd1 vccd1 _27304_/Q sky130_fd_sc_hd__dfxtp_1
X_24516_ _24361_/S _25625_/Q _24515_/X vssd1 vssd1 vccd1 vccd1 _24758_/B sky130_fd_sc_hd__o21a_4
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21728_ _20500_/X _25999_/Q _21732_/S vssd1 vssd1 vccd1 vccd1 _21729_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25496_ _26940_/CLK _25496_/D vssd1 vssd1 vccd1 vccd1 _25496_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_61_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27275_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_235_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24447_ _27019_/Q _24421_/X _24446_/Y _24442_/X vssd1 vssd1 vccd1 vccd1 _27019_/D
+ sky130_fd_sc_hd__o211a_1
X_27235_ _27299_/CLK _27235_/D vssd1 vssd1 vccd1 vccd1 _27235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21659_ _21659_/A vssd1 vssd1 vccd1 vccd1 _25970_/D sky130_fd_sc_hd__clkbuf_1
X_14200_ _13834_/A _14198_/X _14199_/X _13939_/X vssd1 vssd1 vccd1 vccd1 _14204_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27166_ _27166_/CLK _27166_/D vssd1 vssd1 vccd1 vccd1 _27166_/Q sky130_fd_sc_hd__dfxtp_1
X_15180_ _26804_/Q _26448_/Q _16400_/S vssd1 vssd1 vccd1 vccd1 _15180_/X sky130_fd_sc_hd__mux2_1
X_24378_ _24408_/A _24915_/A vssd1 vssd1 vccd1 vccd1 _24378_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14131_ _14131_/A vssd1 vssd1 vccd1 vccd1 _14237_/B sky130_fd_sc_hd__buf_6
X_26117_ _27284_/CLK _26117_/D vssd1 vssd1 vccd1 vccd1 _26117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23329_ _20559_/X _26604_/Q _23335_/S vssd1 vssd1 vccd1 vccd1 _23330_/A sky130_fd_sc_hd__mux2_1
X_27097_ _27228_/CLK _27097_/D vssd1 vssd1 vccd1 vccd1 _27097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14062_ _14453_/A _25834_/Q _26034_/Q _13657_/A _14043_/A vssd1 vssd1 vccd1 vccd1
+ _14062_/X sky130_fd_sc_hd__a221o_1
XFILLER_165_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26048_ _26796_/CLK _26048_/D vssd1 vssd1 vccd1 vccd1 _26048_/Q sky130_fd_sc_hd__dfxtp_1
X_13013_ _13062_/A vssd1 vssd1 vccd1 vccd1 _14272_/S sky130_fd_sc_hd__clkbuf_4
X_18870_ _27147_/Q _19302_/B vssd1 vssd1 vccd1 vccd1 _18870_/X sky130_fd_sc_hd__or2_1
XFILLER_3_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17821_ _13552_/A _17821_/B vssd1 vssd1 vccd1 vccd1 _18676_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_17752_ _27199_/Q _18234_/A _18108_/B _17751_/X vssd1 vssd1 vccd1 vccd1 _17752_/X
+ sky130_fd_sc_hd__a22o_1
X_14964_ _27259_/Q _16501_/B vssd1 vssd1 vccd1 vccd1 _14964_/X sky130_fd_sc_hd__or2_1
XFILLER_236_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16703_ _20800_/B vssd1 vssd1 vccd1 vccd1 _16703_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13915_ _13911_/X _17556_/B _17556_/C _12916_/X _25908_/Q vssd1 vssd1 vccd1 vccd1
+ _13915_/X sky130_fd_sc_hd__o32a_1
XFILLER_207_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17683_ _17683_/A _17683_/B vssd1 vssd1 vccd1 vccd1 _17684_/B sky130_fd_sc_hd__nand2_1
XFILLER_47_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14895_ _15484_/S vssd1 vssd1 vccd1 vccd1 _16262_/S sky130_fd_sc_hd__buf_4
XFILLER_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19422_ _19477_/B _19422_/B vssd1 vssd1 vccd1 vccd1 _19422_/X sky130_fd_sc_hd__or2_2
XFILLER_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_303 _26368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16634_ _18726_/A _18726_/B vssd1 vssd1 vccd1 vccd1 _16635_/D sky130_fd_sc_hd__xnor2_4
XFILLER_35_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13846_ _13813_/X _25836_/Q _26036_/Q _15485_/S _15776_/A vssd1 vssd1 vccd1 vccd1
+ _13846_/X sky130_fd_sc_hd__a221o_1
XFILLER_207_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_314 _19620_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_325 _19616_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_336 _19609_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_347 _19617_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19353_ _25625_/Q _19153_/X _19351_/X _19352_/X vssd1 vssd1 vccd1 vccd1 _25625_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_204_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13777_ _13359_/X _13768_/X _13776_/X _13530_/X vssd1 vssd1 vccd1 vccd1 _13777_/X
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_358 _19612_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16565_ _16565_/A _19327_/A vssd1 vssd1 vccd1 vccd1 _16566_/A sky130_fd_sc_hd__xor2_4
XINSDIODE2_369 _20487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18304_ _18741_/A _18302_/X _18303_/X vssd1 vssd1 vccd1 vccd1 _18306_/B sky130_fd_sc_hd__a21oi_1
XFILLER_204_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15516_ _15516_/A _15516_/B vssd1 vssd1 vccd1 vccd1 _15516_/X sky130_fd_sc_hd__or2_1
X_12728_ _25582_/Q vssd1 vssd1 vccd1 vccd1 _14076_/A sky130_fd_sc_hd__clkinv_2
X_19284_ _19346_/C _19284_/B vssd1 vssd1 vccd1 vccd1 _19284_/X sky130_fd_sc_hd__or2_2
XFILLER_188_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16496_ _16480_/S _16493_/X _16495_/X _14662_/X vssd1 vssd1 vccd1 vccd1 _16496_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_176_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18235_ _27202_/Q _18813_/A vssd1 vssd1 vccd1 vccd1 _18235_/X sky130_fd_sc_hd__and2_1
X_15447_ _26798_/Q _26442_/Q _15471_/S vssd1 vssd1 vccd1 vccd1 _15447_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18166_ _18163_/X _18164_/X _18165_/X _18821_/A _18120_/D vssd1 vssd1 vccd1 vccd1
+ _18166_/X sky130_fd_sc_hd__a221o_1
X_15378_ _25712_/Q _16154_/B vssd1 vssd1 vccd1 vccd1 _15378_/X sky130_fd_sc_hd__or2_1
XFILLER_190_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17117_ _17658_/A _25566_/Q _20646_/A vssd1 vssd1 vccd1 vccd1 _17117_/X sky130_fd_sc_hd__a21o_1
X_14329_ _12767_/A _25760_/Q _14332_/S _26846_/Q _14331_/A vssd1 vssd1 vccd1 vccd1
+ _14330_/C sky130_fd_sc_hd__o221a_1
X_18097_ _18436_/A vssd1 vssd1 vccd1 vccd1 _18555_/A sky130_fd_sc_hd__buf_2
XFILLER_239_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17048_ _17001_/X _16980_/B _16980_/C _17039_/A input238/X vssd1 vssd1 vccd1 vccd1
+ _17048_/X sky130_fd_sc_hd__a32o_4
XFILLER_172_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18999_ _18947_/A _18996_/Y _18998_/X vssd1 vssd1 vccd1 vccd1 _18999_/X sky130_fd_sc_hd__o21a_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_18 _18951_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_29 _19254_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20961_ _23776_/A vssd1 vssd1 vccd1 vccd1 _20961_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22700_ _22700_/A vssd1 vssd1 vccd1 vccd1 _26345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23680_ _26746_/Q _23606_/X _23682_/S vssd1 vssd1 vccd1 vccd1 _23681_/A sky130_fd_sc_hd__mux2_1
X_20892_ _25835_/Q _20891_/X _20901_/S vssd1 vssd1 vccd1 vccd1 _20893_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22631_ _22631_/A _22631_/B vssd1 vssd1 vccd1 vccd1 _22632_/C sky130_fd_sc_hd__nand2_1
XFILLER_241_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25350_ _27275_/Q _23725_/A _25354_/S vssd1 vssd1 vccd1 vccd1 _25351_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22562_ _22553_/X _22560_/Y _22561_/X vssd1 vssd1 vccd1 vccd1 _26300_/D sky130_fd_sc_hd__a21oi_1
XFILLER_210_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24301_ _26991_/Q _26990_/Q _24301_/C vssd1 vssd1 vccd1 vccd1 _24303_/B sky130_fd_sc_hd__and3_1
XFILLER_194_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21513_ _21508_/X _21511_/X _21512_/X vssd1 vssd1 vccd1 vccd1 _21513_/X sky130_fd_sc_hd__a21o_1
X_25281_ _25281_/A vssd1 vssd1 vccd1 vccd1 _27244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22493_ _24630_/A vssd1 vssd1 vccd1 vccd1 _22502_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_222_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27020_ _27022_/CLK _27020_/D vssd1 vssd1 vccd1 vccd1 _27020_/Q sky130_fd_sc_hd__dfxtp_1
X_24232_ _26967_/Q _24233_/C _24231_/Y vssd1 vssd1 vccd1 vccd1 _26967_/D sky130_fd_sc_hd__o21a_1
X_21444_ _25483_/Q _21495_/B vssd1 vssd1 vccd1 vccd1 _21444_/X sky130_fd_sc_hd__or2_1
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24163_ _26945_/Q _24163_/B vssd1 vssd1 vccd1 vccd1 _24169_/C sky130_fd_sc_hd__and2_1
X_21375_ _21354_/X _21355_/X _21374_/Y _21259_/X vssd1 vssd1 vccd1 vccd1 _21375_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_174_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23114_ _23587_/A vssd1 vssd1 vccd1 vccd1 _23114_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20326_ _22522_/A _20225_/X _20318_/X _20325_/Y _20223_/X vssd1 vssd1 vccd1 vccd1
+ _25684_/D sky130_fd_sc_hd__o221a_1
X_24094_ _26915_/Q _23533_/X _24098_/S vssd1 vssd1 vccd1 vccd1 _24095_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23045_ _26490_/Q _23044_/X _23051_/S vssd1 vssd1 vccd1 vccd1 _23046_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20257_ _20448_/A vssd1 vssd1 vccd1 vccd1 _20470_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20188_ _22511_/A _20078_/X _20178_/X _20187_/X _20076_/X vssd1 vssd1 vccd1 vccd1
+ _25679_/D sky130_fd_sc_hd__o221a_1
XFILLER_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26804_ _26931_/CLK _26804_/D vssd1 vssd1 vccd1 vccd1 _26804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24996_ _24994_/X _24995_/X _20973_/A _24986_/Y vssd1 vssd1 vccd1 vccd1 _27166_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_264_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26735_ _27314_/CLK _26735_/D vssd1 vssd1 vccd1 vccd1 _26735_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23947_ _23947_/A vssd1 vssd1 vccd1 vccd1 _26849_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _26528_/Q _26136_/Q _16060_/S vssd1 vssd1 vccd1 vccd1 _13700_/X sky130_fd_sc_hd__mux2_1
XFILLER_245_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _14650_/X _14672_/X _14676_/X _14679_/X vssd1 vssd1 vccd1 vccd1 _14680_/X
+ sky130_fd_sc_hd__o211a_1
X_26666_ _27309_/CLK _26666_/D vssd1 vssd1 vccd1 vccd1 _26666_/Q sky130_fd_sc_hd__dfxtp_1
X_23878_ _23709_/X _26819_/Q _23882_/S vssd1 vssd1 vccd1 vccd1 _23879_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13631_ _15720_/S _13623_/X _13625_/X _13629_/X _13630_/X vssd1 vssd1 vccd1 vccd1
+ _13631_/X sky130_fd_sc_hd__a311o_1
X_22829_ _26396_/Q _22656_/X _22829_/S vssd1 vssd1 vccd1 vccd1 _22830_/A sky130_fd_sc_hd__mux2_1
XFILLER_260_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25617_ _26940_/CLK _25617_/D vssd1 vssd1 vccd1 vccd1 _25617_/Q sky130_fd_sc_hd__dfxtp_2
X_26597_ _27307_/CLK _26597_/D vssd1 vssd1 vccd1 vccd1 _26597_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_198_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13562_ _25927_/Q _13922_/B _13561_/Y _14404_/A vssd1 vssd1 vccd1 vccd1 _13562_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16350_ _16350_/A _16350_/B vssd1 vssd1 vccd1 vccd1 _16350_/X sky130_fd_sc_hd__or2_1
X_25548_ _25553_/CLK _25548_/D vssd1 vssd1 vccd1 vccd1 _25548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15301_ _15298_/X _15299_/X _15301_/S vssd1 vssd1 vccd1 vccd1 _15301_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16281_ _23584_/A _16280_/X _16281_/S vssd1 vssd1 vccd1 vccd1 _16282_/B sky130_fd_sc_hd__mux2_2
X_13493_ _13943_/A vssd1 vssd1 vccd1 vccd1 _14768_/A sky130_fd_sc_hd__buf_4
X_25479_ _26843_/CLK _25479_/D vssd1 vssd1 vccd1 vccd1 _25479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18020_ _25724_/Q vssd1 vssd1 vccd1 vccd1 _20624_/A sky130_fd_sc_hd__buf_4
X_27218_ _27227_/CLK _27218_/D vssd1 vssd1 vccd1 vccd1 _27218_/Q sky130_fd_sc_hd__dfxtp_1
X_15232_ _14803_/A _15227_/X _15231_/X _14818_/A vssd1 vssd1 vccd1 vccd1 _15232_/X
+ sky130_fd_sc_hd__o211a_1
X_15163_ _14649_/A _15157_/X _15162_/X _14679_/A vssd1 vssd1 vccd1 vccd1 _15163_/X
+ sky130_fd_sc_hd__o211a_1
X_27149_ _27227_/CLK _27149_/D vssd1 vssd1 vccd1 vccd1 _27149_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_154_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14114_ _26849_/Q _25763_/Q _14114_/S vssd1 vssd1 vccd1 vccd1 _14114_/X sky130_fd_sc_hd__mux2_1
X_19971_ _19971_/A _20227_/B vssd1 vssd1 vccd1 vccd1 _19971_/Y sky130_fd_sc_hd__nor2_1
X_15094_ _26934_/Q _26418_/Q _15121_/S vssd1 vssd1 vccd1 vccd1 _15094_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14045_ _13653_/S _14041_/X _14044_/X _13966_/A vssd1 vssd1 vccd1 vccd1 _14045_/X
+ sky130_fd_sc_hd__a211o_1
X_18922_ _25516_/Q _18559_/A _18919_/X _18921_/X _18574_/A vssd1 vssd1 vccd1 vccd1
+ _18922_/X sky130_fd_sc_hd__o221a_1
XFILLER_107_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18853_ _18794_/A _18794_/B _18838_/A vssd1 vssd1 vccd1 vccd1 _18855_/C sky130_fd_sc_hd__a21o_1
XFILLER_67_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17804_ _17798_/X _17803_/Y _18482_/A vssd1 vssd1 vccd1 vccd1 _18539_/C sky130_fd_sc_hd__a21oi_2
XFILLER_121_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18784_ _18967_/A _18784_/B vssd1 vssd1 vccd1 vccd1 _18784_/Y sky130_fd_sc_hd__nand2_2
XTAP_5770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15996_ _25577_/Q _16585_/A _15243_/A _15995_/X vssd1 vssd1 vccd1 vccd1 _17828_/A
+ sky130_fd_sc_hd__o22a_4
XTAP_5781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17735_ _17735_/A _17735_/B vssd1 vssd1 vccd1 vccd1 _17736_/D sky130_fd_sc_hd__nand2_1
X_14947_ _26124_/Q _26025_/Q _14970_/S vssd1 vssd1 vccd1 vccd1 _14947_/X sky130_fd_sc_hd__mux2_1
XFILLER_223_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17666_ _19589_/A vssd1 vssd1 vccd1 vccd1 _18377_/A sky130_fd_sc_hd__buf_2
XINSDIODE2_100 _21478_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14878_ _26649_/Q _26745_/Q _14878_/S vssd1 vssd1 vccd1 vccd1 _14878_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_111 _21878_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_122 _23520_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19405_ _25562_/Q _18763_/X _19404_/X _19069_/X _18768_/X vssd1 vssd1 vccd1 vccd1
+ _19405_/X sky130_fd_sc_hd__a221o_1
XFILLER_223_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_133 _12755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16617_ _19034_/A vssd1 vssd1 vccd1 vccd1 _19011_/A sky130_fd_sc_hd__inv_2
XINSDIODE2_144 _14077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13829_ _27302_/Q _26559_/Q _13829_/S vssd1 vssd1 vccd1 vccd1 _13829_/X sky130_fd_sc_hd__mux2_1
X_17597_ _17597_/A vssd1 vssd1 vccd1 vccd1 _17597_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_245_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_155 _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_166 _15805_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_177 _16419_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19336_ _27064_/Q _19055_/X _19333_/X _19335_/X _19066_/X vssd1 vssd1 vccd1 vccd1
+ _19336_/X sky130_fd_sc_hd__o221a_2
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16548_ _20703_/A _19472_/A _18059_/A vssd1 vssd1 vccd1 vccd1 _17927_/A sky130_fd_sc_hd__mux2_4
XINSDIODE2_188 _19769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_199 _19665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19267_ _18437_/X _19257_/X _19266_/X vssd1 vssd1 vccd1 vccd1 _19267_/X sky130_fd_sc_hd__a21o_4
XFILLER_149_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16479_ _16479_/A vssd1 vssd1 vccd1 vccd1 _16480_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_136_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18218_ _18269_/A _18212_/X _18216_/X _19018_/A vssd1 vssd1 vccd1 vccd1 _18218_/X
+ sky130_fd_sc_hd__a211o_1
X_19198_ _27222_/Q _19331_/B vssd1 vssd1 vccd1 vccd1 _19198_/X sky130_fd_sc_hd__and2_1
XFILLER_145_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18149_ _25726_/Q vssd1 vssd1 vccd1 vccd1 _19709_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_145_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21160_ _25925_/Q _21148_/X _21149_/X input25/X vssd1 vssd1 vccd1 vccd1 _21161_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20111_ _22505_/A _20078_/X _20103_/X _20110_/Y _20076_/X vssd1 vssd1 vccd1 vccd1
+ _25676_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21091_ _25906_/Q _21074_/X _21077_/X input36/X vssd1 vssd1 vccd1 vccd1 _21092_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20042_ _20082_/A _20042_/B vssd1 vssd1 vccd1 vccd1 _20042_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24850_ _20668_/A _24848_/X _24715_/Y _24849_/X vssd1 vssd1 vccd1 vccd1 _24850_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23801_ _23858_/S vssd1 vssd1 vccd1 vccd1 _23810_/S sky130_fd_sc_hd__buf_4
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24781_ _24781_/A _24781_/B vssd1 vssd1 vccd1 vccd1 _24781_/Y sky130_fd_sc_hd__nand2_1
X_21993_ _21993_/A vssd1 vssd1 vccd1 vccd1 _26109_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23732_ _23731_/X _26762_/Q _23732_/S vssd1 vssd1 vccd1 vccd1 _23733_/A sky130_fd_sc_hd__mux2_1
X_26520_ _26520_/CLK _26520_/D vssd1 vssd1 vccd1 vccd1 _26520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20944_ _20944_/A vssd1 vssd1 vccd1 vccd1 _25851_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26451_ _26903_/CLK _26451_/D vssd1 vssd1 vccd1 vccd1 _26451_/Q sky130_fd_sc_hd__dfxtp_1
X_23663_ _26738_/Q _23581_/X _23667_/S vssd1 vssd1 vccd1 vccd1 _23664_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20875_ _23690_/A vssd1 vssd1 vccd1 vccd1 _20875_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_198_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22614_ _24835_/A vssd1 vssd1 vccd1 vccd1 _22614_/X sky130_fd_sc_hd__clkbuf_2
X_25402_ _23696_/X _27298_/Q _25404_/S vssd1 vssd1 vccd1 vccd1 _25403_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26382_ _26610_/CLK _26382_/D vssd1 vssd1 vccd1 vccd1 _26382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23594_ _23594_/A vssd1 vssd1 vccd1 vccd1 _23594_/X sky130_fd_sc_hd__clkbuf_2
X_25333_ _25333_/A vssd1 vssd1 vccd1 vccd1 _27267_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22545_ _26295_/Q _22551_/B vssd1 vssd1 vccd1 vccd1 _22545_/Y sky130_fd_sc_hd__nand2_1
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25264_ _25264_/A vssd1 vssd1 vccd1 vccd1 _27236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22476_ _22476_/A _22480_/B vssd1 vssd1 vccd1 vccd1 _22477_/A sky130_fd_sc_hd__and2_1
X_24215_ _26962_/Q _24215_/B vssd1 vssd1 vccd1 vccd1 _24221_/C sky130_fd_sc_hd__and2_1
X_27003_ _27004_/CLK _27003_/D vssd1 vssd1 vccd1 vccd1 _27003_/Q sky130_fd_sc_hd__dfxtp_1
X_21427_ _25949_/Q _21378_/X _21426_/Y _21400_/X vssd1 vssd1 vccd1 vccd1 _25949_/D
+ sky130_fd_sc_hd__a211o_1
X_25195_ _24682_/B _25189_/X _25187_/X _27208_/Q _25191_/X vssd1 vssd1 vccd1 vccd1
+ _27208_/D sky130_fd_sc_hd__o221a_1
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24146_ _26939_/Q _23609_/X _24146_/S vssd1 vssd1 vccd1 vccd1 _24147_/A sky130_fd_sc_hd__mux2_1
X_21358_ _21354_/X _21355_/X _21357_/Y _21259_/X vssd1 vssd1 vccd1 vccd1 _21358_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_151_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20309_ _19246_/A _20355_/A _20308_/Y _20357_/A vssd1 vssd1 vccd1 vccd1 _20353_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_107_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24077_ _24133_/A vssd1 vssd1 vccd1 vccd1 _24146_/S sky130_fd_sc_hd__buf_4
XFILLER_268_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21289_ _21289_/A vssd1 vssd1 vccd1 vccd1 _21290_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23028_ _26485_/Q _22736_/X _23028_/S vssd1 vssd1 vccd1 vccd1 _23029_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ _26794_/Q _26438_/Q _15850_/S vssd1 vssd1 vccd1 vccd1 _15850_/X sky130_fd_sc_hd__mux2_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14802_/A sky130_fd_sc_hd__buf_2
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15781_ _15777_/X _15780_/X _13530_/X vssd1 vssd1 vccd1 vccd1 _15781_/Y sky130_fd_sc_hd__o21ai_1
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _17224_/A _25479_/Q vssd1 vssd1 vccd1 vccd1 _22641_/B sky130_fd_sc_hd__or2b_4
X_24979_ _27161_/Q _24923_/B _24978_/Y _24970_/X vssd1 vssd1 vccd1 vccd1 _27161_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17520_ _25565_/Q _20686_/A _17516_/X _17519_/X vssd1 vssd1 vccd1 vccd1 _17521_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26718_ _26878_/CLK _26718_/D vssd1 vssd1 vccd1 vccd1 _26718_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _15004_/S vssd1 vssd1 vccd1 vccd1 _14733_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _21868_/A _22536_/A vssd1 vssd1 vccd1 vccd1 _17458_/B sky130_fd_sc_hd__or2_1
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26649_ _26905_/CLK _26649_/D vssd1 vssd1 vccd1 vccd1 _26649_/Q sky130_fd_sc_hd__dfxtp_1
X_14663_ _16479_/A _14652_/X _14658_/X _14662_/X vssd1 vssd1 vccd1 vccd1 _14663_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _26647_/Q _26743_/Q _16402_/S vssd1 vssd1 vccd1 vccd1 _16402_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13614_ _13614_/A vssd1 vssd1 vccd1 vccd1 _15819_/S sky130_fd_sc_hd__buf_2
XFILLER_189_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17382_ _17382_/A _17389_/C vssd1 vssd1 vccd1 vccd1 _17382_/Y sky130_fd_sc_hd__nor2_1
X_14594_ _14594_/A vssd1 vssd1 vccd1 vccd1 _14595_/A sky130_fd_sc_hd__clkbuf_2
X_19121_ _19121_/A _19121_/B vssd1 vssd1 vccd1 vccd1 _19121_/Y sky130_fd_sc_hd__xnor2_4
X_16333_ _15290_/A _16332_/X _14718_/A vssd1 vssd1 vccd1 vccd1 _16333_/Y sky130_fd_sc_hd__o21ai_1
X_13545_ _13545_/A vssd1 vssd1 vccd1 vccd1 _14820_/A sky130_fd_sc_hd__buf_8
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19052_ _19358_/A _18732_/Y _19051_/X vssd1 vssd1 vccd1 vccd1 _19052_/X sky130_fd_sc_hd__o21a_1
X_13476_ _13472_/X _25839_/Q _26039_/Q _15496_/S _13762_/A vssd1 vssd1 vccd1 vccd1
+ _13476_/X sky130_fd_sc_hd__a221o_1
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16264_ _15313_/A _16262_/X _16263_/X _15417_/A vssd1 vssd1 vccd1 vccd1 _16264_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18003_ _18003_/A vssd1 vssd1 vccd1 vccd1 _18003_/X sky130_fd_sc_hd__buf_2
X_15215_ _15213_/X _15214_/X _16442_/S vssd1 vssd1 vccd1 vccd1 _15215_/X sky130_fd_sc_hd__mux2_1
XFILLER_275_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16195_ _16193_/X _16194_/X _16195_/S vssd1 vssd1 vccd1 vccd1 _16195_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput307 _16738_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[11] sky130_fd_sc_hd__buf_2
XFILLER_236_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15146_ _26868_/Q _25782_/Q _16387_/S vssd1 vssd1 vccd1 vccd1 _15146_/X sky130_fd_sc_hd__mux2_1
Xoutput318 _16765_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[21] sky130_fd_sc_hd__buf_2
Xoutput329 _16721_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[6] sky130_fd_sc_hd__buf_2
XFILLER_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15077_ _25624_/Q _14597_/X _15076_/X _14618_/X vssd1 vssd1 vccd1 vccd1 _23594_/A
+ sky130_fd_sc_hd__o22a_4
X_19954_ _20017_/C _19940_/Y _19941_/X _19953_/X vssd1 vssd1 vccd1 vccd1 _19954_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_206_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14028_ _13569_/A _14237_/C _15871_/B _14486_/A vssd1 vssd1 vccd1 vccd1 _14028_/X
+ sky130_fd_sc_hd__and4bb_1
X_18905_ _18905_/A _18905_/B vssd1 vssd1 vccd1 vccd1 _18906_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19885_ _19881_/A _19589_/B _20648_/A vssd1 vssd1 vccd1 vccd1 _19885_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_171_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18836_ _18608_/X _18834_/X _18835_/Y vssd1 vssd1 vccd1 vccd1 _18836_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_267_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18767_ _18829_/A vssd1 vssd1 vccd1 vccd1 _18767_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15979_ _15977_/X _15978_/X _15979_/S vssd1 vssd1 vccd1 vccd1 _15979_/X sky130_fd_sc_hd__mux2_1
XFILLER_255_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17718_ _17732_/A _17750_/A _17725_/D _19302_/B vssd1 vssd1 vccd1 vccd1 _18438_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_236_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18698_ _27048_/Q _18503_/X _18694_/X _18697_/X _18519_/X vssd1 vssd1 vccd1 vccd1
+ _18698_/X sky130_fd_sc_hd__o221a_1
XFILLER_224_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17649_ _19916_/A _17635_/X _17608_/A _17648_/Y vssd1 vssd1 vccd1 vccd1 _17650_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_224_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20660_ _20686_/A vssd1 vssd1 vccd1 vccd1 _20660_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_195_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_189_wb_clk_i _26681_/CLK vssd1 vssd1 vccd1 vccd1 _26483_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_220_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19319_ _12721_/A _19218_/X _19317_/Y _19318_/Y _19253_/X vssd1 vssd1 vccd1 vccd1
+ _19319_/X sky130_fd_sc_hd__a221o_2
XFILLER_220_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20591_ _23587_/A vssd1 vssd1 vccd1 vccd1 _23763_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_118_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27000_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_137_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22330_ _22428_/A vssd1 vssd1 vccd1 vccd1 _22330_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22261_ _26199_/Q _22254_/X _22260_/X _22258_/X vssd1 vssd1 vccd1 vccd1 _26199_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24000_ _26874_/Q _23606_/X _24002_/S vssd1 vssd1 vccd1 vccd1 _24001_/A sky130_fd_sc_hd__mux2_1
X_21212_ _21209_/B _21212_/B _24340_/S vssd1 vssd1 vccd1 vccd1 _21562_/D sky130_fd_sc_hd__and3b_1
XFILLER_133_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22192_ _26181_/Q _22186_/X _22179_/X input265/X _22187_/X vssd1 vssd1 vccd1 vccd1
+ _22192_/X sky130_fd_sc_hd__a221o_1
XFILLER_160_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21143_ _21154_/A _21143_/B vssd1 vssd1 vccd1 vccd1 _21144_/A sky130_fd_sc_hd__or2_1
XFILLER_160_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25951_ _25992_/CLK _25951_/D vssd1 vssd1 vccd1 vccd1 _25951_/Q sky130_fd_sc_hd__dfxtp_1
X_21074_ _21112_/A vssd1 vssd1 vccd1 vccd1 _21074_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24902_ _24902_/A vssd1 vssd1 vccd1 vccd1 _24902_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20025_ _20022_/Y _20023_/X _19999_/A _19999_/Y vssd1 vssd1 vccd1 vccd1 _20025_/X
+ sky130_fd_sc_hd__a211o_1
X_25882_ _26601_/CLK _25882_/D vssd1 vssd1 vccd1 vccd1 _25882_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24833_ _27114_/Q _24837_/B vssd1 vssd1 vccd1 vccd1 _24833_/Y sky130_fd_sc_hd__nand2_1
XFILLER_274_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21976_ _21976_/A vssd1 vssd1 vccd1 vccd1 _26101_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24764_ _24764_/A _24764_/B vssd1 vssd1 vccd1 vccd1 _27097_/D sky130_fd_sc_hd__nor2_1
XFILLER_132_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26503_ _27313_/CLK _26503_/D vssd1 vssd1 vccd1 vccd1 _26503_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23715_ _23715_/A vssd1 vssd1 vccd1 vccd1 _23715_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20927_ _25846_/Q _20926_/X _20933_/S vssd1 vssd1 vccd1 vccd1 _20928_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24695_ _24699_/A _24695_/B vssd1 vssd1 vccd1 vccd1 _27081_/D sky130_fd_sc_hd__nor2_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26434_ _26601_/CLK _26434_/D vssd1 vssd1 vccd1 vccd1 _26434_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23646_ _23646_/A vssd1 vssd1 vccd1 vccd1 _26730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20858_ _25825_/Q vssd1 vssd1 vccd1 vccd1 _20859_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_186_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26365_ _26462_/CLK _26365_/D vssd1 vssd1 vccd1 vccd1 _26365_/Q sky130_fd_sc_hd__dfxtp_2
X_23577_ _23577_/A vssd1 vssd1 vccd1 vccd1 _26704_/D sky130_fd_sc_hd__clkbuf_1
X_20789_ _22130_/A vssd1 vssd1 vccd1 vccd1 _22472_/B sky130_fd_sc_hd__clkbuf_4
X_13330_ _13330_/A vssd1 vssd1 vccd1 vccd1 _15333_/A sky130_fd_sc_hd__buf_4
XFILLER_195_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22528_ _22528_/A _22533_/B vssd1 vssd1 vccd1 vccd1 _22529_/A sky130_fd_sc_hd__and2_1
X_25316_ _25316_/A vssd1 vssd1 vccd1 vccd1 _27260_/D sky130_fd_sc_hd__clkbuf_1
X_26296_ _26327_/CLK _26296_/D vssd1 vssd1 vccd1 vccd1 _26296_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_183_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13261_ _13829_/S vssd1 vssd1 vccd1 vccd1 _13262_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22459_ _22459_/A vssd1 vssd1 vccd1 vccd1 _22459_/X sky130_fd_sc_hd__clkbuf_2
X_25247_ _27068_/Q _21873_/A input177/X _25214_/X _25178_/A vssd1 vssd1 vccd1 vccd1
+ _25247_/X sky130_fd_sc_hd__a41o_1
XFILLER_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15000_ _14755_/A _14998_/X _14999_/X _14804_/A vssd1 vssd1 vccd1 vccd1 _15000_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_68_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13192_ _13309_/A _14384_/A vssd1 vssd1 vccd1 vccd1 _14047_/A sky130_fd_sc_hd__nor2_2
XFILLER_157_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25178_ _25178_/A vssd1 vssd1 vccd1 vccd1 _25179_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24129_ _26931_/Q _23584_/X _24131_/S vssd1 vssd1 vccd1 vccd1 _24130_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16951_ _16951_/A vssd1 vssd1 vccd1 vccd1 _16980_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_111_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15902_ _27276_/Q _26469_/Q _15902_/S vssd1 vssd1 vccd1 vccd1 _15902_/X sky130_fd_sc_hd__mux2_1
X_19670_ _19670_/A vssd1 vssd1 vccd1 vccd1 _19671_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16882_ _16463_/X _23558_/A _15747_/X _16860_/B _15388_/X vssd1 vssd1 vccd1 vccd1
+ _16882_/X sky130_fd_sc_hd__o2111a_4
XFILLER_77_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18621_ _25510_/Q _18444_/A _18618_/X _18620_/X _18469_/A vssd1 vssd1 vccd1 vccd1
+ _18621_/X sky130_fd_sc_hd__o221a_1
XFILLER_253_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15833_ _15833_/A vssd1 vssd1 vccd1 vccd1 _23555_/A sky130_fd_sc_hd__buf_8
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ _18552_/A vssd1 vssd1 vccd1 vccd1 _18552_/X sky130_fd_sc_hd__clkbuf_2
X_15764_ _15205_/A _15762_/X _15763_/X _13304_/A vssd1 vssd1 vccd1 vccd1 _15764_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _14401_/A vssd1 vssd1 vccd1 vccd1 _12977_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ _18307_/A vssd1 vssd1 vccd1 vccd1 _17503_/X sky130_fd_sc_hd__buf_4
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14715_ _15830_/A vssd1 vssd1 vccd1 vccd1 _15079_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18483_ _18483_/A _19289_/B vssd1 vssd1 vccd1 vccd1 _18483_/X sky130_fd_sc_hd__or2_1
XFILLER_72_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15695_ _15683_/X _15686_/X _15694_/Y vssd1 vssd1 vccd1 vccd1 _15695_/Y sky130_fd_sc_hd__o21bai_2
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17434_ _25561_/Q _25562_/Q _17434_/C vssd1 vssd1 vccd1 vccd1 _17437_/B sky130_fd_sc_hd__and3_1
XFILLER_33_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14646_ _12777_/A _26422_/Q _16479_/A _14645_/X vssd1 vssd1 vccd1 vccd1 _14646_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17365_ _25541_/Q vssd1 vssd1 vccd1 vccd1 _17365_/X sky130_fd_sc_hd__buf_2
XFILLER_202_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14577_ _18593_/A _16732_/B _18604_/S vssd1 vssd1 vccd1 vccd1 _16735_/B sky130_fd_sc_hd__o21bai_4
X_19104_ _18683_/A _18683_/B _17988_/X _18269_/A vssd1 vssd1 vccd1 vccd1 _19104_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_202_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16316_ _15065_/A _26901_/Q _26773_/Q _16400_/S _15048_/A vssd1 vssd1 vccd1 vccd1
+ _16316_/X sky130_fd_sc_hd__a221o_1
XFILLER_119_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ _13241_/A _13518_/X _13526_/X _15836_/A vssd1 vssd1 vccd1 vccd1 _13528_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17296_ _25519_/Q _17296_/B vssd1 vssd1 vccd1 vccd1 _17303_/C sky130_fd_sc_hd__and2_1
XFILLER_174_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19035_ _18740_/X _19032_/Y _19033_/X _19042_/B _18839_/X vssd1 vssd1 vccd1 vccd1
+ _19035_/X sky130_fd_sc_hd__o32a_2
XFILLER_12_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16247_ _14623_/A _16234_/X _16238_/X _16246_/X _14683_/A vssd1 vssd1 vccd1 vccd1
+ _16247_/X sky130_fd_sc_hd__a311o_1
X_13459_ _14481_/B vssd1 vssd1 vccd1 vccd1 _14560_/S sky130_fd_sc_hd__buf_2
XFILLER_284_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16178_ _26641_/Q _26737_/Q _16178_/S vssd1 vssd1 vccd1 vccd1 _16178_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15129_ _20692_/A _19309_/A _16451_/S vssd1 vssd1 vccd1 vccd1 _17786_/A sky130_fd_sc_hd__mux2_2
XFILLER_142_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19937_ _19905_/X _19928_/X _19936_/X _19718_/X vssd1 vssd1 vccd1 vccd1 _19937_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19868_ _19864_/X _19865_/Y _19867_/Y vssd1 vssd1 vccd1 vccd1 _19868_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18819_ _27114_/Q _18812_/X _18814_/X _18818_/X vssd1 vssd1 vccd1 vccd1 _18819_/X
+ sky130_fd_sc_hd__o22a_2
X_19799_ _25730_/Q vssd1 vssd1 vccd1 vccd1 _20639_/A sky130_fd_sc_hd__buf_8
XFILLER_256_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21830_ _26044_/Q _20919_/X _21838_/S vssd1 vssd1 vccd1 vccd1 _21831_/A sky130_fd_sc_hd__mux2_1
XFILLER_283_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21761_ _20563_/X _26014_/Q _21765_/S vssd1 vssd1 vccd1 vccd1 _21762_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20712_ _20712_/A _20712_/B _20712_/C vssd1 vssd1 vccd1 vccd1 _20712_/X sky130_fd_sc_hd__or3_1
X_23500_ _26680_/Q _23127_/X _23502_/S vssd1 vssd1 vccd1 vccd1 _23501_/A sky130_fd_sc_hd__mux2_1
X_24480_ _24506_/A vssd1 vssd1 vccd1 vccd1 _24480_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21692_ _25985_/Q input197/X _21696_/S vssd1 vssd1 vccd1 vccd1 _21693_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23431_ _23431_/A vssd1 vssd1 vccd1 vccd1 _26649_/D sky130_fd_sc_hd__clkbuf_1
X_20643_ _20643_/A _20643_/B vssd1 vssd1 vccd1 vccd1 _20643_/X sky130_fd_sc_hd__or2_1
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26150_ _26611_/CLK _26150_/D vssd1 vssd1 vccd1 vccd1 _26150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23362_ _23362_/A vssd1 vssd1 vccd1 vccd1 _26619_/D sky130_fd_sc_hd__clkbuf_1
X_20574_ _23574_/A vssd1 vssd1 vccd1 vccd1 _23750_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22313_ _26216_/Q _22310_/X _22300_/X _26317_/Q _22301_/X vssd1 vssd1 vccd1 vccd1
+ _22313_/X sky130_fd_sc_hd__a221o_1
XFILLER_192_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25101_ _27184_/Q _25085_/X _25100_/X vssd1 vssd1 vccd1 vccd1 _27184_/D sky130_fd_sc_hd__o21ba_1
X_26081_ _27330_/A _26081_/D vssd1 vssd1 vccd1 vccd1 _26081_/Q sky130_fd_sc_hd__dfxtp_1
X_23293_ _23361_/S vssd1 vssd1 vccd1 vccd1 _23302_/S sky130_fd_sc_hd__buf_2
XFILLER_164_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25032_ _25114_/A vssd1 vssd1 vccd1 vccd1 _25139_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_22244_ _26193_/Q _22235_/X _22242_/X _22243_/X vssd1 vssd1 vccd1 vccd1 _26193_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22175_ _26175_/Q _22171_/X _22160_/X input274/X _22172_/X vssd1 vssd1 vccd1 vccd1
+ _22175_/X sky130_fd_sc_hd__a221o_1
XFILLER_219_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_86_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26684_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_278_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21126_ _21126_/A vssd1 vssd1 vccd1 vccd1 _25915_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_278_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26983_ _26987_/CLK _26983_/D vssd1 vssd1 vccd1 vccd1 _26983_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_15_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26604_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25934_ _26278_/CLK _25934_/D vssd1 vssd1 vccd1 vccd1 _25934_/Q sky130_fd_sc_hd__dfxtp_1
X_21057_ _25897_/Q _20961_/X _21059_/S vssd1 vssd1 vccd1 vccd1 _21058_/A sky130_fd_sc_hd__mux2_1
XFILLER_274_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20008_ _20008_/A _20055_/B vssd1 vssd1 vccd1 vccd1 _20008_/X sky130_fd_sc_hd__or2_1
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25865_ _25867_/CLK _25865_/D vssd1 vssd1 vccd1 vccd1 _25865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12830_ _25599_/Q vssd1 vssd1 vccd1 vccd1 _12862_/A sky130_fd_sc_hd__inv_2
X_24816_ _24835_/A vssd1 vssd1 vccd1 vccd1 _24816_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25796_ _25796_/CLK _25796_/D vssd1 vssd1 vccd1 vccd1 _25796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24747_ _27093_/Q _24744_/X _24746_/Y _24740_/X vssd1 vssd1 vccd1 vccd1 _24748_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_12761_ _25593_/Q _25592_/Q vssd1 vssd1 vccd1 vccd1 _12790_/C sky130_fd_sc_hd__or2_1
XFILLER_203_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21959_ _20621_/X _26095_/Q _21959_/S vssd1 vssd1 vccd1 vccd1 _21960_/A sky130_fd_sc_hd__mux2_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14500_ _12673_/A _27295_/Q _26552_/Q _14273_/B _13140_/A vssd1 vssd1 vccd1 vccd1
+ _14500_/X sky130_fd_sc_hd__o221a_1
XFILLER_215_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _15462_/X _15479_/X _14590_/A vssd1 vssd1 vccd1 vccd1 _15480_/X sky130_fd_sc_hd__a21o_4
XFILLER_15_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _17679_/A vssd1 vssd1 vccd1 vccd1 _18138_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_230_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24678_ _24678_/A _24678_/B vssd1 vssd1 vccd1 vccd1 _27077_/D sky130_fd_sc_hd__nor2_1
XFILLER_159_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14431_ _14431_/A _14431_/B _14431_/C vssd1 vssd1 vccd1 vccd1 _14431_/X sky130_fd_sc_hd__and3_1
XFILLER_30_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26417_ _26677_/CLK _26417_/D vssd1 vssd1 vccd1 vccd1 _26417_/Q sky130_fd_sc_hd__dfxtp_1
X_23629_ _23629_/A vssd1 vssd1 vccd1 vccd1 _26722_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17150_ _25478_/Q vssd1 vssd1 vccd1 vccd1 _22817_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26348_ _27283_/CLK _26348_/D vssd1 vssd1 vccd1 vccd1 _26348_/Q sky130_fd_sc_hd__dfxtp_1
X_14362_ _14362_/A _14362_/B vssd1 vssd1 vccd1 vccd1 _14362_/Y sky130_fd_sc_hd__nand2_1
Xinput17 core_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16101_ _16097_/X _16100_/X _14817_/A vssd1 vssd1 vccd1 vccd1 _16101_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_128_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput28 core_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_1
X_13313_ _13313_/A vssd1 vssd1 vccd1 vccd1 _13314_/A sky130_fd_sc_hd__buf_6
XFILLER_156_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput39 core_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17081_ _26233_/Q vssd1 vssd1 vccd1 vccd1 _17087_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14293_ _26655_/Q _25695_/Q _14296_/S vssd1 vssd1 vccd1 vccd1 _14293_/X sky130_fd_sc_hd__mux2_1
X_26279_ _26282_/CLK _26279_/D vssd1 vssd1 vccd1 vccd1 _26279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13244_ _13244_/A vssd1 vssd1 vccd1 vccd1 _14223_/S sky130_fd_sc_hd__buf_2
XFILLER_170_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16032_ _16632_/B vssd1 vssd1 vccd1 vccd1 _16035_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_171_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13175_ _13110_/X _13169_/X _14590_/A vssd1 vssd1 vccd1 vccd1 _13175_/X sky130_fd_sc_hd__a21o_2
XFILLER_124_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17983_ _17983_/A vssd1 vssd1 vccd1 vccd1 _18598_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19722_ _20079_/A vssd1 vssd1 vccd1 vccd1 _19722_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16934_ _16907_/X _16983_/C _16933_/X vssd1 vssd1 vccd1 vccd1 _16935_/B sky130_fd_sc_hd__o21a_2
XFILLER_77_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19653_ _20100_/A vssd1 vssd1 vccd1 vccd1 _19941_/A sky130_fd_sc_hd__clkbuf_1
X_16865_ _16865_/A vssd1 vssd1 vccd1 vccd1 _16865_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18604_ _18643_/A _18734_/A _18604_/S vssd1 vssd1 vccd1 vccd1 _18604_/X sky130_fd_sc_hd__mux2_1
X_15816_ _26634_/Q _26730_/Q _15816_/S vssd1 vssd1 vccd1 vccd1 _15816_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19584_ _18214_/A _18369_/A _19584_/S vssd1 vssd1 vccd1 vccd1 _19584_/X sky130_fd_sc_hd__mux2_1
XFILLER_281_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16796_ _21709_/B _17055_/D _16693_/X vssd1 vssd1 vccd1 vccd1 _16796_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_93_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18535_ _13852_/X _18285_/X _18534_/X _18409_/X _25605_/Q vssd1 vssd1 vccd1 vccd1
+ _18536_/B sky130_fd_sc_hd__a32o_1
XFILLER_280_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15747_ _15729_/X _15746_/X _13174_/A vssd1 vssd1 vccd1 vccd1 _15747_/X sky130_fd_sc_hd__a21o_4
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12959_ _12959_/A _25476_/Q vssd1 vssd1 vccd1 vccd1 _12996_/A sky130_fd_sc_hd__or2b_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18466_ _18466_/A vssd1 vssd1 vccd1 vccd1 _18466_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_233_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15678_ _16342_/S _15675_/X _15677_/X _13467_/A vssd1 vssd1 vccd1 vccd1 _15678_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17417_ _17418_/A _17418_/C _25557_/Q vssd1 vssd1 vccd1 vccd1 _17419_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14629_ _14952_/S vssd1 vssd1 vccd1 vccd1 _14700_/S sky130_fd_sc_hd__clkbuf_2
X_18397_ _19790_/A _18952_/B vssd1 vssd1 vccd1 vccd1 _18397_/X sky130_fd_sc_hd__or2_1
XFILLER_159_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17348_ _17347_/X _17351_/C _17318_/X vssd1 vssd1 vccd1 vccd1 _17348_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_158_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17279_ _17278_/X _17282_/C _17269_/X vssd1 vssd1 vccd1 vccd1 _17279_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_146_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19018_ _19018_/A _19018_/B _19018_/C _19018_/D vssd1 vssd1 vccd1 vccd1 _19018_/X
+ sky130_fd_sc_hd__or4_1
X_20290_ _27124_/Q _20248_/X _20276_/X _20289_/Y vssd1 vssd1 vccd1 vccd1 _20290_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_142_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23980_ _23980_/A vssd1 vssd1 vccd1 vccd1 _26864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_257_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22931_ _22931_/A vssd1 vssd1 vccd1 vccd1 _26441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25650_ _25660_/CLK _25650_/D vssd1 vssd1 vccd1 vccd1 _25650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22862_ _26411_/Q _22704_/X _22862_/S vssd1 vssd1 vccd1 vccd1 _22863_/A sky130_fd_sc_hd__mux2_1
XFILLER_283_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24601_ _27056_/Q _24589_/X _24600_/Y _24593_/X vssd1 vssd1 vccd1 vccd1 _27056_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21813_ _21813_/A vssd1 vssd1 vccd1 vccd1 _26036_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25581_ _25598_/CLK _25581_/D vssd1 vssd1 vccd1 vccd1 _25581_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_24_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22793_ _22793_/A vssd1 vssd1 vccd1 vccd1 _26380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_133_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27164_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_145_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27320_ _27324_/CLK _27320_/D vssd1 vssd1 vccd1 vccd1 _27320_/Q sky130_fd_sc_hd__dfxtp_1
X_21744_ _21744_/A vssd1 vssd1 vccd1 vccd1 _26006_/D sky130_fd_sc_hd__clkbuf_1
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24532_ _24768_/B vssd1 vssd1 vccd1 vccd1 _24627_/A sky130_fd_sc_hd__inv_2
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27251_ _27316_/CLK _27251_/D vssd1 vssd1 vccd1 vccd1 _27251_/Q sky130_fd_sc_hd__dfxtp_1
X_21675_ _21675_/A vssd1 vssd1 vccd1 vccd1 _25977_/D sky130_fd_sc_hd__clkbuf_1
X_24463_ _24454_/X _25615_/Q _24462_/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__o21ai_4
XFILLER_12_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26202_ _26307_/CLK _26202_/D vssd1 vssd1 vccd1 vccd1 _26202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20626_ _20626_/A _20630_/B vssd1 vssd1 vccd1 vccd1 _20626_/X sky130_fd_sc_hd__or2_1
X_23414_ _23414_/A vssd1 vssd1 vccd1 vccd1 _26641_/D sky130_fd_sc_hd__clkbuf_1
X_24394_ _24456_/A vssd1 vssd1 vccd1 vccd1 _24394_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27182_ _27188_/CLK _27182_/D vssd1 vssd1 vccd1 vccd1 _27182_/Q sky130_fd_sc_hd__dfxtp_1
X_26133_ _27266_/CLK _26133_/D vssd1 vssd1 vccd1 vccd1 _26133_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23345_ _23345_/A vssd1 vssd1 vccd1 vccd1 _26611_/D sky130_fd_sc_hd__clkbuf_1
X_20557_ _20557_/A vssd1 vssd1 vccd1 vccd1 _25707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_256_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26064_ _26909_/CLK _26064_/D vssd1 vssd1 vccd1 vccd1 _26064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23276_ _23276_/A vssd1 vssd1 vccd1 vccd1 _26580_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_285_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20488_ _20488_/A _21888_/C vssd1 vssd1 vccd1 vccd1 _21793_/B sky130_fd_sc_hd__nor2_4
XFILLER_98_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22227_ _26190_/Q _22222_/X _22206_/A _22226_/X _22155_/A vssd1 vssd1 vccd1 vccd1
+ _22227_/X sky130_fd_sc_hd__a221o_1
X_25015_ _25065_/A vssd1 vssd1 vccd1 vccd1 _25015_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22158_ _26170_/Q _22154_/X _22140_/X input254/X _22155_/X vssd1 vssd1 vccd1 vccd1
+ _22158_/X sky130_fd_sc_hd__a221o_1
XFILLER_152_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21109_ _25911_/Q _21094_/X _21095_/X input41/X vssd1 vssd1 vccd1 vccd1 _21110_/B
+ sky130_fd_sc_hd__o22a_1
X_26966_ _26995_/CLK _26966_/D vssd1 vssd1 vccd1 vccd1 _26966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14980_ _25752_/Q vssd1 vssd1 vccd1 vccd1 _20696_/A sky130_fd_sc_hd__clkinv_4
X_22089_ _22089_/A vssd1 vssd1 vccd1 vccd1 _26152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13931_ _14325_/S vssd1 vssd1 vccd1 vccd1 _14602_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25917_ _27188_/CLK _25917_/D vssd1 vssd1 vccd1 vccd1 _25917_/Q sky130_fd_sc_hd__dfxtp_4
X_26897_ _27252_/CLK _26897_/D vssd1 vssd1 vccd1 vccd1 _26897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16650_ _16639_/Y _16645_/X _16647_/X _16648_/X _24986_/A vssd1 vssd1 vccd1 vccd1
+ _17514_/A sky130_fd_sc_hd__o2111ai_4
X_13862_ _13862_/A vssd1 vssd1 vccd1 vccd1 _13863_/A sky130_fd_sc_hd__clkbuf_4
X_25848_ _26796_/CLK _25848_/D vssd1 vssd1 vccd1 vccd1 _25848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15601_ _16261_/S _15599_/X _15600_/X _13274_/A vssd1 vssd1 vccd1 vccd1 _15601_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_16_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_507 input269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12813_ _12813_/A vssd1 vssd1 vccd1 vccd1 _13636_/B sky130_fd_sc_hd__dlymetal6s2s_1
XINSDIODE2_518 _20990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16581_ _16581_/A _16581_/B vssd1 vssd1 vccd1 vccd1 _17871_/A sky130_fd_sc_hd__and2_1
XFILLER_262_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13793_ _15109_/A _26104_/Q _26005_/Q _15484_/S _13494_/X vssd1 vssd1 vccd1 vccd1
+ _13793_/X sky130_fd_sc_hd__a221o_1
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25779_ _27315_/CLK _25779_/D vssd1 vssd1 vccd1 vccd1 _25779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_529 _17048_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18320_ _18317_/X _18683_/B _18362_/A vssd1 vssd1 vccd1 vccd1 _18321_/B sky130_fd_sc_hd__mux2_1
X_15532_ _25647_/Q _15532_/B vssd1 vssd1 vccd1 vccd1 _15532_/X sky130_fd_sc_hd__and2_1
XFILLER_188_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12744_ _13884_/S vssd1 vssd1 vccd1 vccd1 _12745_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_187_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _18251_/A _18251_/B _18251_/C vssd1 vssd1 vccd1 vccd1 _18252_/B sky130_fd_sc_hd__and3_1
X_15463_ _27313_/Q _26570_/Q _15467_/S vssd1 vssd1 vccd1 vccd1 _15463_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _25596_/Q vssd1 vssd1 vccd1 vccd1 _20189_/A sky130_fd_sc_hd__buf_6
XFILLER_231_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17202_ _18338_/A vssd1 vssd1 vccd1 vccd1 _17222_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_230_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14414_ _14447_/A _14447_/B _13008_/A vssd1 vssd1 vccd1 vccd1 _16813_/B sky130_fd_sc_hd__a21o_4
XFILLER_187_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18182_ _18307_/A _18182_/B vssd1 vssd1 vccd1 vccd1 _18792_/A sky130_fd_sc_hd__or2_2
X_15394_ _15394_/A _15394_/B vssd1 vssd1 vccd1 vccd1 _15394_/X sky130_fd_sc_hd__or2_1
XFILLER_168_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17133_ _17133_/A _20689_/A vssd1 vssd1 vccd1 vccd1 _17133_/X sky130_fd_sc_hd__or2_1
XFILLER_129_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14345_ _13082_/A _26878_/Q _26750_/Q _13993_/A vssd1 vssd1 vccd1 vccd1 _14345_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17064_ _25972_/Q _17061_/X _16992_/X _17063_/X vssd1 vssd1 vccd1 vccd1 _17064_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_128_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14276_ _14273_/X _14274_/X _14275_/X _13889_/A _14089_/S vssd1 vssd1 vccd1 vccd1
+ _14276_/X sky130_fd_sc_hd__a221o_1
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16015_ _16015_/A _16015_/B vssd1 vssd1 vccd1 vccd1 _16015_/X sky130_fd_sc_hd__or2_1
X_13227_ _16110_/S vssd1 vssd1 vccd1 vccd1 _15662_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_171_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _26075_/Q _16067_/S _13723_/A _13157_/X vssd1 vssd1 vccd1 vccd1 _13158_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_285_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13089_ _15971_/S vssd1 vssd1 vccd1 vccd1 _13616_/S sky130_fd_sc_hd__clkbuf_4
X_17966_ _17966_/A vssd1 vssd1 vccd1 vccd1 _18799_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19705_ _19703_/X _19705_/B vssd1 vssd1 vccd1 vccd1 _19712_/A sky130_fd_sc_hd__and2b_1
X_16917_ _16909_/X _16868_/B _16867_/X _16910_/X _16911_/X vssd1 vssd1 vccd1 vccd1
+ _16917_/X sky130_fd_sc_hd__o221a_1
XFILLER_266_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17897_ _17880_/X _17894_/X _18416_/S vssd1 vssd1 vccd1 vccd1 _17897_/X sky130_fd_sc_hd__mux2_1
XFILLER_254_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19636_ _19636_/A _20712_/B vssd1 vssd1 vccd1 vccd1 _20052_/A sky130_fd_sc_hd__nand2_2
XFILLER_65_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16848_ _16906_/A _16848_/B vssd1 vssd1 vccd1 vccd1 _16946_/A sky130_fd_sc_hd__or2_1
XFILLER_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_253_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19567_ _19512_/A _19441_/X _19565_/X _19566_/X vssd1 vssd1 vccd1 vccd1 _25660_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_241_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16779_ _22526_/A _16769_/X _16770_/X _16575_/C vssd1 vssd1 vccd1 vccd1 _16779_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_80_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18518_ _27012_/Q _18514_/X _18517_/X _18455_/X vssd1 vssd1 vccd1 vccd1 _18518_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19498_ _19484_/X _18302_/X _19497_/X _19489_/X vssd1 vssd1 vccd1 vccd1 _25634_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18449_ _18756_/A vssd1 vssd1 vccd1 vccd1 _18449_/X sky130_fd_sc_hd__buf_2
XFILLER_61_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21460_ _20666_/A _21415_/X _21457_/X _21459_/X vssd1 vssd1 vccd1 vccd1 _21460_/X
+ sky130_fd_sc_hd__o211a_1
X_20411_ _27161_/Q _27095_/Q vssd1 vssd1 vccd1 vccd1 _20413_/A sky130_fd_sc_hd__nor2_1
X_21391_ _21364_/X _18702_/X _21365_/X _25808_/Q _21322_/X vssd1 vssd1 vccd1 vccd1
+ _21391_/X sky130_fd_sc_hd__a221o_1
XFILLER_190_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23130_ _23603_/A vssd1 vssd1 vccd1 vccd1 _23130_/X sky130_fd_sc_hd__clkbuf_2
X_20342_ _20342_/A _20342_/B vssd1 vssd1 vccd1 vccd1 _20343_/B sky130_fd_sc_hd__nand2_1
XFILLER_146_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23061_ _26495_/Q _23060_/X _23067_/S vssd1 vssd1 vccd1 vccd1 _23062_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20273_ _19993_/X _20270_/X _20271_/Y _20272_/Y vssd1 vssd1 vccd1 vccd1 _20273_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_103_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22012_ _26118_/Q _20942_/X _22016_/S vssd1 vssd1 vccd1 vccd1 _22013_/A sky130_fd_sc_hd__mux2_1
XFILLER_255_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput207 localMemory_wb_adr_i[3] vssd1 vssd1 vccd1 vccd1 input207/X sky130_fd_sc_hd__clkbuf_1
X_26820_ _26916_/CLK _26820_/D vssd1 vssd1 vccd1 vccd1 _26820_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput218 localMemory_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input218/X sky130_fd_sc_hd__buf_6
Xinput229 localMemory_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 input229/X sky130_fd_sc_hd__buf_8
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26751_ _26751_/CLK _26751_/D vssd1 vssd1 vccd1 vccd1 _26751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23963_ _26857_/Q _23552_/X _23965_/S vssd1 vssd1 vccd1 vccd1 _23964_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25702_ _26601_/CLK _25702_/D vssd1 vssd1 vccd1 vccd1 _25702_/Q sky130_fd_sc_hd__dfxtp_1
X_22914_ _22960_/S vssd1 vssd1 vccd1 vccd1 _22923_/S sky130_fd_sc_hd__buf_2
XFILLER_245_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26682_ _27259_/CLK _26682_/D vssd1 vssd1 vccd1 vccd1 _26682_/Q sky130_fd_sc_hd__dfxtp_1
X_23894_ _23894_/A vssd1 vssd1 vccd1 vccd1 _26826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25633_ _26813_/CLK _25633_/D vssd1 vssd1 vccd1 vccd1 _25633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22845_ _26403_/Q _22679_/X _22851_/S vssd1 vssd1 vccd1 vccd1 _22846_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25564_ _27004_/CLK _25564_/D vssd1 vssd1 vccd1 vccd1 _25564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22776_ _26373_/Q _22685_/X _22778_/S vssd1 vssd1 vccd1 vccd1 _22777_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27303_ _27303_/CLK _27303_/D vssd1 vssd1 vccd1 vccd1 _27303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24515_ _26320_/Q _21881_/X _21883_/X input234/X _24404_/X vssd1 vssd1 vccd1 vccd1
+ _24515_/X sky130_fd_sc_hd__a221o_2
XFILLER_52_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21727_ _21727_/A vssd1 vssd1 vccd1 vccd1 _25998_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25495_ _25796_/CLK _25495_/D vssd1 vssd1 vccd1 vccd1 _25495_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27234_ _27298_/CLK _27234_/D vssd1 vssd1 vccd1 vccd1 _27234_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24446_ _24464_/A _24944_/A vssd1 vssd1 vccd1 vccd1 _24446_/Y sky130_fd_sc_hd__nand2_1
XFILLER_197_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21658_ _25970_/Q input201/X _21662_/S vssd1 vssd1 vccd1 vccd1 _21659_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27165_ _27166_/CLK _27165_/D vssd1 vssd1 vccd1 vccd1 _27165_/Q sky130_fd_sc_hd__dfxtp_1
X_20609_ _23776_/A vssd1 vssd1 vccd1 vccd1 _20609_/X sky130_fd_sc_hd__clkbuf_2
X_24377_ _24472_/A _25601_/Q _24376_/X vssd1 vssd1 vccd1 vccd1 _24915_/A sky130_fd_sc_hd__o21ai_4
X_21589_ _21589_/A vssd1 vssd1 vccd1 vccd1 _21589_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26116_ _26610_/CLK _26116_/D vssd1 vssd1 vccd1 vccd1 _26116_/Q sky130_fd_sc_hd__dfxtp_1
X_14130_ _14443_/A vssd1 vssd1 vccd1 vccd1 _14187_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_23328_ _23328_/A vssd1 vssd1 vccd1 vccd1 _26603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27096_ _27228_/CLK _27096_/D vssd1 vssd1 vccd1 vccd1 _27096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_30_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26913_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14061_ _26785_/Q _26429_/Q _14474_/S vssd1 vssd1 vccd1 vccd1 _14061_/X sky130_fd_sc_hd__mux2_1
X_26047_ _26531_/CLK _26047_/D vssd1 vssd1 vccd1 vccd1 _26047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23259_ _23259_/A vssd1 vssd1 vccd1 vccd1 _26572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13012_ _13012_/A vssd1 vssd1 vccd1 vccd1 _14522_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_180_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17820_ _13691_/A _18593_/C _18634_/A vssd1 vssd1 vccd1 vccd1 _17820_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17751_ _27167_/Q _18615_/A vssd1 vssd1 vccd1 vccd1 _17751_/X sky130_fd_sc_hd__or2_1
X_26949_ _26987_/CLK _26949_/D vssd1 vssd1 vccd1 vccd1 _26949_/Q sky130_fd_sc_hd__dfxtp_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14963_ _26872_/Q _25786_/Q _14963_/S vssd1 vssd1 vccd1 vccd1 _14963_/X sky130_fd_sc_hd__mux2_1
XFILLER_282_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16702_ _25663_/Q vssd1 vssd1 vccd1 vccd1 _22476_/A sky130_fd_sc_hd__buf_2
XFILLER_236_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13914_ input167/X input138/X _14240_/S vssd1 vssd1 vccd1 vccd1 _17556_/C sky130_fd_sc_hd__mux2_8
X_17682_ _17691_/A _17682_/B vssd1 vssd1 vccd1 vccd1 _21214_/B sky130_fd_sc_hd__or2_1
XFILLER_75_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14894_ _14733_/A _14889_/X _14893_/X _14760_/A vssd1 vssd1 vccd1 vccd1 _14904_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_263_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19421_ _20701_/A _19421_/B vssd1 vssd1 vccd1 vccd1 _19422_/B sky130_fd_sc_hd__and2_1
X_16633_ _16633_/A _16633_/B vssd1 vssd1 vccd1 vccd1 _18726_/A sky130_fd_sc_hd__nor2_8
XFILLER_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13845_ _16004_/S vssd1 vssd1 vccd1 vccd1 _15485_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_62_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_304 _25696_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_315 _19620_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_326 _19616_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_337 _19609_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19352_ _19352_/A vssd1 vssd1 vccd1 vccd1 _19352_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16564_ _19325_/A _16567_/B _19294_/S vssd1 vssd1 vccd1 vccd1 _16565_/A sky130_fd_sc_hd__a21oi_2
X_13776_ _13762_/A _13769_/X _13772_/X _15486_/A vssd1 vssd1 vccd1 vccd1 _13776_/X
+ sky130_fd_sc_hd__a211o_1
XINSDIODE2_348 _19617_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_359 input215/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18303_ _19728_/A _17444_/D _18303_/S vssd1 vssd1 vccd1 vccd1 _18303_/X sky130_fd_sc_hd__mux2_1
X_15515_ _25815_/Q _27249_/Q _15515_/S vssd1 vssd1 vccd1 vccd1 _15516_/B sky130_fd_sc_hd__mux2_1
XFILLER_203_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19283_ _19283_/A _19283_/B vssd1 vssd1 vccd1 vccd1 _19284_/B sky130_fd_sc_hd__nor2_1
X_12727_ _25576_/Q vssd1 vssd1 vccd1 vccd1 _17669_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_149_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16495_ _25828_/Q _16493_/S _16499_/S _16494_/X vssd1 vssd1 vccd1 vccd1 _16495_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18234_ _18234_/A vssd1 vssd1 vccd1 vccd1 _18813_/A sky130_fd_sc_hd__clkbuf_2
X_15446_ _25847_/Q _26047_/Q _15459_/S vssd1 vssd1 vccd1 vccd1 _15446_/X sky130_fd_sc_hd__mux2_1
XFILLER_276_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18165_ _27135_/Q _27039_/Q _18615_/A vssd1 vssd1 vccd1 vccd1 _18165_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15377_ _15373_/X _15376_/X _16328_/A vssd1 vssd1 vccd1 vccd1 _15377_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17116_ _17635_/A vssd1 vssd1 vccd1 vccd1 _20646_/A sky130_fd_sc_hd__buf_6
X_14328_ _12767_/A _26394_/Q _14263_/S _26910_/Q _13139_/A vssd1 vssd1 vccd1 vccd1
+ _14330_/B sky130_fd_sc_hd__o221a_1
XFILLER_172_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18096_ _18554_/A vssd1 vssd1 vccd1 vccd1 _18435_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17047_ _17001_/X _16975_/B _16975_/C _17013_/X input236/X vssd1 vssd1 vccd1 vccd1
+ _17047_/X sky130_fd_sc_hd__a32o_4
X_14259_ _26067_/Q _15989_/S _14495_/A _14258_/X vssd1 vssd1 vccd1 vccd1 _14259_/X
+ sky130_fd_sc_hd__o211a_1
X_27328__488 vssd1 vssd1 vccd1 vccd1 _27328__488/HI localMemory_wb_error_o sky130_fd_sc_hd__conb_1
XFILLER_171_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18998_ _18998_/A vssd1 vssd1 vccd1 vccd1 _18998_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_19 _19035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17949_ _17818_/B _16287_/B _17949_/S vssd1 vssd1 vccd1 vccd1 _17949_/X sky130_fd_sc_hd__mux2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20960_ _20960_/A vssd1 vssd1 vccd1 vccd1 _25856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19619_ _27059_/Q _21264_/A input183/X _19616_/X _19618_/X vssd1 vssd1 vccd1 vccd1
+ _19628_/B sky130_fd_sc_hd__a311o_1
X_20891_ _23706_/A vssd1 vssd1 vccd1 vccd1 _20891_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_214_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22630_ _26325_/Q _22630_/B _22638_/D vssd1 vssd1 vccd1 vccd1 _22631_/B sky130_fd_sc_hd__or3b_1
XFILLER_198_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22561_ _22600_/A vssd1 vssd1 vccd1 vccd1 _22561_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_250_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24300_ _26990_/Q _24301_/C _26991_/Q vssd1 vssd1 vccd1 vccd1 _24302_/B sky130_fd_sc_hd__a21oi_1
X_21512_ _21589_/A vssd1 vssd1 vccd1 vccd1 _21512_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25280_ _23728_/X _27244_/Q _25282_/S vssd1 vssd1 vccd1 vccd1 _25281_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22492_ _22492_/A vssd1 vssd1 vccd1 vccd1 _26271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24231_ _24237_/A _24231_/B vssd1 vssd1 vccd1 vccd1 _24231_/Y sky130_fd_sc_hd__nor2_1
X_21443_ _21573_/A vssd1 vssd1 vccd1 vccd1 _21443_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_182_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24162_ _26944_/Q _24159_/A _24161_/Y vssd1 vssd1 vccd1 vccd1 _26944_/D sky130_fd_sc_hd__o21a_1
XFILLER_119_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21374_ _21374_/A vssd1 vssd1 vccd1 vccd1 _21374_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23113_ _23113_/A vssd1 vssd1 vccd1 vccd1 _26511_/D sky130_fd_sc_hd__clkbuf_1
X_20325_ _19905_/X _20324_/X _20052_/X vssd1 vssd1 vccd1 vccd1 _20325_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_190_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24093_ _24093_/A vssd1 vssd1 vccd1 vccd1 _26914_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23044_ _23517_/A vssd1 vssd1 vccd1 vccd1 _23044_/X sky130_fd_sc_hd__buf_2
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20256_ _20426_/A vssd1 vssd1 vccd1 vccd1 _20448_/A sky130_fd_sc_hd__clkbuf_1
XTAP_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20187_ _20179_/X _20185_/X _20186_/X vssd1 vssd1 vccd1 vccd1 _20187_/X sky130_fd_sc_hd__a21o_1
XTAP_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26803_ _27329_/A _26803_/D vssd1 vssd1 vccd1 vccd1 _26803_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24995_ _24994_/B _24671_/Y _19642_/X _24988_/X vssd1 vssd1 vccd1 vccd1 _24995_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26734_ _27308_/CLK _26734_/D vssd1 vssd1 vccd1 vccd1 _26734_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23946_ _26849_/Q _23526_/X _23954_/S vssd1 vssd1 vccd1 vccd1 _23947_/A sky130_fd_sc_hd__mux2_1
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26665_ _26827_/CLK _26665_/D vssd1 vssd1 vccd1 vccd1 _26665_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23877_ _23877_/A vssd1 vssd1 vccd1 vccd1 _26818_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13630_ _13630_/A vssd1 vssd1 vccd1 vccd1 _13630_/X sky130_fd_sc_hd__buf_2
X_25616_ _26940_/CLK _25616_/D vssd1 vssd1 vccd1 vccd1 _25616_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_71_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22828_ _22828_/A vssd1 vssd1 vccd1 vccd1 _26395_/D sky130_fd_sc_hd__clkbuf_1
X_26596_ _27276_/CLK _26596_/D vssd1 vssd1 vccd1 vccd1 _26596_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_204_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25547_ _25547_/CLK _25547_/D vssd1 vssd1 vccd1 vccd1 _25547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13561_ _13561_/A _13561_/B vssd1 vssd1 vccd1 vccd1 _13561_/Y sky130_fd_sc_hd__nor2_1
X_22759_ _26365_/Q _22659_/X _22767_/S vssd1 vssd1 vccd1 vccd1 _22760_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15300_ _15300_/A vssd1 vssd1 vccd1 vccd1 _15301_/S sky130_fd_sc_hd__buf_4
XFILLER_158_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16280_ _16266_/X _16279_/X _16280_/S vssd1 vssd1 vccd1 vccd1 _16280_/X sky130_fd_sc_hd__mux2_2
X_13492_ _15758_/S vssd1 vssd1 vccd1 vccd1 _13492_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_212_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25478_ _26843_/CLK _25478_/D vssd1 vssd1 vccd1 vccd1 _25478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27217_ _27221_/CLK _27217_/D vssd1 vssd1 vccd1 vccd1 _27217_/Q sky130_fd_sc_hd__dfxtp_1
X_15231_ _14753_/A _15228_/X _15230_/X _14792_/A vssd1 vssd1 vccd1 vccd1 _15231_/X
+ sky130_fd_sc_hd__a211o_1
X_24429_ _24434_/A _24936_/A vssd1 vssd1 vccd1 vccd1 _24429_/Y sky130_fd_sc_hd__nand2_1
XFILLER_139_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27148_ _27154_/CLK _27148_/D vssd1 vssd1 vccd1 vccd1 _27148_/Q sky130_fd_sc_hd__dfxtp_4
X_15162_ _16224_/S _15159_/X _15161_/X _14660_/A vssd1 vssd1 vccd1 vccd1 _15162_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14113_ _25802_/Q _27236_/Q _14114_/S vssd1 vssd1 vccd1 vccd1 _14113_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19970_ _25736_/Q vssd1 vssd1 vccd1 vccd1 _20654_/A sky130_fd_sc_hd__clkbuf_16
X_15093_ _27321_/Q _26578_/Q _15121_/S vssd1 vssd1 vccd1 vccd1 _15093_/X sky130_fd_sc_hd__mux2_1
X_27079_ _27198_/CLK _27079_/D vssd1 vssd1 vccd1 vccd1 _27079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14044_ _26069_/Q _14369_/S _14042_/X _14043_/X vssd1 vssd1 vccd1 vccd1 _14044_/X
+ sky130_fd_sc_hd__o211a_1
X_18921_ _25548_/Q _18568_/A _18920_/X _19069_/A _18572_/A vssd1 vssd1 vccd1 vccd1
+ _18921_/X sky130_fd_sc_hd__a221o_1
XFILLER_106_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18852_ _18887_/B _19354_/B vssd1 vssd1 vccd1 vccd1 _18852_/Y sky130_fd_sc_hd__nor2_1
XFILLER_268_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17803_ _17813_/B _17803_/B vssd1 vssd1 vccd1 vccd1 _17803_/Y sky130_fd_sc_hd__nand2_1
XFILLER_269_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18783_ _18723_/X _18780_/X _18781_/X _18782_/X vssd1 vssd1 vccd1 vccd1 _18784_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_5760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15995_ _13010_/A _23549_/A _15994_/Y _13756_/B vssd1 vssd1 vccd1 vccd1 _15995_/X
+ sky130_fd_sc_hd__o211a_2
XTAP_5771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17734_ _17697_/A _17681_/A _17685_/A vssd1 vssd1 vccd1 vccd1 _17762_/A sky130_fd_sc_hd__a21oi_2
XFILLER_85_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14946_ _26548_/Q _26156_/Q _14970_/S vssd1 vssd1 vccd1 vccd1 _14946_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17665_ _19914_/A _19910_/A vssd1 vssd1 vccd1 vccd1 _19589_/A sky130_fd_sc_hd__nand2_2
XFILLER_36_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14877_ _14875_/X _14876_/X _14877_/S vssd1 vssd1 vccd1 vccd1 _14877_/X sky130_fd_sc_hd__mux2_1
XFILLER_223_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_101 _21490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_112 _21946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19404_ _26970_/Q _18764_/X _18765_/X _27002_/Q vssd1 vssd1 vccd1 vccd1 _19404_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_224_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16616_ _19045_/A _19048_/A vssd1 vssd1 vccd1 vccd1 _19046_/A sky130_fd_sc_hd__xnor2_4
XINSDIODE2_123 _23520_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13828_ _15939_/A vssd1 vssd1 vccd1 vccd1 _15509_/A sky130_fd_sc_hd__buf_4
XFILLER_91_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_134 _17592_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17596_ _17634_/A vssd1 vssd1 vccd1 vccd1 _17615_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_145 _13304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_156 _15800_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19335_ _27032_/Q _19063_/X _19334_/X _18565_/X vssd1 vssd1 vccd1 vccd1 _19335_/X
+ sky130_fd_sc_hd__a22o_1
XINSDIODE2_167 _19887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16547_ _14790_/X _23609_/A _16546_/X _16282_/A vssd1 vssd1 vccd1 vccd1 _19472_/A
+ sky130_fd_sc_hd__o211ai_4
XINSDIODE2_178 _15588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13759_ _25877_/Q _16419_/B vssd1 vssd1 vccd1 vccd1 _13759_/X sky130_fd_sc_hd__or2_1
XINSDIODE2_189 _19769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19266_ _17317_/X _18444_/X _19263_/X _19265_/X _18469_/X vssd1 vssd1 vccd1 vccd1
+ _19266_/X sky130_fd_sc_hd__o221a_1
X_16478_ _25860_/Q _26060_/Q _16500_/S vssd1 vssd1 vccd1 vccd1 _16478_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18217_ _19583_/A vssd1 vssd1 vccd1 vccd1 _19018_/A sky130_fd_sc_hd__clkbuf_2
X_15429_ _16360_/S _15427_/X _15428_/X _13467_/A vssd1 vssd1 vccd1 vccd1 _15430_/B
+ sky130_fd_sc_hd__a31o_1
X_19197_ _25524_/Q _18556_/X _18557_/X _17418_/A vssd1 vssd1 vccd1 vccd1 _19197_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_117_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18148_ _18721_/A vssd1 vssd1 vccd1 vccd1 _18968_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18079_ _18369_/A _18603_/A _18079_/S vssd1 vssd1 vccd1 vccd1 _18080_/B sky130_fd_sc_hd__mux2_1
XFILLER_160_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20110_ _19991_/X _20109_/X _20052_/X vssd1 vssd1 vccd1 vccd1 _20110_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_236_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21090_ _21090_/A vssd1 vssd1 vccd1 vccd1 _25905_/D sky130_fd_sc_hd__clkbuf_1
X_20041_ _20007_/B _20038_/X _20040_/X vssd1 vssd1 vccd1 vccd1 _20042_/B sky130_fd_sc_hd__a21oi_1
XFILLER_259_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23800_ _23800_/A vssd1 vssd1 vccd1 vccd1 _26784_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24780_ _27101_/Q _24798_/B vssd1 vssd1 vccd1 vccd1 _24780_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21992_ _26109_/Q _20913_/X _21994_/S vssd1 vssd1 vccd1 vccd1 _21993_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23731_ _23731_/A vssd1 vssd1 vccd1 vccd1 _23731_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_242_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20943_ _25851_/Q _20942_/X _20949_/S vssd1 vssd1 vccd1 vccd1 _20944_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26450_ _26483_/CLK _26450_/D vssd1 vssd1 vccd1 vccd1 _26450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23662_ _23662_/A vssd1 vssd1 vccd1 vccd1 _26737_/D sky130_fd_sc_hd__clkbuf_1
X_20874_ _20874_/A vssd1 vssd1 vccd1 vccd1 _25829_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25401_ _25401_/A vssd1 vssd1 vccd1 vccd1 _27297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22613_ _25027_/A vssd1 vssd1 vccd1 vccd1 _24835_/A sky130_fd_sc_hd__buf_8
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26381_ _26609_/CLK _26381_/D vssd1 vssd1 vccd1 vccd1 _26381_/Q sky130_fd_sc_hd__dfxtp_1
X_23593_ _23593_/A vssd1 vssd1 vccd1 vccd1 _26709_/D sky130_fd_sc_hd__clkbuf_1
X_25332_ _27267_/Q _23699_/A _25332_/S vssd1 vssd1 vccd1 vccd1 _25333_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22544_ _22538_/X _22543_/Y _24770_/A vssd1 vssd1 vccd1 vccd1 _26294_/D sky130_fd_sc_hd__a21oi_1
XFILLER_210_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25263_ _23702_/X _27236_/Q _25271_/S vssd1 vssd1 vccd1 vccd1 _25264_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22475_ _22475_/A vssd1 vssd1 vccd1 vccd1 _26263_/D sky130_fd_sc_hd__clkbuf_1
X_27002_ _27004_/CLK _27002_/D vssd1 vssd1 vccd1 vccd1 _27002_/Q sky130_fd_sc_hd__dfxtp_1
X_24214_ _24222_/A _24214_/B _24215_/B vssd1 vssd1 vccd1 vccd1 _26961_/D sky130_fd_sc_hd__nor3_1
XFILLER_194_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21426_ _21420_/Y _21424_/X _21425_/X vssd1 vssd1 vccd1 vccd1 _21426_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25194_ _24674_/B _25189_/X _25187_/X _27207_/Q _25191_/X vssd1 vssd1 vccd1 vccd1
+ _27207_/D sky130_fd_sc_hd__o221a_1
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21357_ _21357_/A vssd1 vssd1 vccd1 vccd1 _21357_/Y sky130_fd_sc_hd__inv_2
X_24145_ _24145_/A vssd1 vssd1 vccd1 vccd1 _26938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20308_ _19231_/A _20092_/A _19249_/X _20376_/A vssd1 vssd1 vccd1 vccd1 _20308_/Y
+ sky130_fd_sc_hd__a22oi_2
X_21288_ _21284_/X _18246_/X _21286_/X _25800_/Q _21641_/B vssd1 vssd1 vccd1 vccd1
+ _21288_/X sky130_fd_sc_hd__a221o_1
XFILLER_151_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24076_ _25321_/A _25393_/B vssd1 vssd1 vccd1 vccd1 _24133_/A sky130_fd_sc_hd__nor2_2
XFILLER_1_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23027_ _23027_/A vssd1 vssd1 vccd1 vccd1 _26484_/D sky130_fd_sc_hd__clkbuf_1
X_20239_ _20237_/X _20238_/Y _19748_/X vssd1 vssd1 vccd1 vccd1 _20239_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14800_ _15424_/A vssd1 vssd1 vccd1 vccd1 _14801_/A sky130_fd_sc_hd__clkbuf_4
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _13346_/A _15778_/X _15779_/X _13366_/A vssd1 vssd1 vccd1 vccd1 _15780_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_188_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12992_ _12992_/A _13068_/A vssd1 vssd1 vccd1 vccd1 _13012_/A sky130_fd_sc_hd__nor2_4
X_24978_ _24978_/A _24978_/B vssd1 vssd1 vccd1 vccd1 _24978_/Y sky130_fd_sc_hd__nand2_1
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26717_ _26878_/CLK _26717_/D vssd1 vssd1 vccd1 vccd1 _26717_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14731_ _15095_/S vssd1 vssd1 vccd1 vccd1 _15004_/S sky130_fd_sc_hd__buf_2
XFILLER_57_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23929_ _23929_/A vssd1 vssd1 vccd1 vccd1 _26842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _22633_/A _22415_/A vssd1 vssd1 vccd1 vccd1 _22536_/A sky130_fd_sc_hd__nor2_8
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26648_ _26744_/CLK _26648_/D vssd1 vssd1 vccd1 vccd1 _26648_/Q sky130_fd_sc_hd__dfxtp_1
X_14662_ _14662_/A vssd1 vssd1 vccd1 vccd1 _14662_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _16399_/X _16400_/X _16401_/S vssd1 vssd1 vccd1 vccd1 _16401_/X sky130_fd_sc_hd__mux2_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13613_ _14268_/S vssd1 vssd1 vccd1 vccd1 _13614_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_260_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17381_ _25546_/Q _17381_/B vssd1 vssd1 vccd1 vccd1 _17389_/C sky130_fd_sc_hd__and2_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26579_ _26903_/CLK _26579_/D vssd1 vssd1 vccd1 vccd1 _26579_/Q sky130_fd_sc_hd__dfxtp_1
X_14593_ _14593_/A vssd1 vssd1 vccd1 vccd1 _14593_/X sky130_fd_sc_hd__buf_2
XFILLER_186_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19120_ _25618_/Q _18971_/X _19119_/X _19007_/X vssd1 vssd1 vccd1 vccd1 _25618_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_201_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16332_ _15071_/X _16296_/Y _16331_/Y _15830_/A vssd1 vssd1 vccd1 vccd1 _16332_/X
+ sky130_fd_sc_hd__a211o_2
X_13544_ _13532_/X _13536_/X _13542_/X _14816_/A vssd1 vssd1 vccd1 vccd1 _13544_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19051_ _16125_/A _18366_/A _18731_/Y _18602_/A _19050_/X vssd1 vssd1 vccd1 vccd1
+ _19051_/X sky130_fd_sc_hd__o221a_1
XFILLER_200_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16263_ _15110_/A _26611_/Q _15414_/A _26351_/Q _13347_/A vssd1 vssd1 vccd1 vccd1
+ _16263_/X sky130_fd_sc_hd__o221a_1
X_13475_ _13475_/A vssd1 vssd1 vccd1 vccd1 _13762_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_201_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18002_ _18008_/A vssd1 vssd1 vccd1 vccd1 _18003_/A sky130_fd_sc_hd__inv_2
X_15214_ _25853_/Q _26053_/Q _16436_/S vssd1 vssd1 vccd1 vccd1 _15214_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16194_ _27284_/Q _26477_/Q _16194_/S vssd1 vssd1 vccd1 vccd1 _16194_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15145_ _14859_/X _15140_/X _15144_/X _15020_/X vssd1 vssd1 vccd1 vccd1 _15145_/X
+ sky130_fd_sc_hd__a211o_1
Xoutput308 _16740_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[12] sky130_fd_sc_hd__buf_2
XFILLER_127_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput319 _16767_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[22] sky130_fd_sc_hd__buf_2
XFILLER_114_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15076_ _14601_/X _15074_/Y _15075_/X vssd1 vssd1 vccd1 vccd1 _15076_/X sky130_fd_sc_hd__o21a_1
X_19953_ _19879_/X _19951_/Y _19952_/X _19890_/X vssd1 vssd1 vccd1 vccd1 _19953_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_142_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14027_ _12892_/A _14133_/A _14026_/X _14029_/B _25923_/Q vssd1 vssd1 vccd1 vccd1
+ _15871_/B sky130_fd_sc_hd__o32a_2
X_18904_ _18904_/A vssd1 vssd1 vccd1 vccd1 _19049_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19884_ _25733_/Q vssd1 vssd1 vccd1 vccd1 _20648_/A sky130_fd_sc_hd__buf_8
XFILLER_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18835_ _20008_/A _19374_/B vssd1 vssd1 vccd1 vccd1 _18835_/Y sky130_fd_sc_hd__nor2_1
XFILLER_228_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18766_ _26953_/Q _18764_/X _18765_/X _26985_/Q vssd1 vssd1 vccd1 vccd1 _18766_/X
+ sky130_fd_sc_hd__a22o_1
X_15978_ _26792_/Q _26436_/Q _15980_/S vssd1 vssd1 vccd1 vccd1 _15978_/X sky130_fd_sc_hd__mux2_1
XFILLER_282_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17717_ _18757_/A vssd1 vssd1 vccd1 vccd1 _19302_/B sky130_fd_sc_hd__clkbuf_2
X_14929_ _14904_/Y _14911_/Y _14790_/X _14928_/Y vssd1 vssd1 vccd1 vccd1 _14929_/X
+ sky130_fd_sc_hd__o211a_1
X_18697_ _27016_/Q _18514_/X _18696_/X _18455_/X vssd1 vssd1 vccd1 vccd1 _18697_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17648_ _17592_/A _17653_/B _13918_/X _17597_/X _25932_/Q vssd1 vssd1 vccd1 vccd1
+ _17648_/Y sky130_fd_sc_hd__o32ai_4
XFILLER_63_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17579_ _17669_/B _17564_/X _17572_/X _17578_/X vssd1 vssd1 vccd1 vccd1 _17580_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_251_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19318_ _19449_/A _19318_/B vssd1 vssd1 vccd1 vccd1 _19318_/Y sky130_fd_sc_hd__nand2_1
X_20590_ _20590_/A vssd1 vssd1 vccd1 vccd1 _25715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19249_ _19283_/B _19249_/B vssd1 vssd1 vccd1 vccd1 _19249_/X sky130_fd_sc_hd__or2_2
XFILLER_164_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22260_ _26198_/Q _22249_/X _22255_/X _26299_/Q _22256_/X vssd1 vssd1 vccd1 vccd1
+ _22260_/X sky130_fd_sc_hd__a221o_1
XFILLER_192_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21211_ _21870_/A _21562_/C _22536_/A vssd1 vssd1 vccd1 vccd1 _21211_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_158_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27110_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22191_ _26181_/Q _22185_/X _22190_/X _22181_/X vssd1 vssd1 vccd1 vccd1 _26181_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21142_ _25920_/Q _21130_/X _21131_/X input19/X vssd1 vssd1 vccd1 vccd1 _21143_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25950_ _25985_/CLK _25950_/D vssd1 vssd1 vccd1 vccd1 _25950_/Q sky130_fd_sc_hd__dfxtp_1
X_21073_ _21166_/A vssd1 vssd1 vccd1 vccd1 _21112_/A sky130_fd_sc_hd__buf_4
XFILLER_160_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24901_ _24941_/A vssd1 vssd1 vccd1 vccd1 _24902_/A sky130_fd_sc_hd__clkbuf_2
X_20024_ _19999_/A _19999_/Y _20022_/Y _20023_/X vssd1 vssd1 vccd1 vccd1 _20024_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25881_ _27275_/CLK _25881_/D vssd1 vssd1 vccd1 vccd1 _25881_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24832_ _24828_/Y _24831_/X _24816_/X vssd1 vssd1 vccd1 vccd1 _27113_/D sky130_fd_sc_hd__a21oi_1
XFILLER_100_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24763_ _27097_/Q _24744_/X _25155_/A _24720_/A vssd1 vssd1 vccd1 vccd1 _24764_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_21975_ _26101_/Q _20887_/X _21983_/S vssd1 vssd1 vccd1 vccd1 _21976_/A sky130_fd_sc_hd__mux2_1
XFILLER_255_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26502_ _27309_/CLK _26502_/D vssd1 vssd1 vccd1 vccd1 _26502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23714_ _23714_/A vssd1 vssd1 vccd1 vccd1 _26756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20926_ _23741_/A vssd1 vssd1 vccd1 vccd1 _20926_/X sky130_fd_sc_hd__clkbuf_2
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24694_ _27081_/Q _24680_/X _24693_/Y _24676_/X vssd1 vssd1 vccd1 vccd1 _24695_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_215_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26433_ _26433_/CLK _26433_/D vssd1 vssd1 vccd1 vccd1 _26433_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23645_ _26730_/Q _23555_/X _23645_/S vssd1 vssd1 vccd1 vccd1 _23646_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20857_ _20857_/A vssd1 vssd1 vccd1 vccd1 _25824_/D sky130_fd_sc_hd__clkbuf_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26364_ _27267_/CLK _26364_/D vssd1 vssd1 vccd1 vccd1 _26364_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_179_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23576_ _26704_/Q _23574_/X _23588_/S vssd1 vssd1 vccd1 vccd1 _23577_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20788_ _20788_/A vssd1 vssd1 vccd1 vccd1 _25789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25315_ _23779_/X _27260_/Q _25315_/S vssd1 vssd1 vccd1 vccd1 _25316_/A sky130_fd_sc_hd__mux2_1
X_22527_ _22527_/A vssd1 vssd1 vccd1 vccd1 _26287_/D sky130_fd_sc_hd__clkbuf_1
X_26295_ _26297_/CLK _26295_/D vssd1 vssd1 vccd1 vccd1 _26295_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13260_ _15938_/S vssd1 vssd1 vccd1 vccd1 _13829_/S sky130_fd_sc_hd__clkbuf_4
X_25246_ _27229_/Q _25175_/X _25245_/X _19758_/X vssd1 vssd1 vccd1 vccd1 _27229_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22458_ _26207_/Q _22446_/X _22457_/X _22455_/X vssd1 vssd1 vccd1 vccd1 _26255_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21409_ input46/X input81/X _21422_/S vssd1 vssd1 vccd1 vccd1 _21410_/A sky130_fd_sc_hd__mux2_8
X_13191_ _23363_/B _13365_/A _13209_/A _20485_/A _13190_/Y vssd1 vssd1 vccd1 vccd1
+ _13204_/B sky130_fd_sc_hd__o221a_1
X_25177_ _25190_/A vssd1 vssd1 vccd1 vccd1 _25178_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22389_ _22362_/B _22385_/X _22388_/Y vssd1 vssd1 vccd1 vccd1 _22389_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24128_ _24128_/A vssd1 vssd1 vccd1 vccd1 _26930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_269_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24059_ _26900_/Q _23587_/X _24059_/S vssd1 vssd1 vccd1 vccd1 _24060_/A sky130_fd_sc_hd__mux2_1
X_16950_ _16950_/A vssd1 vssd1 vccd1 vccd1 _16950_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15901_ _26077_/Q _25882_/Q _15902_/S vssd1 vssd1 vccd1 vccd1 _15901_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16881_ _16881_/A vssd1 vssd1 vccd1 vccd1 _16881_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_265_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18620_ _25542_/Q _18459_/A _18619_/X _17688_/A _18466_/A vssd1 vssd1 vccd1 vccd1
+ _18620_/X sky130_fd_sc_hd__a221o_1
XFILLER_77_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15832_ _18076_/A _15868_/B _15244_/A _15831_/X vssd1 vssd1 vccd1 vccd1 _17831_/A
+ sky130_fd_sc_hd__o22a_4
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _15491_/A _27278_/Q _26471_/Q _15501_/A _13775_/A vssd1 vssd1 vccd1 vccd1
+ _15763_/X sky130_fd_sc_hd__a221o_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18551_ _18495_/A _18547_/X _18550_/X vssd1 vssd1 vccd1 vccd1 _18551_/Y sky130_fd_sc_hd__o21ai_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _12975_/A _12975_/B _25470_/Q vssd1 vssd1 vccd1 vccd1 _14401_/A sky130_fd_sc_hd__nor3b_2
XFILLER_218_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _15994_/A vssd1 vssd1 vccd1 vccd1 _15830_/A sky130_fd_sc_hd__buf_4
X_17502_ _18036_/A vssd1 vssd1 vccd1 vccd1 _18307_/A sky130_fd_sc_hd__buf_4
XFILLER_205_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18482_ _18482_/A _18482_/B vssd1 vssd1 vccd1 vccd1 _19573_/A sky130_fd_sc_hd__xnor2_2
XFILLER_206_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15694_ _15694_/A _15694_/B vssd1 vssd1 vccd1 vccd1 _15694_/Y sky130_fd_sc_hd__nor2_1
XFILLER_261_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _24239_/A vssd1 vssd1 vccd1 vccd1 _24164_/A sky130_fd_sc_hd__buf_2
XFILLER_72_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14645_ _26938_/Q _16467_/A vssd1 vssd1 vccd1 vccd1 _14645_/X sky130_fd_sc_hd__or2_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17364_ _25540_/Q _17362_/B _17363_/Y vssd1 vssd1 vccd1 vccd1 _25540_/D sky130_fd_sc_hd__o21a_1
XFILLER_242_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14576_ _13801_/Y _16729_/B _18549_/S vssd1 vssd1 vccd1 vccd1 _16732_/B sky130_fd_sc_hd__a21oi_4
XFILLER_202_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16315_ _26677_/Q _25717_/Q _16315_/S vssd1 vssd1 vccd1 vccd1 _16315_/X sky130_fd_sc_hd__mux2_1
X_19103_ _19234_/A _19103_/B _19103_/C vssd1 vssd1 vccd1 vccd1 _19103_/X sky130_fd_sc_hd__or3_4
X_13527_ _15859_/A vssd1 vssd1 vccd1 vccd1 _15836_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17295_ _24966_/A vssd1 vssd1 vccd1 vccd1 _17334_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_201_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19034_ _19034_/A _19034_/B vssd1 vssd1 vccd1 vccd1 _19042_/B sky130_fd_sc_hd__xnor2_4
X_16246_ _15020_/X _16241_/X _16245_/X _14679_/A vssd1 vssd1 vccd1 vccd1 _16246_/X
+ sky130_fd_sc_hd__o211a_1
X_13458_ _25595_/Q _13756_/B vssd1 vssd1 vccd1 vccd1 _13458_/X sky130_fd_sc_hd__or2_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16177_ _16175_/X _16176_/X _16183_/S vssd1 vssd1 vccd1 vccd1 _16177_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13389_ _13389_/A _13389_/B vssd1 vssd1 vccd1 vccd1 _13389_/Y sky130_fd_sc_hd__nor2_1
XFILLER_182_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15128_ _14790_/X _23594_/A _15126_/X _16282_/A vssd1 vssd1 vccd1 vccd1 _19309_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_114_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15059_ _25855_/Q _26055_/Q _16223_/S vssd1 vssd1 vccd1 vccd1 _15059_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19936_ _19930_/A _19870_/B _19935_/X _24810_/A vssd1 vssd1 vccd1 vccd1 _19936_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_123_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19867_ _19839_/A _27074_/Q _19866_/X vssd1 vssd1 vccd1 vccd1 _19867_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18818_ _27082_/Q _18815_/X _18816_/X _27180_/Q _18817_/X vssd1 vssd1 vccd1 vccd1
+ _18818_/X sky130_fd_sc_hd__a221o_1
XFILLER_228_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19798_ _19798_/A _20249_/B vssd1 vssd1 vccd1 vccd1 _19823_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18749_ _18813_/A vssd1 vssd1 vccd1 vccd1 _19462_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_209_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21760_ _21760_/A vssd1 vssd1 vccd1 vccd1 _26013_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_252_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20711_ _27102_/Q _19691_/X _20710_/X vssd1 vssd1 vccd1 vccd1 _20712_/C sky130_fd_sc_hd__o21ai_1
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21691_ _21691_/A vssd1 vssd1 vccd1 vccd1 _25984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23430_ _26649_/Q _23130_/X _23430_/S vssd1 vssd1 vccd1 vccd1 _23431_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20642_ _26268_/Q _20633_/X _20641_/X _20631_/X vssd1 vssd1 vccd1 vccd1 _25731_/D
+ sky130_fd_sc_hd__o211a_1
X_23361_ _20621_/X _26619_/Q _23361_/S vssd1 vssd1 vccd1 vccd1 _23362_/A sky130_fd_sc_hd__mux2_1
X_20573_ _20573_/A vssd1 vssd1 vccd1 vccd1 _25711_/D sky130_fd_sc_hd__clkbuf_1
X_25100_ _24715_/Y _25097_/X _25099_/Y _25082_/X vssd1 vssd1 vccd1 vccd1 _25100_/X
+ sky130_fd_sc_hd__a31o_1
X_22312_ _26216_/Q _22299_/X _22311_/X _22304_/X vssd1 vssd1 vccd1 vccd1 _26216_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26080_ _27282_/CLK _26080_/D vssd1 vssd1 vccd1 vccd1 _26080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23292_ _23348_/A vssd1 vssd1 vccd1 vccd1 _23361_/S sky130_fd_sc_hd__buf_6
XFILLER_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25031_ _25138_/A vssd1 vssd1 vccd1 vccd1 _25031_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22243_ _22288_/A vssd1 vssd1 vccd1 vccd1 _22243_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22174_ _26175_/Q _22169_/X _22173_/X _22164_/X vssd1 vssd1 vccd1 vccd1 _26175_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21125_ _21136_/A _21125_/B vssd1 vssd1 vccd1 vccd1 _21126_/A sky130_fd_sc_hd__or2_1
X_26982_ _27001_/CLK _26982_/D vssd1 vssd1 vccd1 vccd1 _26982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25933_ _27221_/CLK _25933_/D vssd1 vssd1 vccd1 vccd1 _25933_/Q sky130_fd_sc_hd__dfxtp_2
X_21056_ _21056_/A vssd1 vssd1 vccd1 vccd1 _25896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20007_ _20007_/A _20007_/B vssd1 vssd1 vccd1 vccd1 _20014_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25864_ _25867_/CLK _25864_/D vssd1 vssd1 vccd1 vccd1 _25864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_55_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27305_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_207_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24815_ _20643_/A _24810_/X _24674_/Y _24811_/X vssd1 vssd1 vccd1 vccd1 _24815_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25795_ _25796_/CLK _25795_/D vssd1 vssd1 vccd1 vccd1 _25795_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24746_ _24768_/A _24746_/B vssd1 vssd1 vccd1 vccd1 _24746_/Y sky130_fd_sc_hd__nand2_4
X_12760_ _17443_/A _12760_/B _17444_/D _20487_/A vssd1 vssd1 vccd1 vccd1 _12762_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_261_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21958_ _21958_/A vssd1 vssd1 vccd1 vccd1 _26094_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_opt_8_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_8_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_270_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20909_ _20909_/A vssd1 vssd1 vccd1 vccd1 _25840_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24677_ _27077_/Q _24657_/X _24674_/Y _24676_/X vssd1 vssd1 vccd1 vccd1 _24678_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_12691_ _17504_/A _17971_/A _18006_/B vssd1 vssd1 vccd1 vccd1 _17679_/A sky130_fd_sc_hd__or3_1
X_21889_ _25249_/B _23788_/B vssd1 vssd1 vccd1 vccd1 _21946_/A sky130_fd_sc_hd__or2_4
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _13082_/A _26685_/Q _26813_/Q _14095_/A _13121_/B vssd1 vssd1 vccd1 vccd1
+ _14431_/C sky130_fd_sc_hd__a221o_1
X_26416_ _27287_/CLK _26416_/D vssd1 vssd1 vccd1 vccd1 _26416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23628_ _26722_/Q _23530_/X _23634_/S vssd1 vssd1 vccd1 vccd1 _23629_/A sky130_fd_sc_hd__mux2_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14361_ _14443_/A _16816_/B _14360_/Y _14362_/B vssd1 vssd1 vccd1 vccd1 _14361_/X
+ sky130_fd_sc_hd__a211o_1
X_26347_ _26796_/CLK _26347_/D vssd1 vssd1 vccd1 vccd1 _26347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23559_ _23591_/A vssd1 vssd1 vccd1 vccd1 _23572_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_183_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 core_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_1
X_16100_ _14729_/A _16098_/X _16099_/X _13467_/A vssd1 vssd1 vccd1 vccd1 _16100_/X
+ sky130_fd_sc_hd__a31o_1
X_13312_ _13543_/A vssd1 vssd1 vccd1 vccd1 _13313_/A sky130_fd_sc_hd__buf_4
X_17080_ _26235_/Q _26234_/Q vssd1 vssd1 vccd1 vccd1 _17091_/C sky130_fd_sc_hd__or2_1
Xinput29 core_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_1
X_14292_ _14535_/A _14292_/B _14292_/C vssd1 vssd1 vccd1 vccd1 _14292_/X sky130_fd_sc_hd__or3_1
X_26278_ _26278_/CLK _26278_/D vssd1 vssd1 vccd1 vccd1 _26278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16031_ _25736_/Q _19971_/A _16031_/S vssd1 vssd1 vccd1 vccd1 _16632_/B sky130_fd_sc_hd__mux2_1
X_25229_ _27059_/Q _21874_/A input183/X _25214_/X _25178_/A vssd1 vssd1 vccd1 vccd1
+ _25229_/X sky130_fd_sc_hd__a41o_1
X_13243_ _14791_/A _13229_/X _13236_/X _13242_/X vssd1 vssd1 vccd1 vccd1 _13276_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13174_ _13174_/A vssd1 vssd1 vccd1 vccd1 _14590_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_123_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17982_ _18416_/S _17977_/X _17981_/Y vssd1 vssd1 vccd1 vccd1 _18487_/B sky130_fd_sc_hd__o21ai_1
XFILLER_112_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19721_ _20225_/A vssd1 vssd1 vccd1 vccd1 _19721_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_278_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16933_ _16909_/X _16883_/B _16882_/X _16910_/X _16911_/X vssd1 vssd1 vccd1 vccd1
+ _16933_/X sky130_fd_sc_hd__o221a_1
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19652_ _19652_/A vssd1 vssd1 vccd1 vccd1 _20100_/A sky130_fd_sc_hd__buf_2
X_16864_ _16864_/A _16864_/B vssd1 vssd1 vccd1 vccd1 _16865_/A sky130_fd_sc_hd__and2_1
XFILLER_253_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18603_ _18603_/A vssd1 vssd1 vccd1 vccd1 _18643_/A sky130_fd_sc_hd__buf_2
XFILLER_92_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15815_ _15813_/X _15814_/X _15826_/S vssd1 vssd1 vccd1 vccd1 _15815_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16795_ _17856_/A _16887_/A _16794_/Y _16853_/A _16697_/D vssd1 vssd1 vccd1 vccd1
+ _17055_/D sky130_fd_sc_hd__a221o_4
X_19583_ _19583_/A _19583_/B vssd1 vssd1 vccd1 vccd1 _19583_/Y sky130_fd_sc_hd__nand2_1
XFILLER_234_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15746_ _14713_/A _15733_/X _15737_/X _15745_/X _13876_/X vssd1 vssd1 vccd1 vccd1
+ _15746_/X sky130_fd_sc_hd__a311o_1
X_18534_ _19256_/A _18483_/A _18501_/X _18533_/X vssd1 vssd1 vccd1 vccd1 _18534_/X
+ sky130_fd_sc_hd__a211o_1
X_12958_ _12959_/A _25475_/Q vssd1 vssd1 vccd1 vccd1 _20868_/A sky130_fd_sc_hd__nor2b_4
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18465_ _18465_/A vssd1 vssd1 vccd1 vccd1 _18466_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15677_ _15676_/X _27279_/Q _26472_/Q _15674_/X _13281_/A vssd1 vssd1 vccd1 vccd1
+ _15677_/X sky130_fd_sc_hd__a221o_1
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12889_ _12941_/A _13569_/C _13569_/A vssd1 vssd1 vccd1 vccd1 _15706_/C sky130_fd_sc_hd__a21oi_1
XFILLER_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17416_ _17418_/A _17418_/C _17415_/Y vssd1 vssd1 vccd1 vccd1 _25556_/D sky130_fd_sc_hd__o21a_1
XFILLER_221_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14628_ _14969_/S vssd1 vssd1 vccd1 vccd1 _14952_/S sky130_fd_sc_hd__buf_2
X_18396_ _27138_/Q vssd1 vssd1 vccd1 vccd1 _19790_/A sky130_fd_sc_hd__buf_4
XFILLER_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17347_ _25535_/Q vssd1 vssd1 vccd1 vccd1 _17347_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14559_ _13465_/A _23508_/A _14558_/X _13683_/A vssd1 vssd1 vccd1 vccd1 _14559_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_158_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17278_ _25514_/Q vssd1 vssd1 vccd1 vccd1 _17278_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16229_ _14881_/A _16224_/X _16228_/Y _15187_/X vssd1 vssd1 vccd1 vccd1 _16229_/X
+ sky130_fd_sc_hd__o211a_1
X_19017_ _18861_/X _19016_/X _15529_/A vssd1 vssd1 vccd1 vccd1 _19018_/D sky130_fd_sc_hd__a21oi_2
XFILLER_174_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19919_ _19889_/A _19919_/B vssd1 vssd1 vccd1 vccd1 _19923_/A sky130_fd_sc_hd__and2b_1
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22930_ _26441_/Q _22698_/X _22934_/S vssd1 vssd1 vccd1 vccd1 _22931_/A sky130_fd_sc_hd__mux2_1
XFILLER_257_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22861_ _22861_/A vssd1 vssd1 vccd1 vccd1 _26410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24600_ _24600_/A _24608_/B vssd1 vssd1 vccd1 vccd1 _24600_/Y sky130_fd_sc_hd__nand2_1
X_21812_ _26036_/Q _20894_/X _21816_/S vssd1 vssd1 vccd1 vccd1 _21813_/A sky130_fd_sc_hd__mux2_1
X_25580_ _26684_/CLK _25580_/D vssd1 vssd1 vccd1 vccd1 _25580_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22792_ _26380_/Q _22707_/X _22800_/S vssd1 vssd1 vccd1 vccd1 _22793_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24531_ _24472_/X _25628_/Q _24530_/X vssd1 vssd1 vccd1 vccd1 _24768_/B sky130_fd_sc_hd__o21a_4
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21743_ _20529_/X _26006_/Q _21743_/S vssd1 vssd1 vccd1 vccd1 _21744_/A sky130_fd_sc_hd__mux2_1
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27250_ _27311_/CLK _27250_/D vssd1 vssd1 vccd1 vccd1 _27250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24462_ _26310_/Q _24455_/X _24456_/X input223/X _24457_/X vssd1 vssd1 vccd1 vccd1
+ _24462_/X sky130_fd_sc_hd__a221o_1
XFILLER_40_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21674_ _25977_/Q input212/X _21674_/S vssd1 vssd1 vccd1 vccd1 _21675_/A sky130_fd_sc_hd__mux2_1
XFILLER_269_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26201_ _26307_/CLK _26201_/D vssd1 vssd1 vccd1 vccd1 _26201_/Q sky130_fd_sc_hd__dfxtp_1
X_23413_ _26641_/Q _23105_/X _23419_/S vssd1 vssd1 vccd1 vccd1 _23414_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20625_ _26261_/Q _17190_/X _20624_/X _19965_/X vssd1 vssd1 vccd1 vccd1 _25724_/D
+ sky130_fd_sc_hd__o211a_1
X_27181_ _27196_/CLK _27181_/D vssd1 vssd1 vccd1 vccd1 _27181_/Q sky130_fd_sc_hd__dfxtp_1
X_24393_ _24455_/A vssd1 vssd1 vccd1 vccd1 _24393_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_102_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26186_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_26132_ _26592_/CLK _26132_/D vssd1 vssd1 vccd1 vccd1 _26132_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_138_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23344_ _20588_/X _26611_/Q _23346_/S vssd1 vssd1 vccd1 vccd1 _23345_/A sky130_fd_sc_hd__mux2_1
X_20556_ _20554_/X _25707_/Q _20572_/S vssd1 vssd1 vccd1 vccd1 _20557_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26063_ _26063_/CLK _26063_/D vssd1 vssd1 vccd1 vccd1 _26063_/Q sky130_fd_sc_hd__dfxtp_1
X_23275_ _26580_/Q _23127_/X _23277_/S vssd1 vssd1 vccd1 vccd1 _23276_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20487_ _20487_/A _20487_/B _20487_/C vssd1 vssd1 vccd1 vccd1 _21888_/C sky130_fd_sc_hd__or3_2
XFILLER_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25014_ _25142_/A vssd1 vssd1 vccd1 vccd1 _25014_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22226_ input8/X input283/X _22226_/S vssd1 vssd1 vccd1 vccd1 _22226_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22157_ _26170_/Q _22152_/X _22156_/X _22148_/X vssd1 vssd1 vccd1 vccd1 _26170_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_267_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput480 _25732_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[8] sky130_fd_sc_hd__buf_2
XFILLER_120_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21108_ _21108_/A vssd1 vssd1 vccd1 vccd1 _25910_/D sky130_fd_sc_hd__clkbuf_1
X_26965_ _26995_/CLK _26965_/D vssd1 vssd1 vccd1 vccd1 _26965_/Q sky130_fd_sc_hd__dfxtp_1
X_22088_ _26152_/Q _20948_/X _22088_/S vssd1 vssd1 vccd1 vccd1 _22089_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13930_ _14485_/B _14606_/C _13925_/Y _13929_/X vssd1 vssd1 vccd1 vccd1 _13930_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25916_ _27188_/CLK _25916_/D vssd1 vssd1 vccd1 vccd1 _25916_/Q sky130_fd_sc_hd__dfxtp_4
X_21039_ _21050_/A vssd1 vssd1 vccd1 vccd1 _21048_/S sky130_fd_sc_hd__clkbuf_4
X_26896_ _27253_/CLK _26896_/D vssd1 vssd1 vccd1 vccd1 _26896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13861_ _25804_/Q _15797_/B _13134_/A _13860_/X vssd1 vssd1 vccd1 vccd1 _13861_/X
+ sky130_fd_sc_hd__o211a_1
X_25847_ _26531_/CLK _25847_/D vssd1 vssd1 vccd1 vccd1 _25847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15600_ _15676_/A _26113_/Q _26014_/Q _16178_/S _15670_/A vssd1 vssd1 vccd1 vccd1
+ _15600_/X sky130_fd_sc_hd__a221o_1
X_12812_ _18001_/A _16594_/A vssd1 vssd1 vccd1 vccd1 _12813_/A sky130_fd_sc_hd__or2_1
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16580_ _16580_/A vssd1 vssd1 vccd1 vccd1 _17998_/A sky130_fd_sc_hd__clkbuf_4
XINSDIODE2_508 input270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13792_ _26528_/Q _26136_/Q _13792_/S vssd1 vssd1 vccd1 vccd1 _13792_/X sky130_fd_sc_hd__mux2_1
X_25778_ _27315_/CLK _25778_/D vssd1 vssd1 vccd1 vccd1 _25778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_519 _17023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15531_ _15245_/A _13567_/Y _14603_/A vssd1 vssd1 vccd1 vccd1 _15531_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12743_ _14431_/A vssd1 vssd1 vccd1 vccd1 _13884_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24729_ _24739_/A _24729_/B vssd1 vssd1 vccd1 vccd1 _24729_/Y sky130_fd_sc_hd__nand2_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ _19196_/A _18250_/B _18250_/C vssd1 vssd1 vccd1 vccd1 _18250_/X sky130_fd_sc_hd__or3_2
X_15462_ _15187_/A _15452_/X _15461_/X _13717_/A vssd1 vssd1 vccd1 vccd1 _15462_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_179_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12674_ _12674_/A vssd1 vssd1 vccd1 vccd1 _17444_/C sky130_fd_sc_hd__buf_4
XFILLER_231_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17201_ _17201_/A vssd1 vssd1 vccd1 vccd1 _25493_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14413_ _14409_/Y _14412_/X _12981_/A vssd1 vssd1 vccd1 vccd1 _14447_/B sky130_fd_sc_hd__o21ai_1
X_18181_ _18805_/A _18181_/B _18181_/C vssd1 vssd1 vccd1 vccd1 _18181_/X sky130_fd_sc_hd__or3_2
XFILLER_156_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15393_ _26640_/Q _26736_/Q _16086_/S vssd1 vssd1 vccd1 vccd1 _15394_/B sky130_fd_sc_hd__mux2_1
XFILLER_11_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17132_ _25473_/Q _17114_/X _17131_/Y _17120_/X vssd1 vssd1 vccd1 vccd1 _25473_/D
+ sky130_fd_sc_hd__o211a_1
X_14344_ _26654_/Q _25694_/Q _14344_/S vssd1 vssd1 vccd1 vccd1 _14344_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17063_ _17063_/A vssd1 vssd1 vccd1 vccd1 _17063_/X sky130_fd_sc_hd__buf_2
X_14275_ _13890_/A _26879_/Q _26751_/Q _14497_/A vssd1 vssd1 vccd1 vccd1 _14275_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16014_ _26532_/Q _26140_/Q _16014_/S vssd1 vssd1 vccd1 vccd1 _16015_/B sky130_fd_sc_hd__mux2_1
X_13226_ _15923_/S vssd1 vssd1 vccd1 vccd1 _16110_/S sky130_fd_sc_hd__buf_2
XFILLER_170_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13157_ _25880_/Q _16061_/B vssd1 vssd1 vccd1 vccd1 _13157_/X sky130_fd_sc_hd__or2_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13088_ _15904_/S vssd1 vssd1 vccd1 vccd1 _15971_/S sky130_fd_sc_hd__buf_4
X_17965_ _18683_/A _17918_/X _17964_/X vssd1 vssd1 vccd1 vccd1 _19454_/B sky130_fd_sc_hd__a21oi_2
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19704_ _19704_/A _19704_/B vssd1 vssd1 vccd1 vccd1 _19705_/B sky130_fd_sc_hd__or2_1
XFILLER_238_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16916_ _16916_/A _16927_/B vssd1 vssd1 vccd1 vccd1 _16968_/C sky130_fd_sc_hd__nor2_1
XFILLER_254_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17896_ _18347_/S vssd1 vssd1 vccd1 vccd1 _18416_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19635_ _19652_/A _19779_/A _24641_/A _17514_/A vssd1 vssd1 vccd1 vccd1 _20712_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_254_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16847_ _16847_/A vssd1 vssd1 vccd1 vccd1 _16847_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19566_ _20644_/A vssd1 vssd1 vccd1 vccd1 _19566_/X sky130_fd_sc_hd__buf_6
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16778_ _25686_/Q vssd1 vssd1 vccd1 vccd1 _22526_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_34_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18517_ _19839_/A _19261_/B vssd1 vssd1 vccd1 vccd1 _18517_/X sky130_fd_sc_hd__or2_1
XFILLER_209_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15729_ _13608_/X _15720_/X _15728_/X _14713_/C vssd1 vssd1 vccd1 vccd1 _15729_/X
+ sky130_fd_sc_hd__a211o_1
X_19497_ _25634_/Q _19497_/B vssd1 vssd1 vccd1 vccd1 _19497_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_0_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27287_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18448_ _27205_/Q _19364_/B _18447_/X vssd1 vssd1 vccd1 vccd1 _18448_/X sky130_fd_sc_hd__a21o_1
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18379_ _19772_/A _18432_/C vssd1 vssd1 vccd1 vccd1 _19768_/A sky130_fd_sc_hd__nand2_1
XFILLER_187_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20410_ _27129_/Q _19765_/X _20276_/X _20409_/Y vssd1 vssd1 vccd1 vccd1 _20410_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21390_ _22817_/A _21416_/B vssd1 vssd1 vccd1 vccd1 _21390_/X sky130_fd_sc_hd__or2_1
XFILLER_105_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20341_ _27158_/Q _27092_/Q vssd1 vssd1 vccd1 vccd1 _20342_/B sky130_fd_sc_hd__or2_1
XFILLER_161_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23060_ _23533_/A vssd1 vssd1 vccd1 vccd1 _23060_/X sky130_fd_sc_hd__clkbuf_4
X_20272_ _27155_/Q _20323_/B vssd1 vssd1 vccd1 vccd1 _20272_/Y sky130_fd_sc_hd__nand2_1
XFILLER_190_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22011_ _22011_/A vssd1 vssd1 vccd1 vccd1 _26117_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput208 localMemory_wb_adr_i[4] vssd1 vssd1 vccd1 vccd1 input208/X sky130_fd_sc_hd__clkbuf_1
Xinput219 localMemory_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input219/X sky130_fd_sc_hd__buf_6
XFILLER_271_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26750_ _26878_/CLK _26750_/D vssd1 vssd1 vccd1 vccd1 _26750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23962_ _23962_/A vssd1 vssd1 vccd1 vccd1 _26856_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25701_ _26595_/CLK _25701_/D vssd1 vssd1 vccd1 vccd1 _25701_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_84_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22913_ _22913_/A vssd1 vssd1 vccd1 vccd1 _26433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_257_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26681_ _26681_/CLK _26681_/D vssd1 vssd1 vccd1 vccd1 _26681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23893_ _23731_/X _26826_/Q _23893_/S vssd1 vssd1 vccd1 vccd1 _23894_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25632_ _26813_/CLK _25632_/D vssd1 vssd1 vccd1 vccd1 _25632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22844_ _22844_/A vssd1 vssd1 vccd1 vccd1 _26402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_271_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25563_ _27004_/CLK _25563_/D vssd1 vssd1 vccd1 vccd1 _25563_/Q sky130_fd_sc_hd__dfxtp_1
X_22775_ _22775_/A vssd1 vssd1 vccd1 vccd1 _26372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27302_ _27304_/CLK _27302_/D vssd1 vssd1 vccd1 vccd1 _27302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24514_ _27031_/Q _24506_/X _24513_/Y _24499_/X vssd1 vssd1 vccd1 vccd1 _27031_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21726_ _20496_/X _25998_/Q _21732_/S vssd1 vssd1 vccd1 vccd1 _21727_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25494_ _26940_/CLK _25494_/D vssd1 vssd1 vccd1 vccd1 _25494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27233_ _27297_/CLK _27233_/D vssd1 vssd1 vccd1 vccd1 _27233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24445_ _24472_/A _25612_/Q _24444_/X vssd1 vssd1 vccd1 vccd1 _24944_/A sky130_fd_sc_hd__o21ai_4
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21657_ _21657_/A vssd1 vssd1 vccd1 vccd1 _25969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27164_ _27164_/CLK _27164_/D vssd1 vssd1 vccd1 vccd1 _27164_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_149_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20608_ _23600_/A vssd1 vssd1 vccd1 vccd1 _23776_/A sky130_fd_sc_hd__clkbuf_4
X_24376_ _26296_/Q _24473_/A _24474_/A input240/X _24501_/A vssd1 vssd1 vccd1 vccd1
+ _24376_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21588_ _21586_/X _19308_/X _21587_/X _25823_/Q _21547_/X vssd1 vssd1 vccd1 vccd1
+ _21588_/X sky130_fd_sc_hd__a221o_1
XFILLER_137_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26115_ _26673_/CLK _26115_/D vssd1 vssd1 vccd1 vccd1 _26115_/Q sky130_fd_sc_hd__dfxtp_1
X_23327_ _20554_/X _26603_/Q _23335_/S vssd1 vssd1 vccd1 vccd1 _23328_/A sky130_fd_sc_hd__mux2_1
X_20539_ _20538_/X _25703_/Q _20551_/S vssd1 vssd1 vccd1 vccd1 _20540_/A sky130_fd_sc_hd__mux2_1
X_27095_ _27228_/CLK _27095_/D vssd1 vssd1 vccd1 vccd1 _27095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14060_ _14060_/A vssd1 vssd1 vccd1 vccd1 _14474_/S sky130_fd_sc_hd__buf_2
X_26046_ _27330_/A _26046_/D vssd1 vssd1 vccd1 vccd1 _26046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23258_ _26572_/Q _23101_/X _23266_/S vssd1 vssd1 vccd1 vccd1 _23259_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13011_ _13011_/A vssd1 vssd1 vccd1 vccd1 _15073_/A sky130_fd_sc_hd__buf_4
X_22209_ _26186_/Q _22200_/X _22208_/X _22195_/X vssd1 vssd1 vccd1 vccd1 _26186_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23189_ _23189_/A vssd1 vssd1 vccd1 vccd1 _26541_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_70_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26433_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_121_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17750_ _17750_/A _18111_/C vssd1 vssd1 vccd1 vccd1 _18108_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14962_ _14952_/S _14959_/X _14961_/X _14650_/X vssd1 vssd1 vccd1 vccd1 _14962_/X
+ sky130_fd_sc_hd__a211o_1
X_26948_ _26980_/CLK _26948_/D vssd1 vssd1 vccd1 vccd1 _26948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_282_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16701_ _22474_/A _16693_/X _18151_/B _16864_/A vssd1 vssd1 vccd1 vccd1 _16701_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13913_ _14489_/A vssd1 vssd1 vccd1 vccd1 _17556_/B sky130_fd_sc_hd__buf_2
XFILLER_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17681_ _17681_/A vssd1 vssd1 vccd1 vccd1 _19552_/A sky130_fd_sc_hd__clkbuf_4
X_14893_ _14890_/X _25858_/Q _26058_/Q _14984_/S _14754_/A vssd1 vssd1 vccd1 vccd1
+ _14893_/X sky130_fd_sc_hd__a221o_1
XFILLER_235_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26879_ _26880_/CLK _26879_/D vssd1 vssd1 vccd1 vccd1 _26879_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_262_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19420_ _20701_/A _19421_/B vssd1 vssd1 vccd1 vccd1 _19477_/B sky130_fd_sc_hd__nor2_1
XFILLER_262_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13844_ _13363_/A _13840_/X _13843_/X _13339_/A vssd1 vssd1 vccd1 vccd1 _13844_/X
+ sky130_fd_sc_hd__o211a_1
X_16632_ _17828_/A _16632_/B vssd1 vssd1 vccd1 vccd1 _16633_/A sky130_fd_sc_hd__and2_1
XFILLER_262_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_305 _25902_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_316 _19620_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_327 _19616_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19351_ _17444_/A _18972_/X _18973_/X _19350_/Y vssd1 vssd1 vccd1 vccd1 _19351_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_262_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13775_ _13775_/A vssd1 vssd1 vccd1 vccd1 _15486_/A sky130_fd_sc_hd__buf_2
XINSDIODE2_338 _19609_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16563_ _19385_/B vssd1 vssd1 vccd1 vccd1 _16575_/A sky130_fd_sc_hd__inv_2
XINSDIODE2_349 _19612_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18302_ _18806_/A _18290_/X _18301_/X vssd1 vssd1 vccd1 vccd1 _18302_/X sky130_fd_sc_hd__a21o_4
X_15514_ _27313_/Q _26570_/Q _15514_/S vssd1 vssd1 vccd1 vccd1 _15514_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12726_ _17992_/A vssd1 vssd1 vccd1 vccd1 _17995_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_128_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19282_ _19283_/A _19283_/B vssd1 vssd1 vccd1 vccd1 _19346_/C sky130_fd_sc_hd__and2_2
X_16494_ _27262_/Q _16501_/B vssd1 vssd1 vccd1 vccd1 _16494_/X sky130_fd_sc_hd__or2_1
XFILLER_128_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15445_ _25616_/Q _14595_/A _15444_/X _14616_/A vssd1 vssd1 vccd1 vccd1 _23568_/A
+ sky130_fd_sc_hd__o22a_4
X_18233_ _18812_/A vssd1 vssd1 vccd1 vccd1 _19056_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_90_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18164_ _27007_/Q _18116_/B _18161_/C _17742_/Y vssd1 vssd1 vccd1 vccd1 _18164_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_30_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15376_ _15374_/X _15375_/X _15376_/S vssd1 vssd1 vccd1 vccd1 _15376_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14327_ _14610_/A _14325_/X _14326_/Y vssd1 vssd1 vccd1 vccd1 _23517_/A sky130_fd_sc_hd__o21ai_4
XFILLER_184_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17115_ _17210_/A vssd1 vssd1 vccd1 vccd1 _17635_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_183_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18095_ _18805_/A vssd1 vssd1 vccd1 vccd1 _19196_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17046_ _17042_/X _16970_/B _16970_/C _17013_/X input235/X vssd1 vssd1 vccd1 vccd1
+ _17046_/X sky130_fd_sc_hd__a32o_4
X_14258_ _25872_/Q _14273_/B vssd1 vssd1 vccd1 vccd1 _14258_/X sky130_fd_sc_hd__or2_1
XFILLER_171_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13209_ _13209_/A vssd1 vssd1 vccd1 vccd1 _13210_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14189_ _14189_/A vssd1 vssd1 vccd1 vccd1 _17856_/A sky130_fd_sc_hd__buf_4
XFILLER_258_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _17673_/X _18995_/X _18996_/Y vssd1 vssd1 vccd1 vccd1 _18997_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _17946_/X _17947_/X _18067_/S vssd1 vssd1 vccd1 vccd1 _17948_/X sky130_fd_sc_hd__mux2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17879_ _17975_/A vssd1 vssd1 vccd1 vccd1 _18050_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_285_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19618_ _27053_/Q _21264_/A input171/X _19617_/X vssd1 vssd1 vccd1 vccd1 _19618_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20890_ _20890_/A vssd1 vssd1 vccd1 vccd1 _25834_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19549_ _25654_/Q _19549_/B vssd1 vssd1 vccd1 vccd1 _19549_/X sky130_fd_sc_hd__or2_1
XFILLER_41_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22560_ _26300_/Q _22565_/B vssd1 vssd1 vccd1 vccd1 _22560_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21511_ _21509_/X _19099_/X _21510_/X _25817_/Q _21483_/X vssd1 vssd1 vccd1 vccd1
+ _21511_/X sky130_fd_sc_hd__a221o_1
XFILLER_210_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22491_ _22491_/A _22491_/B vssd1 vssd1 vccd1 vccd1 _22492_/A sky130_fd_sc_hd__and2_1
XFILLER_166_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24230_ _26967_/Q _24233_/C vssd1 vssd1 vccd1 vccd1 _24231_/B sky130_fd_sc_hd__and2_1
Xclkbuf_4_15_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_15_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
X_21442_ _25950_/Q _21378_/X _21441_/Y _21400_/X vssd1 vssd1 vccd1 vccd1 _25950_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_148_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24161_ _24164_/A _24163_/B vssd1 vssd1 vccd1 vccd1 _24161_/Y sky130_fd_sc_hd__nor2_1
XFILLER_181_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21373_ input106/X input78/X _21422_/S vssd1 vssd1 vccd1 vccd1 _21374_/A sky130_fd_sc_hd__mux2_8
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23112_ _26511_/Q _23111_/X _23115_/S vssd1 vssd1 vccd1 vccd1 _23113_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20324_ _20219_/B _20321_/X _20339_/B _20323_/Y vssd1 vssd1 vccd1 vccd1 _20324_/X
+ sky130_fd_sc_hd__o31a_2
X_24092_ _26914_/Q _23530_/X _24098_/S vssd1 vssd1 vccd1 vccd1 _24093_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23043_ _23043_/A vssd1 vssd1 vccd1 vccd1 _26489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20255_ _20277_/A _20303_/B vssd1 vssd1 vccd1 vccd1 _20300_/C sky130_fd_sc_hd__xnor2_2
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20186_ _20186_/A vssd1 vssd1 vccd1 vccd1 _20186_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26802_ _27317_/CLK _26802_/D vssd1 vssd1 vccd1 vccd1 _26802_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24994_ _27166_/Q _24994_/B vssd1 vssd1 vccd1 vccd1 _24994_/X sky130_fd_sc_hd__and2_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26733_ _27308_/CLK _26733_/D vssd1 vssd1 vccd1 vccd1 _26733_/Q sky130_fd_sc_hd__dfxtp_1
X_23945_ _24002_/S vssd1 vssd1 vccd1 vccd1 _23954_/S sky130_fd_sc_hd__clkbuf_4
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26664_ _27276_/CLK _26664_/D vssd1 vssd1 vccd1 vccd1 _26664_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23876_ _23706_/X _26818_/Q _23882_/S vssd1 vssd1 vccd1 vccd1 _23877_/A sky130_fd_sc_hd__mux2_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25615_ _26940_/CLK _25615_/D vssd1 vssd1 vccd1 vccd1 _25615_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22827_ _26395_/Q _22653_/X _22829_/S vssd1 vssd1 vccd1 vccd1 _22828_/A sky130_fd_sc_hd__mux2_1
XFILLER_272_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26595_ _26595_/CLK _26595_/D vssd1 vssd1 vccd1 vccd1 _26595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25546_ _25547_/CLK _25546_/D vssd1 vssd1 vccd1 vccd1 _25546_/Q sky130_fd_sc_hd__dfxtp_1
X_13560_ input124/X input159/X _14320_/S vssd1 vssd1 vccd1 vccd1 _13561_/B sky130_fd_sc_hd__mux2_8
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22758_ _22815_/S vssd1 vssd1 vccd1 vccd1 _22767_/S sky130_fd_sc_hd__buf_2
XFILLER_213_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21709_ _21709_/A _21709_/B vssd1 vssd1 vccd1 vccd1 _25993_/D sky130_fd_sc_hd__nor2_1
X_13491_ _15759_/S vssd1 vssd1 vccd1 vccd1 _15758_/S sky130_fd_sc_hd__buf_2
XFILLER_157_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25477_ _26881_/CLK _25477_/D vssd1 vssd1 vccd1 vccd1 _25477_/Q sky130_fd_sc_hd__dfxtp_1
X_22689_ _26342_/Q _22688_/X _22689_/S vssd1 vssd1 vccd1 vccd1 _22690_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15230_ _14743_/A _26612_/Q _16354_/S _26352_/Q _16360_/S vssd1 vssd1 vccd1 vccd1
+ _15230_/X sky130_fd_sc_hd__o221a_1
X_24428_ _24392_/X _25609_/Q _24427_/X vssd1 vssd1 vccd1 vccd1 _24936_/A sky130_fd_sc_hd__o21ai_4
X_27216_ _27221_/CLK _27216_/D vssd1 vssd1 vccd1 vccd1 _27216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27147_ _27160_/CLK _27147_/D vssd1 vssd1 vccd1 vccd1 _27147_/Q sky130_fd_sc_hd__dfxtp_2
X_15161_ _26088_/Q _16242_/S _16308_/S _15160_/X vssd1 vssd1 vccd1 vccd1 _15161_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24359_ _24454_/A vssd1 vssd1 vccd1 vccd1 _24472_/A sky130_fd_sc_hd__buf_2
XFILLER_176_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14112_ _14107_/X _14108_/X _14110_/X _14111_/X vssd1 vssd1 vccd1 vccd1 _14112_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15092_ _16441_/S vssd1 vssd1 vccd1 vccd1 _15121_/S sky130_fd_sc_hd__buf_2
XFILLER_4_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27078_ _27176_/CLK _27078_/D vssd1 vssd1 vccd1 vccd1 _27078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18920_ _26956_/Q _18569_/A _18570_/A _26988_/Q vssd1 vssd1 vccd1 vccd1 _18920_/X
+ sky130_fd_sc_hd__a22o_1
X_26029_ _27265_/CLK _26029_/D vssd1 vssd1 vccd1 vccd1 _26029_/Q sky130_fd_sc_hd__dfxtp_2
X_14043_ _14043_/A vssd1 vssd1 vccd1 vccd1 _14043_/X sky130_fd_sc_hd__buf_2
XFILLER_268_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18851_ _18855_/A _18851_/B vssd1 vssd1 vccd1 vccd1 _18887_/B sky130_fd_sc_hd__xor2_4
XFILLER_268_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17802_ _17802_/A _17802_/B vssd1 vssd1 vccd1 vccd1 _17803_/B sky130_fd_sc_hd__or2_1
XFILLER_94_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18782_ _19003_/A vssd1 vssd1 vccd1 vccd1 _18782_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_282_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15994_ _15994_/A _15994_/B vssd1 vssd1 vccd1 vccd1 _15994_/Y sky130_fd_sc_hd__nor2_2
XTAP_5761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17733_ _25533_/Q _18458_/A _17731_/X _18172_/A _18465_/A vssd1 vssd1 vccd1 vccd1
+ _17733_/X sky130_fd_sc_hd__a221o_1
XFILLER_208_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14945_ _15014_/S vssd1 vssd1 vccd1 vccd1 _14970_/S sky130_fd_sc_hd__clkbuf_2
XTAP_5794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17664_ _19769_/B vssd1 vssd1 vccd1 vccd1 _19910_/A sky130_fd_sc_hd__buf_2
XFILLER_62_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14876_ _25858_/Q _26058_/Q _14876_/S vssd1 vssd1 vccd1 vccd1 _14876_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_102 _21504_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19403_ _27066_/Q _19055_/X _19400_/X _19402_/X _19066_/X vssd1 vssd1 vccd1 vccd1
+ _19403_/X sky130_fd_sc_hd__o221a_2
X_16615_ _19034_/A _19034_/B _19016_/S vssd1 vssd1 vccd1 vccd1 _19045_/A sky130_fd_sc_hd__o21ai_4
XFILLER_51_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_113 _21946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13827_ _13827_/A vssd1 vssd1 vccd1 vccd1 _15939_/A sky130_fd_sc_hd__buf_2
XINSDIODE2_124 _23556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_135 _17592_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17595_ _17595_/A _17595_/B vssd1 vssd1 vccd1 vccd1 _25580_/D sky130_fd_sc_hd__nor2_1
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_146 _13304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_157 _14725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19334_ _27160_/Q _19334_/B vssd1 vssd1 vccd1 vccd1 _19334_/X sky130_fd_sc_hd__or2_1
XFILLER_16_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13758_ _27271_/Q _26464_/Q _13792_/S vssd1 vssd1 vccd1 vccd1 _13758_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_168 _13641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16546_ _14787_/X _16521_/X _16529_/X _14724_/X _16545_/X vssd1 vssd1 vccd1 vccd1
+ _16546_/X sky130_fd_sc_hd__a311o_1
XFILLER_250_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_179 _19882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ _25590_/Q vssd1 vssd1 vccd1 vccd1 _19774_/A sky130_fd_sc_hd__buf_6
X_19265_ _25558_/Q _18459_/X _19264_/X _18436_/A _18466_/X vssd1 vssd1 vccd1 vccd1
+ _19265_/X sky130_fd_sc_hd__a221o_1
XFILLER_31_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13689_ _13689_/A _17819_/B vssd1 vssd1 vccd1 vccd1 _13690_/B sky130_fd_sc_hd__nor2_1
X_16477_ _26811_/Q _26455_/Q _16500_/S vssd1 vssd1 vccd1 vccd1 _16477_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18216_ _14562_/X _17997_/A _18215_/Y _16706_/A vssd1 vssd1 vccd1 vccd1 _18216_/X
+ sky130_fd_sc_hd__a22o_1
X_15428_ _13255_/X _26864_/Q _25778_/Q _16347_/S _15424_/A vssd1 vssd1 vccd1 vccd1
+ _15428_/X sky130_fd_sc_hd__a221o_1
XFILLER_176_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19196_ _19196_/A vssd1 vssd1 vccd1 vccd1 _19196_/X sky130_fd_sc_hd__clkbuf_2
X_15359_ _25817_/Q _16240_/S _15265_/X _15358_/X vssd1 vssd1 vccd1 vccd1 _15359_/X
+ sky130_fd_sc_hd__o211a_1
X_18147_ _18147_/A vssd1 vssd1 vccd1 vccd1 _25599_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18078_ _18078_/A vssd1 vssd1 vccd1 vccd1 _18603_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17029_ _17028_/X _16885_/B _17025_/X input221/X vssd1 vssd1 vccd1 vccd1 _17029_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_116_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20040_ _20007_/A _20038_/X _20039_/X vssd1 vssd1 vccd1 vccd1 _20040_/X sky130_fd_sc_hd__a21o_1
XFILLER_259_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21991_ _21991_/A vssd1 vssd1 vccd1 vccd1 _26108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23730_ _23730_/A vssd1 vssd1 vccd1 vccd1 _26761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ _23757_/A vssd1 vssd1 vccd1 vccd1 _20942_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_254_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23661_ _26737_/Q _23578_/X _23667_/S vssd1 vssd1 vccd1 vccd1 _23662_/A sky130_fd_sc_hd__mux2_1
X_20873_ _25829_/Q _20866_/X _20885_/S vssd1 vssd1 vccd1 vccd1 _20874_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25400_ _23693_/X _27297_/Q _25404_/S vssd1 vssd1 vccd1 vccd1 _25401_/A sky130_fd_sc_hd__mux2_1
X_22612_ _26320_/Q _22618_/B vssd1 vssd1 vccd1 vccd1 _22612_/Y sky130_fd_sc_hd__nand2_1
XFILLER_242_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26380_ _26609_/CLK _26380_/D vssd1 vssd1 vccd1 vccd1 _26380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23592_ _26709_/Q _23590_/X _23604_/S vssd1 vssd1 vccd1 vccd1 _23593_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25331_ _25331_/A vssd1 vssd1 vccd1 vccd1 _27266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22543_ _26294_/Q _22551_/B vssd1 vssd1 vccd1 vccd1 _22543_/Y sky130_fd_sc_hd__nand2_1
XFILLER_194_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25262_ _25319_/S vssd1 vssd1 vccd1 vccd1 _25271_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_210_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22474_ _22474_/A _22480_/B vssd1 vssd1 vccd1 vccd1 _22475_/A sky130_fd_sc_hd__and2_1
X_27001_ _27001_/CLK _27001_/D vssd1 vssd1 vccd1 vccd1 _27001_/Q sky130_fd_sc_hd__dfxtp_1
X_24213_ _26961_/Q _26960_/Q _24213_/C vssd1 vssd1 vccd1 vccd1 _24215_/B sky130_fd_sc_hd__and3_1
XFILLER_148_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21425_ _21556_/A vssd1 vssd1 vccd1 vccd1 _21425_/X sky130_fd_sc_hd__buf_4
XFILLER_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25193_ _24671_/B _25189_/X _25187_/X _27206_/Q _25191_/X vssd1 vssd1 vccd1 vccd1
+ _27206_/D sky130_fd_sc_hd__o221a_1
XFILLER_147_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24144_ _26938_/Q _23606_/X _24146_/S vssd1 vssd1 vccd1 vccd1 _24145_/A sky130_fd_sc_hd__mux2_1
X_21356_ input105/X input77/X _21356_/S vssd1 vssd1 vccd1 vccd1 _21357_/A sky130_fd_sc_hd__mux2_8
XFILLER_151_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20307_ _20205_/B _20301_/Y _20306_/X vssd1 vssd1 vccd1 vccd1 _20352_/A sky130_fd_sc_hd__a21oi_2
XFILLER_135_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24075_ _24075_/A vssd1 vssd1 vccd1 vccd1 _26907_/D sky130_fd_sc_hd__clkbuf_1
X_21287_ _21346_/A vssd1 vssd1 vccd1 vccd1 _21641_/B sky130_fd_sc_hd__clkbuf_2
X_23026_ _26484_/Q _22733_/X _23028_/S vssd1 vssd1 vccd1 vccd1 _23027_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20238_ _27122_/Q _20707_/D vssd1 vssd1 vccd1 vccd1 _20238_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20169_ _20092_/A _19082_/X _20092_/B _20168_/X vssd1 vssd1 vccd1 vccd1 _20169_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _25589_/Q vssd1 vssd1 vccd1 vccd1 _13068_/A sky130_fd_sc_hd__inv_2
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24977_ _27160_/Q _24957_/X _24976_/Y vssd1 vssd1 vccd1 vccd1 _27160_/D sky130_fd_sc_hd__o21a_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26716_ _26878_/CLK _26716_/D vssd1 vssd1 vccd1 vccd1 _26716_/Q sky130_fd_sc_hd__dfxtp_1
X_14730_ _15227_/S vssd1 vssd1 vccd1 vccd1 _15095_/S sky130_fd_sc_hd__buf_2
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23928_ _23782_/X _26842_/Q _23930_/S vssd1 vssd1 vccd1 vccd1 _23929_/A sky130_fd_sc_hd__mux2_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _14661_/A vssd1 vssd1 vccd1 vccd1 _14662_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23859_ _23859_/A vssd1 vssd1 vccd1 vccd1 _26811_/D sky130_fd_sc_hd__clkbuf_1
X_26647_ _26903_/CLK _26647_/D vssd1 vssd1 vccd1 vccd1 _26647_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _13585_/X _26885_/Q _26757_/Q _13441_/S _15716_/S vssd1 vssd1 vccd1 vccd1
+ _13612_/X sky130_fd_sc_hd__a221o_1
X_16400_ _26807_/Q _26451_/Q _16400_/S vssd1 vssd1 vccd1 vccd1 _16400_/X sky130_fd_sc_hd__mux2_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ _17380_/A _17380_/B _17381_/B vssd1 vssd1 vccd1 vccd1 _25545_/D sky130_fd_sc_hd__nor3_1
X_14592_ _15071_/A vssd1 vssd1 vccd1 vccd1 _14593_/A sky130_fd_sc_hd__buf_2
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26578_ _27321_/CLK _26578_/D vssd1 vssd1 vccd1 vccd1 _26578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13543_ _13543_/A vssd1 vssd1 vccd1 vccd1 _14816_/A sky130_fd_sc_hd__buf_4
X_16331_ _16314_/X _16330_/X _15071_/A vssd1 vssd1 vccd1 vccd1 _16331_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_111_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25529_ _25553_/CLK _25529_/D vssd1 vssd1 vccd1 vccd1 _25529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16262_ _26511_/Q _26383_/Q _16262_/S vssd1 vssd1 vccd1 vccd1 _16262_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19050_ _16124_/Y _18371_/A _18368_/A _19048_/A _18307_/A vssd1 vssd1 vccd1 vccd1
+ _19050_/X sky130_fd_sc_hd__o221a_1
X_13474_ _15937_/S vssd1 vssd1 vccd1 vccd1 _15496_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_158_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15213_ _26804_/Q _26448_/Q _16441_/S vssd1 vssd1 vccd1 vccd1 _15213_/X sky130_fd_sc_hd__mux2_1
X_18001_ _18001_/A _18001_/B vssd1 vssd1 vccd1 vccd1 _18008_/A sky130_fd_sc_hd__or2_2
XFILLER_185_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16193_ _26085_/Q _25890_/Q _16193_/S vssd1 vssd1 vccd1 vccd1 _16193_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15144_ _15065_/X _26416_/Q _15142_/X _15143_/X vssd1 vssd1 vccd1 vccd1 _15144_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_275_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput309 _16744_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[13] sky130_fd_sc_hd__buf_2
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15075_ _25656_/Q _14609_/A _14613_/X vssd1 vssd1 vccd1 vccd1 _15075_/X sky130_fd_sc_hd__a21o_1
XFILLER_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19952_ _19951_/A _19951_/B _19951_/C vssd1 vssd1 vccd1 vccd1 _19952_/X sky130_fd_sc_hd__a21o_1
XFILLER_126_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14026_ input120/X input155/X _14132_/S vssd1 vssd1 vccd1 vccd1 _14026_/X sky130_fd_sc_hd__mux2_8
XFILLER_141_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18903_ _18903_/A _18903_/B vssd1 vssd1 vccd1 vccd1 _18903_/Y sky130_fd_sc_hd__nor2_1
XFILLER_268_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19883_ _20252_/B _18590_/X _19600_/X _19882_/Y vssd1 vssd1 vccd1 vccd1 _19883_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_268_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18834_ _18806_/X _18809_/X _18833_/X vssd1 vssd1 vccd1 vccd1 _18834_/X sky130_fd_sc_hd__a21o_4
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18765_ _18827_/A vssd1 vssd1 vccd1 vccd1 _18765_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_255_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15977_ _25841_/Q _26041_/Q _15980_/S vssd1 vssd1 vccd1 vccd1 _15977_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17716_ _18615_/A vssd1 vssd1 vccd1 vccd1 _18757_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_270_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14928_ _14920_/X _14927_/X _17179_/A vssd1 vssd1 vccd1 vccd1 _14928_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_270_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18696_ _19957_/A _19261_/B vssd1 vssd1 vccd1 vccd1 _18696_/X sky130_fd_sc_hd__or2_1
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17647_ _17650_/A _17647_/B vssd1 vssd1 vccd1 vccd1 _25594_/D sky130_fd_sc_hd__nor2_1
XFILLER_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14859_ _16401_/S vssd1 vssd1 vccd1 vccd1 _14859_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_91_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17578_ _25913_/Q _17568_/X _12937_/Y _17577_/X vssd1 vssd1 vccd1 vccd1 _17578_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19317_ _19317_/A _19317_/B vssd1 vssd1 vccd1 vccd1 _19317_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16529_ _14760_/X _16525_/X _16528_/X _20119_/A vssd1 vssd1 vccd1 vccd1 _16529_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_177_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19248_ _20683_/A _19246_/C _19246_/A vssd1 vssd1 vccd1 vccd1 _19249_/B sky130_fd_sc_hd__a21oi_1
XFILLER_164_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19179_ _25746_/Q _19179_/B vssd1 vssd1 vccd1 vccd1 _19180_/B sky130_fd_sc_hd__nor2_1
XFILLER_247_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21210_ _21219_/B _21210_/B vssd1 vssd1 vccd1 vccd1 _21866_/C sky130_fd_sc_hd__nor2_1
XFILLER_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22190_ _26180_/Q _22186_/X _22179_/X input279/X _22187_/X vssd1 vssd1 vccd1 vccd1
+ _22190_/X sky130_fd_sc_hd__a221o_1
XFILLER_172_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21141_ _21141_/A vssd1 vssd1 vccd1 vccd1 _25919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_198_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26931_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21072_ _25935_/Q _21075_/A _25934_/Q vssd1 vssd1 vccd1 vccd1 _21166_/A sky130_fd_sc_hd__a21oi_4
XFILLER_59_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_127_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27022_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_24900_ _24543_/B _24341_/A _24900_/C _24900_/D vssd1 vssd1 vccd1 vccd1 _24941_/A
+ sky130_fd_sc_hd__and4bb_2
X_20023_ _27146_/Q _27080_/Q vssd1 vssd1 vccd1 vccd1 _20023_/X sky130_fd_sc_hd__or2_1
X_25880_ _26599_/CLK _25880_/D vssd1 vssd1 vccd1 vccd1 _25880_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_258_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24831_ _20654_/A _24829_/X _24693_/Y _24830_/X vssd1 vssd1 vccd1 vccd1 _24831_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_101_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24762_ _24781_/A _24762_/B vssd1 vssd1 vccd1 vccd1 _25155_/A sky130_fd_sc_hd__nand2_4
X_21974_ _22031_/S vssd1 vssd1 vccd1 vccd1 _21983_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26501_ _27304_/CLK _26501_/D vssd1 vssd1 vccd1 vccd1 _26501_/Q sky130_fd_sc_hd__dfxtp_2
X_23713_ _23712_/X _26756_/Q _23716_/S vssd1 vssd1 vccd1 vccd1 _23714_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20925_ _20925_/A vssd1 vssd1 vccd1 vccd1 _25845_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24693_ _24703_/A _24693_/B vssd1 vssd1 vccd1 vccd1 _24693_/Y sky130_fd_sc_hd__nand2_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26432_ _26465_/CLK _26432_/D vssd1 vssd1 vccd1 vccd1 _26432_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_242_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23644_ _23644_/A vssd1 vssd1 vccd1 vccd1 _26729_/D sky130_fd_sc_hd__clkbuf_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20856_ _25824_/Q vssd1 vssd1 vccd1 vccd1 _20857_/A sky130_fd_sc_hd__clkbuf_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26363_ _26462_/CLK _26363_/D vssd1 vssd1 vccd1 vccd1 _26363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23575_ _23591_/A vssd1 vssd1 vccd1 vccd1 _23588_/S sky130_fd_sc_hd__buf_4
X_20787_ _20621_/X _25789_/Q _20787_/S vssd1 vssd1 vccd1 vccd1 _20788_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25314_ _25314_/A vssd1 vssd1 vccd1 vccd1 _27259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22526_ _22526_/A _22533_/B vssd1 vssd1 vccd1 vccd1 _22527_/A sky130_fd_sc_hd__and2_1
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26294_ _26297_/CLK _26294_/D vssd1 vssd1 vccd1 vccd1 _26294_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_211_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25245_ _25208_/A _19616_/X _24771_/A _24768_/B _25219_/A vssd1 vssd1 vccd1 vccd1
+ _25245_/X sky130_fd_sc_hd__a221o_1
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22457_ _26255_/Q _22457_/B vssd1 vssd1 vccd1 vccd1 _22457_/X sky130_fd_sc_hd__or2_1
XFILLER_194_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21408_ _21342_/X _21406_/X _21407_/X vssd1 vssd1 vccd1 vccd1 _21408_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_157_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13190_ _20868_/A _14452_/S vssd1 vssd1 vccd1 vccd1 _13190_/Y sky130_fd_sc_hd__xnor2_1
X_25176_ _25176_/A _25218_/A vssd1 vssd1 vccd1 vccd1 _25190_/A sky130_fd_sc_hd__nor2_1
XFILLER_124_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22388_ _22388_/A _22416_/C vssd1 vssd1 vccd1 vccd1 _22388_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24127_ _26930_/Q _23581_/X _24131_/S vssd1 vssd1 vccd1 vccd1 _24128_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21339_ _21271_/A _21338_/X _21259_/A vssd1 vssd1 vccd1 vccd1 _21339_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_150_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24058_ _24058_/A vssd1 vssd1 vccd1 vccd1 _26899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15900_ _13857_/A _15896_/X _15899_/X _13112_/A vssd1 vssd1 vccd1 vccd1 _15900_/X
+ sky130_fd_sc_hd__o211a_1
X_23009_ _26476_/Q _22707_/X _23017_/S vssd1 vssd1 vccd1 vccd1 _23010_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16880_ _16893_/A _16880_/B vssd1 vssd1 vccd1 vccd1 _16881_/A sky130_fd_sc_hd__and2_1
XFILLER_104_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831_ _13010_/A _15833_/A _15830_/Y _13756_/B vssd1 vssd1 vccd1 vccd1 _15831_/X
+ sky130_fd_sc_hd__o211a_2
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18550_ _18548_/X _18549_/X _16728_/B vssd1 vssd1 vccd1 vccd1 _18550_/X sky130_fd_sc_hd__a21o_1
X_15762_ _15491_/A _26343_/Q _26603_/Q _15501_/A _15939_/A vssd1 vssd1 vccd1 vccd1
+ _15762_/X sky130_fd_sc_hd__a221o_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ _14610_/B vssd1 vssd1 vccd1 vccd1 _14401_/B sky130_fd_sc_hd__inv_2
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17501_ _18077_/A _17772_/B vssd1 vssd1 vccd1 vccd1 _18036_/A sky130_fd_sc_hd__nand2_1
X_14713_ _14713_/A _14713_/B _14713_/C _14713_/D vssd1 vssd1 vccd1 vccd1 _15994_/A
+ sky130_fd_sc_hd__and4_2
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18481_ _17813_/B _18423_/B _17798_/X vssd1 vssd1 vccd1 vccd1 _18482_/B sky130_fd_sc_hd__a21bo_1
XFILLER_206_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _15301_/S _15691_/X _15692_/X _13367_/X vssd1 vssd1 vccd1 vccd1 _15694_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _24208_/A vssd1 vssd1 vccd1 vccd1 _24239_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_205_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14644_ _14692_/S vssd1 vssd1 vccd1 vccd1 _16467_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17363_ _17382_/A _17370_/C vssd1 vssd1 vccd1 vccd1 _17363_/Y sky130_fd_sc_hd__nor2_1
X_14575_ _14575_/A _17818_/B vssd1 vssd1 vccd1 vccd1 _18549_/S sky130_fd_sc_hd__and2_1
XFILLER_198_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19102_ _18383_/A _19100_/Y _18998_/A vssd1 vssd1 vccd1 vccd1 _19103_/C sky130_fd_sc_hd__o21a_1
XFILLER_9_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16314_ _14622_/A _16300_/X _16304_/X _16313_/X _14682_/A vssd1 vssd1 vccd1 vccd1
+ _16314_/X sky130_fd_sc_hd__a311o_1
X_13526_ _15488_/A _25768_/Q _15841_/S _26854_/Q _13834_/A vssd1 vssd1 vccd1 vccd1
+ _13526_/X sky130_fd_sc_hd__o221a_1
XFILLER_202_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17294_ _17332_/A _17294_/B _17296_/B vssd1 vssd1 vccd1 vccd1 _25518_/D sky130_fd_sc_hd__nor3_1
X_19033_ _18775_/X _19031_/Y _18382_/A vssd1 vssd1 vccd1 vccd1 _19033_/X sky130_fd_sc_hd__o21ba_1
XFILLER_158_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16245_ _15060_/S _16242_/X _16244_/X _15040_/X vssd1 vssd1 vccd1 vccd1 _16245_/X
+ sky130_fd_sc_hd__a211o_1
X_13457_ _14124_/B vssd1 vssd1 vccd1 vccd1 _13756_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_185_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13388_ input116/X input152/X _13741_/S vssd1 vssd1 vccd1 vccd1 _13389_/B sky130_fd_sc_hd__mux2_8
X_16176_ _26117_/Q _26018_/Q _16176_/S vssd1 vssd1 vccd1 vccd1 _16176_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15127_ _15127_/A vssd1 vssd1 vccd1 vccd1 _16282_/A sky130_fd_sc_hd__buf_6
XFILLER_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15058_ _16319_/S vssd1 vssd1 vccd1 vccd1 _16223_/S sky130_fd_sc_hd__clkbuf_4
X_19935_ _20000_/A _19935_/B _19935_/C vssd1 vssd1 vccd1 vccd1 _19935_/X sky130_fd_sc_hd__or3_1
XFILLER_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14009_ _26494_/Q _26366_/Q _14009_/S vssd1 vssd1 vccd1 vccd1 _14009_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19866_ _27140_/Q _27074_/Q _19841_/B vssd1 vssd1 vccd1 vccd1 _19866_/X sky130_fd_sc_hd__a21o_1
XFILLER_256_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18817_ _18817_/A vssd1 vssd1 vccd1 vccd1 _18817_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19797_ _20189_/B vssd1 vssd1 vccd1 vccd1 _20249_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18748_ _18812_/A vssd1 vssd1 vccd1 vccd1 _18748_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18679_ _19235_/B _19574_/B _18678_/X _18037_/X vssd1 vssd1 vccd1 vccd1 _18679_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20710_ _19657_/X _19606_/Y _19607_/X _24986_/B vssd1 vssd1 vccd1 vccd1 _20710_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_224_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21690_ _25984_/Q input196/X _21696_/S vssd1 vssd1 vccd1 vccd1 _21691_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20641_ _20641_/A _20643_/B vssd1 vssd1 vccd1 vccd1 _20641_/X sky130_fd_sc_hd__or2_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23360_ _23360_/A vssd1 vssd1 vccd1 vccd1 _26618_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20572_ _20571_/X _25711_/Q _20572_/S vssd1 vssd1 vccd1 vccd1 _20573_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22311_ _26215_/Q _22310_/X _22300_/X _26316_/Q _22301_/X vssd1 vssd1 vccd1 vccd1
+ _22311_/X sky130_fd_sc_hd__a221o_1
X_23291_ _23860_/A _23291_/B vssd1 vssd1 vccd1 vccd1 _23348_/A sky130_fd_sc_hd__or2_4
XFILLER_191_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25030_ _25159_/B vssd1 vssd1 vccd1 vccd1 _25030_/X sky130_fd_sc_hd__clkbuf_2
X_22242_ input188/X _22222_/X _22238_/X _26293_/Q _22241_/X vssd1 vssd1 vccd1 vccd1
+ _22242_/X sky130_fd_sc_hd__a221o_1
XFILLER_106_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22173_ _26174_/Q _22171_/X _22160_/X input273/X _22172_/X vssd1 vssd1 vccd1 vccd1
+ _22173_/X sky130_fd_sc_hd__a221o_1
XFILLER_274_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21124_ _25915_/Q _21112_/X _21113_/X input14/X vssd1 vssd1 vccd1 vccd1 _21125_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26981_ _27001_/CLK _26981_/D vssd1 vssd1 vccd1 vccd1 _26981_/Q sky130_fd_sc_hd__dfxtp_1
X_25932_ _27227_/CLK _25932_/D vssd1 vssd1 vccd1 vccd1 _25932_/Q sky130_fd_sc_hd__dfxtp_4
X_21055_ _25896_/Q _20958_/X _21059_/S vssd1 vssd1 vccd1 vccd1 _21056_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20006_ _20006_/A _20006_/B vssd1 vssd1 vccd1 vccd1 _20007_/A sky130_fd_sc_hd__and2_1
XFILLER_219_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25863_ _26063_/CLK _25863_/D vssd1 vssd1 vccd1 vccd1 _25863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24814_ _27109_/Q _24818_/B vssd1 vssd1 vccd1 vccd1 _24814_/Y sky130_fd_sc_hd__nand2_1
XFILLER_246_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25794_ _25796_/CLK _25794_/D vssd1 vssd1 vccd1 vccd1 _25794_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24745_ _24969_/A vssd1 vssd1 vccd1 vccd1 _24746_/B sky130_fd_sc_hd__inv_2
XFILLER_61_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21957_ _20617_/X _26094_/Q _21959_/S vssd1 vssd1 vccd1 vccd1 _21958_/A sky130_fd_sc_hd__mux2_1
XFILLER_265_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_95_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26520_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20908_ _25840_/Q _20907_/X _20917_/S vssd1 vssd1 vccd1 vccd1 _20909_/A sky130_fd_sc_hd__mux2_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24676_ _24720_/A vssd1 vssd1 vccd1 vccd1 _24676_/X sky130_fd_sc_hd__clkbuf_2
X_12690_ _17504_/B _12799_/A vssd1 vssd1 vccd1 vccd1 _18006_/B sky130_fd_sc_hd__nand2_1
X_21888_ _21888_/A _21888_/B _21888_/C vssd1 vssd1 vccd1 vccd1 _23788_/B sky130_fd_sc_hd__or3_4
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26938_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23627_ _23627_/A vssd1 vssd1 vccd1 vccd1 _26721_/D sky130_fd_sc_hd__clkbuf_1
X_26415_ _26611_/CLK _26415_/D vssd1 vssd1 vccd1 vccd1 _26415_/Q sky130_fd_sc_hd__dfxtp_2
X_20839_ _20839_/A vssd1 vssd1 vccd1 vccd1 _25815_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14360_ _25574_/Q _21195_/B vssd1 vssd1 vccd1 vccd1 _14360_/Y sky130_fd_sc_hd__nor2_1
XFILLER_211_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26346_ _27281_/CLK _26346_/D vssd1 vssd1 vccd1 vccd1 _26346_/Q sky130_fd_sc_hd__dfxtp_1
X_23558_ _23558_/A vssd1 vssd1 vccd1 vccd1 _23558_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_196_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13311_ _13311_/A vssd1 vssd1 vccd1 vccd1 _13543_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_210_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22509_ _22509_/A _22513_/B vssd1 vssd1 vccd1 vccd1 _22510_/A sky130_fd_sc_hd__and2_1
XFILLER_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 core_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_1
X_14291_ _13484_/A _14289_/X _14290_/X _13945_/X vssd1 vssd1 vccd1 vccd1 _14292_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26277_ _26278_/CLK _26277_/D vssd1 vssd1 vccd1 vccd1 _26277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23489_ _26675_/Q _23111_/X _23491_/S vssd1 vssd1 vccd1 vccd1 _23490_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16030_ _13466_/A _15959_/A _16029_/Y vssd1 vssd1 vccd1 vccd1 _19971_/A sky130_fd_sc_hd__o21a_4
X_13242_ _13291_/A vssd1 vssd1 vccd1 vccd1 _13242_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25228_ _25228_/A vssd1 vssd1 vccd1 vccd1 _25228_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13173_ _13173_/A vssd1 vssd1 vccd1 vccd1 _13174_/A sky130_fd_sc_hd__buf_4
X_25159_ _25159_/A _25159_/B vssd1 vssd1 vccd1 vccd1 _25159_/Y sky130_fd_sc_hd__nand2_1
XFILLER_151_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17981_ _17973_/A _18904_/A _18202_/A vssd1 vssd1 vccd1 vccd1 _17981_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_69_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19720_ _22476_/A _19638_/X _19719_/X _19566_/X vssd1 vssd1 vccd1 vccd1 _25663_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16932_ _16932_/A _16932_/B vssd1 vssd1 vccd1 vccd1 _16983_/C sky130_fd_sc_hd__nor2_1
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19651_ _20186_/A vssd1 vssd1 vccd1 vccd1 _19651_/X sky130_fd_sc_hd__buf_2
XFILLER_265_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16863_ _16836_/X _16860_/X _16862_/X _16842_/X vssd1 vssd1 vccd1 vccd1 _16864_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_238_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18602_ _18602_/A vssd1 vssd1 vccd1 vccd1 _18602_/X sky130_fd_sc_hd__clkbuf_2
X_15814_ _25843_/Q _26043_/Q _15816_/S vssd1 vssd1 vccd1 vccd1 _15814_/X sky130_fd_sc_hd__mux2_1
XFILLER_219_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19582_ _19581_/X _19582_/B _19582_/C vssd1 vssd1 vccd1 vccd1 _19583_/B sky130_fd_sc_hd__and3b_1
XFILLER_92_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16794_ _16962_/A _16794_/B vssd1 vssd1 vccd1 vccd1 _16794_/Y sky130_fd_sc_hd__nand2_1
XFILLER_281_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18533_ _17671_/X _18527_/X _18528_/Y _18532_/Y vssd1 vssd1 vccd1 vccd1 _18533_/X
+ sky130_fd_sc_hd__a31o_1
X_15745_ _13126_/A _15740_/X _15744_/X _13163_/A vssd1 vssd1 vccd1 vccd1 _15745_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12957_ _13197_/A _13002_/A vssd1 vssd1 vccd1 vccd1 _21887_/B sky130_fd_sc_hd__nand2_2
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18464_ _26947_/Q _18461_/X _18463_/X _26979_/Q vssd1 vssd1 vccd1 vccd1 _18464_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15676_ _15676_/A vssd1 vssd1 vccd1 vccd1 _15676_/X sky130_fd_sc_hd__buf_2
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _25598_/Q _12933_/B vssd1 vssd1 vccd1 vccd1 _13569_/C sky130_fd_sc_hd__or2_1
XFILLER_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _17418_/A _17418_/C _17414_/X vssd1 vssd1 vccd1 vccd1 _17415_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14627_ _16386_/S vssd1 vssd1 vccd1 vccd1 _14969_/S sky130_fd_sc_hd__clkbuf_2
X_18395_ _27106_/Q _18504_/A _18390_/X _18394_/X vssd1 vssd1 vccd1 vccd1 _18395_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_159_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17346_ _25534_/Q _17344_/B _17345_/Y vssd1 vssd1 vccd1 vccd1 _25534_/D sky130_fd_sc_hd__o21a_1
XFILLER_158_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14558_ _13304_/A _14535_/X _14542_/X _13508_/A _14557_/X vssd1 vssd1 vccd1 vccd1
+ _14558_/X sky130_fd_sc_hd__a311o_2
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13509_ _13509_/A vssd1 vssd1 vccd1 vccd1 _14722_/A sky130_fd_sc_hd__buf_8
X_17277_ _25513_/Q _17275_/B _17276_/Y vssd1 vssd1 vccd1 vccd1 _25513_/D sky130_fd_sc_hd__o21a_1
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14489_ _14489_/A _14489_/B vssd1 vssd1 vccd1 vccd1 _14489_/Y sky130_fd_sc_hd__nor2_1
X_19016_ _18371_/A _18368_/A _19016_/S vssd1 vssd1 vccd1 vccd1 _19016_/X sky130_fd_sc_hd__mux2_1
X_16228_ _16405_/A _16228_/B vssd1 vssd1 vccd1 vccd1 _16228_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16159_ _26541_/Q _26149_/Q _16161_/S vssd1 vssd1 vccd1 vccd1 _16160_/B sky130_fd_sc_hd__mux2_1
XFILLER_170_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19918_ _19918_/A _19918_/B vssd1 vssd1 vccd1 vccd1 _19919_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19849_ _19849_/A _19910_/A vssd1 vssd1 vccd1 vccd1 _19849_/X sky130_fd_sc_hd__or2_1
XFILLER_229_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22860_ _26410_/Q _22701_/X _22862_/S vssd1 vssd1 vccd1 vccd1 _22861_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21811_ _21811_/A vssd1 vssd1 vccd1 vccd1 _26035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22791_ _22802_/A vssd1 vssd1 vccd1 vccd1 _22800_/S sky130_fd_sc_hd__clkbuf_4
X_24530_ _26323_/Q _24473_/X _24474_/X input238/X _21885_/A vssd1 vssd1 vccd1 vccd1
+ _24530_/X sky130_fd_sc_hd__a221o_2
X_21742_ _21742_/A vssd1 vssd1 vccd1 vccd1 _26005_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24461_ _27021_/Q _24448_/X _24460_/Y _24442_/X vssd1 vssd1 vccd1 vccd1 _27021_/D
+ sky130_fd_sc_hd__o211a_1
X_21673_ _21673_/A vssd1 vssd1 vccd1 vccd1 _25976_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26200_ _26250_/CLK _26200_/D vssd1 vssd1 vccd1 vccd1 _26200_/Q sky130_fd_sc_hd__dfxtp_1
X_23412_ _23412_/A vssd1 vssd1 vccd1 vccd1 _26640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_269_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20624_ _20624_/A _20630_/B vssd1 vssd1 vccd1 vccd1 _20624_/X sky130_fd_sc_hd__or2_1
X_27180_ _27196_/CLK _27180_/D vssd1 vssd1 vccd1 vccd1 _27180_/Q sky130_fd_sc_hd__dfxtp_1
X_24392_ _24454_/A vssd1 vssd1 vccd1 vccd1 _24392_/X sky130_fd_sc_hd__buf_4
X_26131_ _26909_/CLK _26131_/D vssd1 vssd1 vccd1 vccd1 _26131_/Q sky130_fd_sc_hd__dfxtp_1
X_23343_ _23343_/A vssd1 vssd1 vccd1 vccd1 _26610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20555_ _20597_/A vssd1 vssd1 vccd1 vccd1 _20572_/S sky130_fd_sc_hd__buf_4
XFILLER_138_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26062_ _27137_/CLK _26062_/D vssd1 vssd1 vccd1 vccd1 _26062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23274_ _23274_/A vssd1 vssd1 vccd1 vccd1 _26579_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20486_ _22817_/B _23363_/A _25249_/A vssd1 vssd1 vccd1 vccd1 _24004_/A sky130_fd_sc_hd__nand3_4
XFILLER_285_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25013_ _27168_/Q _25000_/X _25012_/X vssd1 vssd1 vccd1 vccd1 _27168_/D sky130_fd_sc_hd__o21ba_1
X_22225_ _26190_/Q _22152_/A _22224_/X _22217_/X vssd1 vssd1 vccd1 vccd1 _26190_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_142_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27327_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_279_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22156_ _26169_/Q _22154_/X _22140_/X input263/X _22155_/X vssd1 vssd1 vccd1 vccd1
+ _22156_/X sky130_fd_sc_hd__a221o_1
XFILLER_106_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput470 _25752_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[28] sky130_fd_sc_hd__buf_2
XFILLER_133_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput481 _25733_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[9] sky130_fd_sc_hd__buf_2
X_21107_ _21118_/A _21107_/B vssd1 vssd1 vccd1 vccd1 _21108_/A sky130_fd_sc_hd__or2_1
XFILLER_78_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26964_ _26995_/CLK _26964_/D vssd1 vssd1 vccd1 vccd1 _26964_/Q sky130_fd_sc_hd__dfxtp_1
X_22087_ _22087_/A vssd1 vssd1 vccd1 vccd1 _26151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25915_ _27117_/CLK _25915_/D vssd1 vssd1 vccd1 vccd1 _25915_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21038_ _21038_/A vssd1 vssd1 vccd1 vccd1 _25888_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26895_ _27314_/CLK _26895_/D vssd1 vssd1 vccd1 vccd1 _26895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_274_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13860_ _27238_/Q _15808_/B vssd1 vssd1 vccd1 vccd1 _13860_/X sky130_fd_sc_hd__or2_1
X_25846_ _27330_/A _25846_/D vssd1 vssd1 vccd1 vccd1 _25846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_270_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12811_ _19076_/A _14443_/A vssd1 vssd1 vccd1 vccd1 _16594_/A sky130_fd_sc_hd__nand2_2
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_509 input280/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22989_ _26467_/Q _22679_/X _22995_/S vssd1 vssd1 vccd1 vccd1 _22990_/A sky130_fd_sc_hd__mux2_1
X_13791_ _13791_/A vssd1 vssd1 vccd1 vccd1 _16336_/A sky130_fd_sc_hd__clkbuf_8
X_25777_ _27282_/CLK _25777_/D vssd1 vssd1 vccd1 vccd1 _25777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ _19016_/S _15530_/B vssd1 vssd1 vccd1 vccd1 _19034_/A sky130_fd_sc_hd__nand2_4
X_12742_ _25586_/Q vssd1 vssd1 vccd1 vccd1 _14431_/A sky130_fd_sc_hd__buf_2
X_24728_ _24960_/A vssd1 vssd1 vccd1 vccd1 _24729_/B sky130_fd_sc_hd__clkinv_2
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12673_ _12673_/A vssd1 vssd1 vccd1 vccd1 _12674_/A sky130_fd_sc_hd__buf_12
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15461_ _15455_/X _15457_/X _15460_/X _15646_/A _14362_/A vssd1 vssd1 vccd1 vccd1
+ _15461_/X sky130_fd_sc_hd__o221a_1
XFILLER_179_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24659_ _24682_/A _24659_/B vssd1 vssd1 vccd1 vccd1 _24659_/Y sky130_fd_sc_hd__nand2_2
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17200_ _17200_/A _17200_/B vssd1 vssd1 vccd1 vccd1 _17201_/A sky130_fd_sc_hd__and2_1
X_14412_ _13562_/X _14410_/Y _14411_/X _13556_/A _14407_/X vssd1 vssd1 vccd1 vccd1
+ _14412_/X sky130_fd_sc_hd__o2111a_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18180_ _18910_/A _18178_/X _18381_/A vssd1 vssd1 vccd1 vccd1 _18181_/C sky130_fd_sc_hd__o21ba_1
X_15392_ _26672_/Q _25712_/Q _16436_/S vssd1 vssd1 vccd1 vccd1 _15392_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17131_ _17504_/C _17131_/B vssd1 vssd1 vccd1 vccd1 _17131_/Y sky130_fd_sc_hd__nand2_1
X_26329_ _27267_/CLK _26329_/D vssd1 vssd1 vccd1 vccd1 _26329_/Q sky130_fd_sc_hd__dfxtp_2
X_14343_ _13582_/A _26686_/Q _26814_/Q _13993_/A vssd1 vssd1 vccd1 vccd1 _14343_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14274_ _26655_/Q _14497_/A _13048_/A vssd1 vssd1 vccd1 vccd1 _14274_/X sky130_fd_sc_hd__o21a_1
X_17062_ _25971_/Q _17061_/X _16991_/X _17051_/X vssd1 vssd1 vccd1 vccd1 _17062_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16013_ _26792_/Q _26436_/Q _16013_/S vssd1 vssd1 vccd1 vccd1 _16013_/X sky130_fd_sc_hd__mux2_1
X_13225_ _14296_/S vssd1 vssd1 vccd1 vccd1 _15923_/S sky130_fd_sc_hd__buf_4
XFILLER_171_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13156_ _15468_/B vssd1 vssd1 vccd1 vccd1 _16061_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13087_ _14176_/S vssd1 vssd1 vccd1 vccd1 _15904_/S sky130_fd_sc_hd__clkbuf_8
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _17920_/X _17944_/X _17961_/X _18685_/S vssd1 vssd1 vccd1 vccd1 _17964_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19703_ _19704_/A _19704_/B vssd1 vssd1 vccd1 vccd1 _19703_/X sky130_fd_sc_hd__and2_1
X_16915_ _16915_/A vssd1 vssd1 vccd1 vccd1 _16915_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_239_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17895_ _17941_/A vssd1 vssd1 vccd1 vccd1 _18347_/S sky130_fd_sc_hd__buf_2
XFILLER_93_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19634_ _19640_/A _19634_/B _19634_/C vssd1 vssd1 vccd1 vccd1 _24641_/A sky130_fd_sc_hd__and3b_4
XFILLER_66_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16846_ _16846_/A _16859_/A vssd1 vssd1 vccd1 vccd1 _16847_/A sky130_fd_sc_hd__nand2_2
XFILLER_253_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19565_ _25660_/Q _19568_/B vssd1 vssd1 vccd1 vccd1 _19565_/X sky130_fd_sc_hd__or2_1
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16777_ _22524_/A _16769_/X _16770_/X _19256_/B vssd1 vssd1 vccd1 vccd1 _16777_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_281_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13989_ _15983_/S _13988_/X _12700_/A vssd1 vssd1 vccd1 vccd1 _13989_/X sky130_fd_sc_hd__o21a_1
X_18516_ _18952_/B vssd1 vssd1 vccd1 vccd1 _19261_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15728_ _15722_/X _15724_/X _15727_/X _15819_/S _13630_/X vssd1 vssd1 vccd1 vccd1
+ _15728_/X sky130_fd_sc_hd__o221a_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19496_ _19484_/X _18246_/X _19495_/X _19489_/X vssd1 vssd1 vccd1 vccd1 _25633_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18447_ _27075_/Q _18815_/A _18816_/A _27173_/Q _18817_/A vssd1 vssd1 vccd1 vccd1
+ _18447_/X sky130_fd_sc_hd__a221o_1
XFILLER_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15659_ _15659_/A _16889_/A vssd1 vssd1 vccd1 vccd1 _15659_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18378_ _25729_/Q vssd1 vssd1 vccd1 vccd1 _19772_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_187_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17329_ _17327_/X _17331_/C _17328_/Y vssd1 vssd1 vccd1 vccd1 _25529_/D sky130_fd_sc_hd__o21a_1
XFILLER_175_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20340_ _27158_/Q _27092_/Q vssd1 vssd1 vccd1 vccd1 _20342_/A sky130_fd_sc_hd__nand2_1
XFILLER_162_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20271_ _20240_/Y _20242_/Y _20268_/X _20269_/Y vssd1 vssd1 vccd1 vccd1 _20271_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_255_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22010_ _26117_/Q _20939_/X _22016_/S vssd1 vssd1 vccd1 vccd1 _22011_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput209 localMemory_wb_adr_i[5] vssd1 vssd1 vccd1 vccd1 input209/X sky130_fd_sc_hd__clkbuf_1
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23961_ _26856_/Q _23549_/X _23965_/S vssd1 vssd1 vccd1 vccd1 _23962_/A sky130_fd_sc_hd__mux2_1
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25700_ _27276_/CLK _25700_/D vssd1 vssd1 vccd1 vccd1 _25700_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_112_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22912_ _26433_/Q _22672_/X _22912_/S vssd1 vssd1 vccd1 vccd1 _22913_/A sky130_fd_sc_hd__mux2_1
X_23892_ _23892_/A vssd1 vssd1 vccd1 vccd1 _26825_/D sky130_fd_sc_hd__clkbuf_1
X_26680_ _26744_/CLK _26680_/D vssd1 vssd1 vccd1 vccd1 _26680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22843_ _26402_/Q _22675_/X _22851_/S vssd1 vssd1 vccd1 vccd1 _22844_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25631_ _26813_/CLK _25631_/D vssd1 vssd1 vccd1 vccd1 _25631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22774_ _26372_/Q _22682_/X _22778_/S vssd1 vssd1 vccd1 vccd1 _22775_/A sky130_fd_sc_hd__mux2_1
X_25562_ _27000_/CLK _25562_/D vssd1 vssd1 vccd1 vccd1 _25562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27301_ _27301_/CLK _27301_/D vssd1 vssd1 vccd1 vccd1 _27301_/Q sky130_fd_sc_hd__dfxtp_1
X_21725_ _21725_/A vssd1 vssd1 vccd1 vccd1 _25997_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24513_ _24518_/A _24974_/A vssd1 vssd1 vccd1 vccd1 _24513_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25493_ _27327_/CLK _25493_/D vssd1 vssd1 vccd1 vccd1 _25493_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27232_ _27295_/CLK _27232_/D vssd1 vssd1 vccd1 vccd1 _27232_/Q sky130_fd_sc_hd__dfxtp_1
X_24444_ _26307_/Q _24473_/A _24474_/A input220/X _24395_/X vssd1 vssd1 vccd1 vccd1
+ _24444_/X sky130_fd_sc_hd__a221o_1
X_21656_ _25969_/Q input190/X _21662_/S vssd1 vssd1 vccd1 vccd1 _21657_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20607_ _20607_/A vssd1 vssd1 vccd1 vccd1 _25719_/D sky130_fd_sc_hd__clkbuf_1
X_24375_ _24494_/A vssd1 vssd1 vccd1 vccd1 _24408_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_27163_ _27164_/CLK _27163_/D vssd1 vssd1 vccd1 vccd1 _27163_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21587_ _21587_/A vssd1 vssd1 vccd1 vccd1 _21587_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26114_ _26531_/CLK _26114_/D vssd1 vssd1 vccd1 vccd1 _26114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23326_ _23348_/A vssd1 vssd1 vccd1 vccd1 _23335_/S sky130_fd_sc_hd__buf_4
X_20538_ _23722_/A vssd1 vssd1 vccd1 vccd1 _20538_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_181_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27094_ _27176_/CLK _27094_/D vssd1 vssd1 vccd1 vccd1 _27094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23257_ _23268_/A vssd1 vssd1 vccd1 vccd1 _23266_/S sky130_fd_sc_hd__clkbuf_4
X_26045_ _26796_/CLK _26045_/D vssd1 vssd1 vccd1 vccd1 _26045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20469_ _20703_/A _20355_/X _20468_/X _20357_/X vssd1 vssd1 vccd1 vccd1 _20470_/B
+ sky130_fd_sc_hd__o22a_1
X_13010_ _13010_/A vssd1 vssd1 vccd1 vccd1 _13011_/A sky130_fd_sc_hd__buf_2
XFILLER_134_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22208_ _26185_/Q _22201_/X _22206_/X _22207_/X _22203_/X vssd1 vssd1 vccd1 vccd1
+ _22208_/X sky130_fd_sc_hd__a221o_1
XFILLER_152_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23188_ _26541_/Q _23105_/X _23194_/S vssd1 vssd1 vccd1 vccd1 _23189_/A sky130_fd_sc_hd__mux2_1
XFILLER_279_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22139_ _26165_/Q _22136_/X _22138_/X _22132_/X vssd1 vssd1 vccd1 vccd1 _26165_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_267_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26947_ _26980_/CLK _26947_/D vssd1 vssd1 vccd1 vccd1 _26947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14961_ _12776_/A _26420_/Q _14948_/S _14960_/X vssd1 vssd1 vccd1 vccd1 _14961_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16700_ _16951_/A vssd1 vssd1 vccd1 vccd1 _16864_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13912_ _14403_/A vssd1 vssd1 vccd1 vccd1 _14489_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17680_ _20487_/A _18094_/A vssd1 vssd1 vccd1 vccd1 _17681_/A sky130_fd_sc_hd__nor2_4
X_26878_ _26878_/CLK _26878_/D vssd1 vssd1 vccd1 vccd1 _26878_/Q sky130_fd_sc_hd__dfxtp_1
X_14892_ _15005_/S vssd1 vssd1 vccd1 vccd1 _14984_/S sky130_fd_sc_hd__buf_2
XFILLER_235_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16631_ _16631_/A _18838_/B vssd1 vssd1 vccd1 vccd1 _16635_/C sky130_fd_sc_hd__xnor2_4
XFILLER_75_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25829_ _26240_/CLK _25829_/D vssd1 vssd1 vccd1 vccd1 _25829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13843_ _16015_/A _13843_/B vssd1 vssd1 vccd1 vccd1 _13843_/X sky130_fd_sc_hd__or2_1
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_262_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_306 _25912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_317 _19620_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19350_ _18144_/A _16566_/A _19349_/X vssd1 vssd1 vccd1 vccd1 _19350_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_328 _19616_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16562_ _16562_/A _19356_/A vssd1 vssd1 vccd1 vccd1 _19385_/B sky130_fd_sc_hd__xnor2_4
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13774_ _13966_/A vssd1 vssd1 vccd1 vccd1 _13775_/A sky130_fd_sc_hd__buf_2
XINSDIODE2_339 _19609_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18301_ _25505_/Q _18810_/A _18298_/X _18300_/X _18832_/A vssd1 vssd1 vccd1 vccd1
+ _18301_/X sky130_fd_sc_hd__o221a_1
XFILLER_43_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15513_ _13347_/A _15511_/X _15512_/X _14228_/X vssd1 vssd1 vccd1 vccd1 _15513_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19281_ _25749_/Q vssd1 vssd1 vccd1 vccd1 _19283_/A sky130_fd_sc_hd__buf_8
X_12725_ _25577_/Q vssd1 vssd1 vccd1 vccd1 _17992_/A sky130_fd_sc_hd__buf_4
XFILLER_231_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16493_ _26875_/Q _25789_/Q _16493_/S vssd1 vssd1 vccd1 vccd1 _16493_/X sky130_fd_sc_hd__mux2_1
XFILLER_231_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18232_ _18232_/A vssd1 vssd1 vccd1 vccd1 _18812_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15444_ _14599_/A _15442_/Y _15443_/X _14612_/A vssd1 vssd1 vccd1 vccd1 _15444_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_176_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18163_ _18160_/X _18162_/X _18238_/A vssd1 vssd1 vccd1 vccd1 _18163_/X sky130_fd_sc_hd__a21o_1
X_15375_ _15167_/A _26704_/Q _26832_/Q _16163_/S vssd1 vssd1 vccd1 vccd1 _15375_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17114_ _17224_/B vssd1 vssd1 vccd1 vccd1 _17114_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14326_ _25632_/Q _13933_/A _13577_/A _25600_/Q vssd1 vssd1 vccd1 vccd1 _14326_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_128_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18094_ _18094_/A vssd1 vssd1 vccd1 vccd1 _18805_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17045_ _17042_/X _16965_/B _16965_/C _17013_/X input234/X vssd1 vssd1 vccd1 vccd1
+ _17045_/X sky130_fd_sc_hd__a32o_4
X_14257_ _14257_/A vssd1 vssd1 vccd1 vccd1 _15989_/S sky130_fd_sc_hd__buf_4
XFILLER_172_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13208_ _13309_/A vssd1 vssd1 vccd1 vccd1 _18028_/A sky130_fd_sc_hd__buf_4
XFILLER_152_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14188_ _14188_/A vssd1 vssd1 vccd1 vccd1 _19455_/B sky130_fd_sc_hd__buf_2
XFILLER_135_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13139_ _13139_/A vssd1 vssd1 vccd1 vccd1 _13140_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ _20120_/A _19442_/B vssd1 vssd1 vccd1 vccd1 _18996_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ _17824_/B _15438_/B _17947_/S vssd1 vssd1 vccd1 vccd1 _17947_/X sky130_fd_sc_hd__mux2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17878_ _17875_/X _17876_/X _17958_/S vssd1 vssd1 vccd1 vccd1 _17878_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19617_ _27058_/Q _19617_/B _19617_/C vssd1 vssd1 vccd1 vccd1 _19617_/X sky130_fd_sc_hd__and3_1
X_16829_ _16829_/A vssd1 vssd1 vccd1 vccd1 _16829_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_226_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19548_ _19538_/X _19207_/X _19547_/X _19541_/X vssd1 vssd1 vccd1 vccd1 _25653_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19479_ _18144_/A _25166_/A _19478_/X vssd1 vssd1 vccd1 vccd1 _19479_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21510_ _21587_/A vssd1 vssd1 vccd1 vccd1 _21510_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22490_ _22490_/A vssd1 vssd1 vccd1 vccd1 _26270_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21441_ _21436_/Y _21440_/X _21425_/X vssd1 vssd1 vccd1 vccd1 _21441_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24160_ _26944_/Q _26943_/Q _24160_/C vssd1 vssd1 vccd1 vccd1 _24163_/B sky130_fd_sc_hd__and3_1
XFILLER_163_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21372_ _21646_/S vssd1 vssd1 vccd1 vccd1 _21422_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_147_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23111_ _23584_/A vssd1 vssd1 vccd1 vccd1 _23111_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20323_ _27157_/Q _20323_/B vssd1 vssd1 vccd1 vccd1 _20323_/Y sky130_fd_sc_hd__nand2_1
X_24091_ _24091_/A vssd1 vssd1 vccd1 vccd1 _26913_/D sky130_fd_sc_hd__clkbuf_1
X_23042_ _26489_/Q _23041_/X _23051_/S vssd1 vssd1 vccd1 vccd1 _23043_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20254_ _20681_/A _19727_/X _20253_/X _19920_/A vssd1 vssd1 vccd1 vccd1 _20303_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20185_ _27152_/Q _20184_/Y _20371_/S vssd1 vssd1 vccd1 vccd1 _20185_/X sky130_fd_sc_hd__mux2_2
XFILLER_276_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26801_ _27316_/CLK _26801_/D vssd1 vssd1 vccd1 vccd1 _26801_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24993_ _27166_/Q _24986_/Y _24992_/X _24970_/X vssd1 vssd1 vccd1 vccd1 _27165_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26732_ _27314_/CLK _26732_/D vssd1 vssd1 vccd1 vccd1 _26732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_285_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23944_ _23944_/A vssd1 vssd1 vccd1 vccd1 _26848_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26663_ _27330_/A _26663_/D vssd1 vssd1 vccd1 vccd1 _26663_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23875_ _23875_/A vssd1 vssd1 vccd1 vccd1 _26817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25614_ _25660_/CLK _25614_/D vssd1 vssd1 vccd1 vccd1 _25614_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22826_ _22826_/A vssd1 vssd1 vccd1 vccd1 _26394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26594_ _26594_/CLK _26594_/D vssd1 vssd1 vccd1 vccd1 _26594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25545_ _25545_/CLK _25545_/D vssd1 vssd1 vccd1 vccd1 _25545_/Q sky130_fd_sc_hd__dfxtp_1
X_22757_ _22757_/A vssd1 vssd1 vccd1 vccd1 _26364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21708_ _21708_/A vssd1 vssd1 vccd1 vccd1 _25992_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13490_ _14307_/S vssd1 vssd1 vccd1 vccd1 _15759_/S sky130_fd_sc_hd__clkbuf_4
X_22688_ _23731_/A vssd1 vssd1 vccd1 vccd1 _22688_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_212_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25476_ _26843_/CLK _25476_/D vssd1 vssd1 vccd1 vccd1 _25476_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_200_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27215_ _27221_/CLK _27215_/D vssd1 vssd1 vccd1 vccd1 _27215_/Q sky130_fd_sc_hd__dfxtp_1
X_21639_ _25966_/Q _21273_/A _21638_/Y _21597_/X vssd1 vssd1 vccd1 vccd1 _25966_/D
+ sky130_fd_sc_hd__a211o_1
X_24427_ _26304_/Q _24393_/X _24394_/X input217/X _24395_/X vssd1 vssd1 vccd1 vccd1
+ _24427_/X sky130_fd_sc_hd__a221o_1
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27146_ _27160_/CLK _27146_/D vssd1 vssd1 vccd1 vccd1 _27146_/Q sky130_fd_sc_hd__dfxtp_4
X_15160_ _25893_/Q _16243_/B vssd1 vssd1 vccd1 vccd1 _15160_/X sky130_fd_sc_hd__or2_1
XFILLER_5_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24358_ _24390_/A vssd1 vssd1 vccd1 vccd1 _24372_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_165_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14111_ _14111_/A vssd1 vssd1 vccd1 vccd1 _14111_/X sky130_fd_sc_hd__buf_2
XFILLER_158_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23309_ _20521_/X _26595_/Q _23313_/S vssd1 vssd1 vccd1 vccd1 _23310_/A sky130_fd_sc_hd__mux2_1
X_15091_ _15422_/S vssd1 vssd1 vccd1 vccd1 _16441_/S sky130_fd_sc_hd__buf_4
X_24289_ _26987_/Q _24293_/C _24271_/X vssd1 vssd1 vccd1 vccd1 _24289_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_153_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27077_ _27176_/CLK _27077_/D vssd1 vssd1 vccd1 vccd1 _27077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14042_ _25874_/Q _14449_/B vssd1 vssd1 vccd1 vccd1 _14042_/X sky130_fd_sc_hd__or2_1
X_26028_ _26843_/CLK _26028_/D vssd1 vssd1 vccd1 vccd1 _26028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18850_ _25611_/Q _18719_/X _18849_/X _18790_/X vssd1 vssd1 vccd1 vccd1 _25611_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17801_ _14127_/B _17801_/B vssd1 vssd1 vccd1 vccd1 _17802_/B sky130_fd_sc_hd__and2b_1
XFILLER_268_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18781_ _25736_/Q _18781_/B vssd1 vssd1 vccd1 vccd1 _18781_/X sky130_fd_sc_hd__xor2_4
XTAP_5740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15993_ _15976_/X _15992_/X _13174_/A vssd1 vssd1 vccd1 vccd1 _15994_/B sky130_fd_sc_hd__a21oi_4
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17732_ _17732_/A _17732_/B vssd1 vssd1 vccd1 vccd1 _18465_/A sky130_fd_sc_hd__and2_1
XTAP_5773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14944_ _12751_/A _14942_/X _14943_/X vssd1 vssd1 vccd1 vccd1 _14944_/X sky130_fd_sc_hd__o21a_1
XTAP_5784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17663_ _19583_/A _18182_/B vssd1 vssd1 vccd1 vccd1 _19769_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14875_ _26809_/Q _26453_/Q _14878_/S vssd1 vssd1 vccd1 vccd1 _14875_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19402_ _27034_/Q _19063_/X _19401_/X _18759_/X vssd1 vssd1 vccd1 vccd1 _19402_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_103 _21504_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16614_ _16621_/B _16614_/B vssd1 vssd1 vccd1 vccd1 _19034_/B sky130_fd_sc_hd__or2_4
X_13826_ _13822_/X _13825_/X _13313_/A vssd1 vssd1 vccd1 vccd1 _13826_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_63_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_114 _22815_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17594_ _16513_/X _17551_/X _17553_/X _17593_/Y vssd1 vssd1 vccd1 vccd1 _17595_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_63_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_125 _23645_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_136 _12937_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_147 _13304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19333_ _27128_/Q _19056_/X _19331_/X _19332_/X vssd1 vssd1 vccd1 vccd1 _19333_/X
+ sky130_fd_sc_hd__o22a_2
X_16545_ _16537_/X _16544_/X _17179_/A vssd1 vssd1 vccd1 vccd1 _16545_/X sky130_fd_sc_hd__o21a_1
XINSDIODE2_158 _14725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13757_ _15482_/A _16839_/A _13756_/X _15526_/S vssd1 vssd1 vccd1 vccd1 _14575_/A
+ sky130_fd_sc_hd__o211a_1
XINSDIODE2_169 _14449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19264_ _26966_/Q _18461_/X _18463_/X _26998_/Q vssd1 vssd1 vccd1 vccd1 _19264_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12708_ _19798_/A vssd1 vssd1 vccd1 vccd1 _12721_/A sky130_fd_sc_hd__buf_6
X_16476_ _16472_/X _16475_/X _16476_/S vssd1 vssd1 vccd1 vccd1 _16476_/X sky130_fd_sc_hd__mux2_1
X_13688_ _13688_/A vssd1 vssd1 vccd1 vccd1 _17819_/B sky130_fd_sc_hd__clkbuf_2
X_18215_ _14562_/X _18213_/X _18548_/A vssd1 vssd1 vccd1 vccd1 _18215_/Y sky130_fd_sc_hd__o21ai_1
X_15427_ _13255_/X _26928_/Q _26412_/Q _16347_/S _15333_/A vssd1 vssd1 vccd1 vccd1
+ _15427_/X sky130_fd_sc_hd__a221o_1
XFILLER_176_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19195_ _18792_/X _19190_/X _19193_/X _19194_/X vssd1 vssd1 vccd1 vccd1 _19195_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_12_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18146_ _18336_/A _18146_/B vssd1 vssd1 vccd1 vccd1 _18147_/A sky130_fd_sc_hd__and2_1
X_15358_ _27251_/Q _16154_/B vssd1 vssd1 vccd1 vccd1 _15358_/X sky130_fd_sc_hd__or2_1
XFILLER_172_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14309_ _14307_/X _14308_/X _14309_/S vssd1 vssd1 vccd1 vccd1 _14309_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18077_ _18077_/A _18077_/B vssd1 vssd1 vccd1 vccd1 _18078_/A sky130_fd_sc_hd__or2_1
XFILLER_117_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15289_ _15071_/X _15250_/Y _15288_/Y _15830_/A vssd1 vssd1 vccd1 vccd1 _16927_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17028_ _17063_/A vssd1 vssd1 vccd1 vccd1 _17028_/X sky130_fd_sc_hd__buf_2
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ _19575_/A _16637_/C _19453_/S vssd1 vssd1 vccd1 vccd1 _18979_/X sky130_fd_sc_hd__mux2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21990_ _26108_/Q _20910_/X _21994_/S vssd1 vssd1 vccd1 vccd1 _21991_/A sky130_fd_sc_hd__mux2_1
X_20941_ _20941_/A vssd1 vssd1 vccd1 vccd1 _25850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_282_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20872_ _20971_/S vssd1 vssd1 vccd1 vccd1 _20885_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_226_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23660_ _23660_/A vssd1 vssd1 vccd1 vccd1 _26736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_281_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22611_ _22606_/X _22610_/Y _22600_/X vssd1 vssd1 vccd1 vccd1 _26319_/D sky130_fd_sc_hd__a21oi_1
XFILLER_81_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23591_ _23591_/A vssd1 vssd1 vccd1 vccd1 _23604_/S sky130_fd_sc_hd__buf_6
XFILLER_201_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25330_ _27266_/Q _23696_/A _25332_/S vssd1 vssd1 vccd1 vccd1 _25331_/A sky130_fd_sc_hd__mux2_1
X_22542_ _22538_/X _22541_/Y _24770_/A vssd1 vssd1 vccd1 vccd1 _26293_/D sky130_fd_sc_hd__a21oi_1
XFILLER_194_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25261_ _25261_/A vssd1 vssd1 vccd1 vccd1 _27235_/D sky130_fd_sc_hd__clkbuf_1
X_22473_ _22473_/A vssd1 vssd1 vccd1 vccd1 _26262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27000_ _27000_/CLK _27000_/D vssd1 vssd1 vccd1 vccd1 _27000_/Q sky130_fd_sc_hd__dfxtp_1
X_24212_ _26960_/Q _24213_/C _26961_/Q vssd1 vssd1 vccd1 vccd1 _24214_/B sky130_fd_sc_hd__a21oi_1
X_21424_ _21421_/X _25863_/Q _21423_/Y _21386_/X vssd1 vssd1 vccd1 vccd1 _21424_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_147_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25192_ _24668_/B _25189_/X _25187_/X _27205_/Q _25191_/X vssd1 vssd1 vccd1 vccd1
+ _27205_/D sky130_fd_sc_hd__o221a_1
XFILLER_277_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24143_ _24143_/A vssd1 vssd1 vccd1 vccd1 _26937_/D sky130_fd_sc_hd__clkbuf_1
X_21355_ _25863_/Q vssd1 vssd1 vccd1 vccd1 _21355_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_49_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27313_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20306_ _20206_/B _20302_/Y _20305_/X vssd1 vssd1 vccd1 vccd1 _20306_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24074_ _26907_/Q _23609_/X _24074_/S vssd1 vssd1 vccd1 vccd1 _24075_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21286_ _21286_/A vssd1 vssd1 vccd1 vccd1 _21286_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23025_ _23025_/A vssd1 vssd1 vccd1 vccd1 _26483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_277_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20237_ _19740_/X _20231_/X _20232_/Y _20235_/X _20707_/D vssd1 vssd1 vccd1 vccd1
+ _20237_/X sky130_fd_sc_hd__a311o_1
XFILLER_89_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20168_ _20168_/A _20194_/B vssd1 vssd1 vccd1 vccd1 _20168_/X sky130_fd_sc_hd__or2_1
XFILLER_89_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _12992_/A _25585_/Q vssd1 vssd1 vccd1 vccd1 _13590_/A sky130_fd_sc_hd__or2b_2
X_24976_ _24621_/A _24902_/A _24966_/X vssd1 vssd1 vccd1 vccd1 _24976_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20099_ _25675_/Q _20098_/C _22505_/A vssd1 vssd1 vccd1 vccd1 _20099_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_92_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26715_ _26715_/CLK _26715_/D vssd1 vssd1 vccd1 vccd1 _26715_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23927_ _23927_/A vssd1 vssd1 vccd1 vccd1 _26841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26646_ _27321_/CLK _26646_/D vssd1 vssd1 vccd1 vccd1 _26646_/Q sky130_fd_sc_hd__dfxtp_1
X_14660_ _14660_/A vssd1 vssd1 vccd1 vccd1 _14661_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23858_ _23785_/X _26811_/Q _23858_/S vssd1 vssd1 vccd1 vccd1 _23859_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13611_ _13611_/A vssd1 vssd1 vccd1 vccd1 _15716_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22809_ _26388_/Q _22733_/X _22811_/S vssd1 vssd1 vccd1 vccd1 _22810_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26577_ _27258_/CLK _26577_/D vssd1 vssd1 vccd1 vccd1 _26577_/Q sky130_fd_sc_hd__dfxtp_1
X_14591_ _14591_/A vssd1 vssd1 vccd1 vccd1 _15071_/A sky130_fd_sc_hd__buf_4
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23789_ _23845_/A vssd1 vssd1 vccd1 vccd1 _23858_/S sky130_fd_sc_hd__buf_6
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16330_ _12704_/A _16321_/X _16329_/X _14709_/A vssd1 vssd1 vccd1 vccd1 _16330_/X
+ sky130_fd_sc_hd__a211o_1
X_25528_ _25992_/CLK _25528_/D vssd1 vssd1 vccd1 vccd1 _25528_/Q sky130_fd_sc_hd__dfxtp_1
X_13542_ _13241_/A _13537_/X _13538_/X _15401_/A vssd1 vssd1 vccd1 vccd1 _13542_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_197_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16261_ _16259_/X _16260_/X _16261_/S vssd1 vssd1 vccd1 vccd1 _16261_/X sky130_fd_sc_hd__mux2_1
X_13473_ _15938_/S vssd1 vssd1 vccd1 vccd1 _15937_/S sky130_fd_sc_hd__clkbuf_4
X_25459_ _23779_/X _27324_/Q _25459_/S vssd1 vssd1 vccd1 vccd1 _25460_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18000_ _19358_/A _19454_/B _17989_/Y _19454_/A _17999_/X vssd1 vssd1 vccd1 vccd1
+ _18000_/X sky130_fd_sc_hd__o221a_1
X_15212_ _14764_/A _15209_/X _15211_/X vssd1 vssd1 vccd1 vccd1 _15212_/X sky130_fd_sc_hd__o21a_1
XFILLER_173_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16192_ _13242_/X _16189_/X _16191_/X _15333_/X vssd1 vssd1 vccd1 vccd1 _16192_/X
+ sky130_fd_sc_hd__a211o_1
X_15143_ _26932_/Q _16223_/S vssd1 vssd1 vccd1 vccd1 _15143_/X sky130_fd_sc_hd__or2_1
X_27129_ _27130_/CLK _27129_/D vssd1 vssd1 vccd1 vccd1 _27129_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_126_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15074_ _15074_/A _16409_/B vssd1 vssd1 vccd1 vccd1 _15074_/Y sky130_fd_sc_hd__nor2_1
X_19951_ _19951_/A _19951_/B _19951_/C vssd1 vssd1 vccd1 vccd1 _19951_/Y sky130_fd_sc_hd__nand3_1
XFILLER_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14025_ _14025_/A _14025_/B vssd1 vssd1 vccd1 vccd1 _14237_/C sky130_fd_sc_hd__or2_1
X_18902_ _18548_/X _18901_/X _15789_/B vssd1 vssd1 vccd1 vccd1 _18903_/B sky130_fd_sc_hd__a21oi_1
XFILLER_45_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19882_ _19882_/A _19882_/B vssd1 vssd1 vccd1 vccd1 _19882_/Y sky130_fd_sc_hd__nand2_1
XFILLER_150_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18833_ _17278_/X _18810_/X _18824_/X _18831_/X _18832_/X vssd1 vssd1 vccd1 vccd1
+ _18833_/X sky130_fd_sc_hd__o221a_1
XFILLER_150_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18764_ _18826_/A vssd1 vssd1 vccd1 vccd1 _18764_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_255_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15976_ _14713_/A _15963_/X _15967_/X _15975_/X _13876_/X vssd1 vssd1 vccd1 vccd1
+ _15976_/X sky130_fd_sc_hd__a311o_1
XFILLER_64_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17715_ _18161_/B vssd1 vssd1 vccd1 vccd1 _18615_/A sky130_fd_sc_hd__buf_2
X_14927_ _14804_/A _14923_/X _14926_/X _14818_/X vssd1 vssd1 vccd1 vccd1 _14927_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18695_ _27144_/Q vssd1 vssd1 vccd1 vccd1 _19957_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17646_ _19887_/A _17612_/X _17516_/X _17645_/Y vssd1 vssd1 vccd1 vccd1 _17647_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14858_ _16144_/S vssd1 vssd1 vccd1 vccd1 _16401_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_24_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13809_ _13827_/A vssd1 vssd1 vccd1 vccd1 _16015_/A sky130_fd_sc_hd__buf_2
XFILLER_205_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17577_ _25794_/Q vssd1 vssd1 vccd1 vccd1 _17577_/X sky130_fd_sc_hd__clkbuf_1
X_14789_ _14789_/A vssd1 vssd1 vccd1 vccd1 _16281_/S sky130_fd_sc_hd__buf_6
XFILLER_177_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19316_ _19087_/X _19313_/X _19315_/Y _18891_/X vssd1 vssd1 vccd1 vccd1 _19317_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16528_ _16517_/X _16526_/X _16527_/X _12758_/A vssd1 vssd1 vccd1 vccd1 _16528_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_189_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19247_ _25747_/Q vssd1 vssd1 vccd1 vccd1 _20683_/A sky130_fd_sc_hd__buf_8
X_16459_ _17851_/A _17850_/A vssd1 vssd1 vccd1 vccd1 _16561_/B sky130_fd_sc_hd__nor2_2
XFILLER_191_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19178_ _25746_/Q _19179_/B vssd1 vssd1 vccd1 vccd1 _19246_/C sky130_fd_sc_hd__and2_1
XFILLER_117_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18129_ _18465_/A vssd1 vssd1 vccd1 vccd1 _18572_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21140_ _21154_/A _21140_/B vssd1 vssd1 vccd1 vccd1 _21141_/A sky130_fd_sc_hd__or2_1
XFILLER_133_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21071_ input9/X vssd1 vssd1 vccd1 vccd1 _21075_/A sky130_fd_sc_hd__inv_2
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20022_ _27146_/Q _27080_/Q vssd1 vssd1 vccd1 vccd1 _20022_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24830_ _24874_/A vssd1 vssd1 vccd1 vccd1 _24830_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_167_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25690_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_67_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24761_ _24978_/A vssd1 vssd1 vccd1 vccd1 _24762_/B sky130_fd_sc_hd__clkinv_2
X_21973_ _21973_/A vssd1 vssd1 vccd1 vccd1 _26100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26500_ _26920_/CLK _26500_/D vssd1 vssd1 vccd1 vccd1 _26500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23712_ _23712_/A vssd1 vssd1 vccd1 vccd1 _23712_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20924_ _25845_/Q _20923_/X _20933_/S vssd1 vssd1 vccd1 vccd1 _20925_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24692_ _24699_/A _24692_/B vssd1 vssd1 vccd1 vccd1 _27080_/D sky130_fd_sc_hd__nor2_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26431_ _26433_/CLK _26431_/D vssd1 vssd1 vccd1 vccd1 _26431_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_270_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23643_ _26729_/Q _23552_/X _23645_/S vssd1 vssd1 vccd1 vccd1 _23644_/A sky130_fd_sc_hd__mux2_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20855_ _20855_/A vssd1 vssd1 vccd1 vccd1 _25823_/D sky130_fd_sc_hd__clkbuf_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26362_ _27266_/CLK _26362_/D vssd1 vssd1 vccd1 vccd1 _26362_/Q sky130_fd_sc_hd__dfxtp_2
X_23574_ _23574_/A vssd1 vssd1 vccd1 vccd1 _23574_/X sky130_fd_sc_hd__clkbuf_2
X_20786_ _20786_/A vssd1 vssd1 vccd1 vccd1 _25788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25313_ _23776_/X _27259_/Q _25315_/S vssd1 vssd1 vccd1 vccd1 _25314_/A sky130_fd_sc_hd__mux2_1
X_22525_ _22525_/A vssd1 vssd1 vccd1 vccd1 _26286_/D sky130_fd_sc_hd__clkbuf_1
X_26293_ _26297_/CLK _26293_/D vssd1 vssd1 vccd1 vccd1 _26293_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_211_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25244_ _27228_/Q _25225_/X _25228_/X _24765_/B _25243_/X vssd1 vssd1 vccd1 vccd1
+ _27228_/D sky130_fd_sc_hd__o221a_1
X_22456_ _26206_/Q _22446_/X _22454_/X _22455_/X vssd1 vssd1 vccd1 vccd1 _26254_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21407_ _21407_/A vssd1 vssd1 vccd1 vccd1 _21407_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22387_ _22387_/A _22387_/B vssd1 vssd1 vccd1 vccd1 _22416_/C sky130_fd_sc_hd__nor2_1
X_25175_ _25217_/A vssd1 vssd1 vccd1 vccd1 _25175_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21338_ input104/X input75/X _21356_/S vssd1 vssd1 vccd1 vccd1 _21338_/X sky130_fd_sc_hd__mux2_8
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24126_ _24126_/A vssd1 vssd1 vccd1 vccd1 _26929_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21269_ _21873_/A _17482_/B _21866_/B _21275_/A _21268_/X vssd1 vssd1 vccd1 vccd1
+ _21269_/X sky130_fd_sc_hd__a311o_1
XFILLER_151_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24057_ _26899_/Q _23584_/X _24059_/S vssd1 vssd1 vccd1 vccd1 _24058_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23008_ _23019_/A vssd1 vssd1 vccd1 vccd1 _23017_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_173_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ _15830_/A _15830_/B vssd1 vssd1 vccd1 vccd1 _15830_/Y sky130_fd_sc_hd__nor2_2
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15761_ _15486_/A _15758_/X _15760_/X _15311_/A vssd1 vssd1 vccd1 vccd1 _15761_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24959_ _27152_/Q _24957_/X _24958_/Y vssd1 vssd1 vccd1 vccd1 _27152_/D sky130_fd_sc_hd__o21a_1
X_12973_ _12973_/A _12973_/B _13916_/B vssd1 vssd1 vccd1 vccd1 _14610_/B sky130_fd_sc_hd__or3b_4
XFILLER_46_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _25568_/Q _17500_/B _18028_/B vssd1 vssd1 vccd1 vccd1 _17662_/B sky130_fd_sc_hd__nand3_4
XFILLER_246_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _14684_/X _14711_/X _14593_/X vssd1 vssd1 vccd1 vccd1 _14712_/Y sky130_fd_sc_hd__a21oi_2
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ _18480_/A vssd1 vssd1 vccd1 vccd1 _25604_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _14741_/A _26860_/Q _25774_/Q _16259_/S _13335_/A vssd1 vssd1 vccd1 vccd1
+ _15692_/X sky130_fd_sc_hd__a221o_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _25561_/Q _17434_/C _17430_/Y vssd1 vssd1 vccd1 vccd1 _25561_/D sky130_fd_sc_hd__o21a_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26629_ _27303_/CLK _26629_/D vssd1 vssd1 vccd1 vccd1 _26629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14643_ _14693_/S vssd1 vssd1 vccd1 vccd1 _16479_/A sky130_fd_sc_hd__buf_2
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17362_ _25540_/Q _17362_/B vssd1 vssd1 vccd1 vccd1 _17370_/C sky130_fd_sc_hd__and2_1
XFILLER_199_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14574_ _18482_/A _16723_/B _18498_/S vssd1 vssd1 vccd1 vccd1 _16729_/B sky130_fd_sc_hd__a21o_2
X_19101_ _18608_/X _19099_/X _19100_/Y vssd1 vssd1 vccd1 vccd1 _19103_/B sky130_fd_sc_hd__a21oi_1
XFILLER_203_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16313_ _15020_/A _16308_/X _16312_/X _14678_/A vssd1 vssd1 vccd1 vccd1 _16313_/X
+ sky130_fd_sc_hd__o211a_1
X_13525_ _13653_/S vssd1 vssd1 vccd1 vccd1 _13834_/A sky130_fd_sc_hd__clkbuf_4
X_17293_ _25517_/Q _25518_/Q _17293_/C vssd1 vssd1 vccd1 vccd1 _17296_/B sky130_fd_sc_hd__and3_1
XFILLER_158_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19032_ _18741_/X _19030_/X _19031_/Y vssd1 vssd1 vccd1 vccd1 _19032_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_185_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16244_ _26087_/Q _16301_/S _16308_/S _16243_/X vssd1 vssd1 vccd1 vccd1 _16244_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13456_ _18001_/A _16594_/A vssd1 vssd1 vccd1 vccd1 _14124_/B sky130_fd_sc_hd__nor2_4
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16175_ _26541_/Q _26149_/Q _16176_/S vssd1 vssd1 vccd1 vccd1 _16175_/X sky130_fd_sc_hd__mux2_1
X_13387_ _14834_/A _14834_/B _14323_/A vssd1 vssd1 vccd1 vccd1 _15074_/A sky130_fd_sc_hd__nor3_1
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15126_ _16350_/A _15103_/X _15125_/X vssd1 vssd1 vccd1 vccd1 _15126_/X sky130_fd_sc_hd__a21o_2
XFILLER_217_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15057_ _26806_/Q _26450_/Q _16242_/S vssd1 vssd1 vccd1 vccd1 _15057_/X sky130_fd_sc_hd__mux2_1
X_19934_ _19933_/A _19933_/B _19933_/C vssd1 vssd1 vccd1 vccd1 _19935_/C sky130_fd_sc_hd__a21oi_1
XFILLER_269_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14008_ _26334_/Q _26594_/Q _14008_/S vssd1 vssd1 vccd1 vccd1 _14008_/X sky130_fd_sc_hd__mux2_1
XFILLER_229_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19865_ _19870_/A _27075_/Q vssd1 vssd1 vccd1 vccd1 _19865_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18816_ _18816_/A vssd1 vssd1 vccd1 vccd1 _18816_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_283_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19796_ _19879_/A vssd1 vssd1 vccd1 vccd1 _19796_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18747_ _18811_/A vssd1 vssd1 vccd1 vccd1 _18747_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15959_ _15959_/A vssd1 vssd1 vccd1 vccd1 _23549_/A sky130_fd_sc_hd__buf_6
XFILLER_37_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18678_ _18678_/A _19290_/A vssd1 vssd1 vccd1 vccd1 _18678_/X sky130_fd_sc_hd__or2_1
XFILLER_252_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17629_ _16476_/S _17612_/X _17608_/X _17628_/Y vssd1 vssd1 vccd1 vccd1 _17630_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_211_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20640_ _26267_/Q _20633_/X _20639_/X _20631_/X vssd1 vssd1 vccd1 vccd1 _25730_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_211_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20571_ _23747_/A vssd1 vssd1 vccd1 vccd1 _20571_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22310_ _22310_/A vssd1 vssd1 vccd1 vccd1 _22310_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23290_ _23290_/A vssd1 vssd1 vccd1 vccd1 _26587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22241_ _22271_/A vssd1 vssd1 vccd1 vccd1 _22241_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22172_ _22203_/A vssd1 vssd1 vccd1 vccd1 _22172_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21123_ _21123_/A vssd1 vssd1 vccd1 vccd1 _25914_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26980_ _26980_/CLK _26980_/D vssd1 vssd1 vccd1 vccd1 _26980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25931_ _27221_/CLK _25931_/D vssd1 vssd1 vccd1 vccd1 _25931_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21054_ _21054_/A vssd1 vssd1 vccd1 vccd1 _25895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20005_ _22496_/A _19876_/X _19989_/X _20004_/Y _19874_/X vssd1 vssd1 vccd1 vccd1
+ _25672_/D sky130_fd_sc_hd__o221a_1
XFILLER_86_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25862_ _26063_/CLK _25862_/D vssd1 vssd1 vccd1 vccd1 _25862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24813_ _24809_/Y _24812_/X _24796_/X vssd1 vssd1 vccd1 vccd1 _27108_/D sky130_fd_sc_hd__a21oi_1
XFILLER_274_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_15_0_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_15_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_101_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25793_ _25796_/CLK _25793_/D vssd1 vssd1 vccd1 vccd1 _25793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24744_ _24744_/A vssd1 vssd1 vccd1 vccd1 _24744_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_227_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21956_ _21956_/A vssd1 vssd1 vccd1 vccd1 _26093_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _23722_/A vssd1 vssd1 vccd1 vccd1 _20907_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24675_ _24740_/A vssd1 vssd1 vccd1 vccd1 _24720_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_243_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21887_ _25249_/A _21887_/B vssd1 vssd1 vccd1 vccd1 _21888_/A sky130_fd_sc_hd__nor2_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26414_ _26610_/CLK _26414_/D vssd1 vssd1 vccd1 vccd1 _26414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23626_ _26721_/Q _23526_/X _23634_/S vssd1 vssd1 vccd1 vccd1 _23627_/A sky130_fd_sc_hd__mux2_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20838_ _25815_/Q vssd1 vssd1 vccd1 vccd1 _20839_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_70_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26345_ _27280_/CLK _26345_/D vssd1 vssd1 vccd1 vccd1 _26345_/Q sky130_fd_sc_hd__dfxtp_1
X_23557_ _23557_/A vssd1 vssd1 vccd1 vccd1 _26698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20769_ _20769_/A vssd1 vssd1 vccd1 vccd1 _25780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_64_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26920_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13310_ _13310_/A vssd1 vssd1 vccd1 vccd1 _13311_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_196_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22508_ _22508_/A vssd1 vssd1 vccd1 vccd1 _26278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14290_ _13252_/A _26687_/Q _26815_/Q _16020_/S _13943_/X vssd1 vssd1 vccd1 vccd1
+ _14290_/X sky130_fd_sc_hd__a221o_1
X_26276_ _26282_/CLK _26276_/D vssd1 vssd1 vccd1 vccd1 _26276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23488_ _23488_/A vssd1 vssd1 vccd1 vccd1 _26674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13241_ _13241_/A vssd1 vssd1 vccd1 vccd1 _13291_/A sky130_fd_sc_hd__buf_2
X_25227_ _27220_/Q _25225_/X _25207_/X _24732_/B _25226_/X vssd1 vssd1 vccd1 vccd1
+ _27220_/D sky130_fd_sc_hd__o221a_1
X_22439_ _26200_/Q _22432_/X _22438_/X _22428_/X vssd1 vssd1 vccd1 vccd1 _26248_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13172_ _13172_/A vssd1 vssd1 vccd1 vccd1 _13173_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_136_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25158_ _20699_/A _25138_/X _25157_/X vssd1 vssd1 vccd1 vccd1 _25158_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24109_ _26922_/Q _23555_/X _24109_/S vssd1 vssd1 vccd1 vccd1 _24110_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_272_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17980_ _17979_/Y _17971_/X _17978_/A _17219_/A vssd1 vssd1 vccd1 vccd1 _18904_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_124_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25089_ _20664_/A _25086_/X _25088_/X vssd1 vssd1 vccd1 vccd1 _25089_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_81_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16931_ _16931_/A vssd1 vssd1 vccd1 vccd1 _16931_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_266_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19650_ _19650_/A _20712_/B vssd1 vssd1 vccd1 vccd1 _20186_/A sky130_fd_sc_hd__and2_2
X_16862_ _16868_/A _16862_/B vssd1 vssd1 vccd1 vccd1 _16862_/X sky130_fd_sc_hd__or2_1
XFILLER_265_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15813_ _26794_/Q _26438_/Q _15825_/S vssd1 vssd1 vccd1 vccd1 _15813_/X sky130_fd_sc_hd__mux2_1
XFILLER_219_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18601_ _18362_/X _18415_/X _18364_/X vssd1 vssd1 vccd1 vccd1 _18601_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19581_ _19581_/A _19581_/B _19581_/C _19327_/X vssd1 vssd1 vccd1 vccd1 _19581_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_65_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16793_ _16785_/Y _16792_/X _16693_/X vssd1 vssd1 vccd1 vccd1 _16793_/X sky130_fd_sc_hd__a21o_1
XFILLER_281_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18532_ _18027_/A _18531_/X _18059_/A vssd1 vssd1 vccd1 vccd1 _18532_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_218_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15744_ _13065_/A _15741_/X _15743_/X _13142_/A vssd1 vssd1 vccd1 vccd1 _15744_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12956_ _12959_/A _25478_/Q vssd1 vssd1 vccd1 vccd1 _13002_/A sky130_fd_sc_hd__or2b_2
XFILLER_92_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _18463_/A vssd1 vssd1 vccd1 vccd1 _18463_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_233_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _15406_/A _26344_/Q _26604_/Q _15674_/X _15672_/A vssd1 vssd1 vccd1 vccd1
+ _15675_/X sky130_fd_sc_hd__a221o_1
XFILLER_18_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12887_ _15706_/B vssd1 vssd1 vccd1 vccd1 _14834_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17414_ _17414_/A vssd1 vssd1 vccd1 vccd1 _17414_/X sky130_fd_sc_hd__buf_4
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14626_ _15263_/S vssd1 vssd1 vccd1 vccd1 _16386_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18394_ _27074_/Q _18508_/A _18509_/A _27172_/Q _18510_/A vssd1 vssd1 vccd1 vccd1
+ _18394_/X sky130_fd_sc_hd__a221o_1
XFILLER_187_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _17382_/A _17351_/C vssd1 vssd1 vccd1 vccd1 _17345_/Y sky130_fd_sc_hd__nor2_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _14549_/X _14556_/X _13976_/A vssd1 vssd1 vccd1 vccd1 _14557_/X sky130_fd_sc_hd__o21a_1
XFILLER_187_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13508_ _13508_/A vssd1 vssd1 vccd1 vccd1 _13509_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17276_ _17285_/A _17282_/C vssd1 vssd1 vccd1 vccd1 _17276_/Y sky130_fd_sc_hd__nor2_1
X_14488_ input107/X input132/X _14488_/S vssd1 vssd1 vccd1 vccd1 _14489_/B sky130_fd_sc_hd__mux2_8
XFILLER_146_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19015_ _18362_/X _18798_/X _18799_/Y _18682_/A vssd1 vssd1 vccd1 vccd1 _19018_/C
+ sky130_fd_sc_hd__o211a_1
X_16227_ _12750_/A _16225_/X _16226_/X vssd1 vssd1 vccd1 vccd1 _16228_/B sky130_fd_sc_hd__o21ai_1
X_13439_ _13437_/X _13438_/X _13698_/A vssd1 vssd1 vccd1 vccd1 _13439_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16158_ _14694_/A _16153_/X _16157_/X _14706_/A vssd1 vssd1 vccd1 vccd1 _16167_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15109_ _15109_/A vssd1 vssd1 vccd1 vccd1 _15110_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16089_ _14791_/A _16086_/X _16088_/X _13291_/X vssd1 vssd1 vccd1 vccd1 _16093_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19917_ _19978_/A _19978_/B vssd1 vssd1 vccd1 vccd1 _19980_/C sky130_fd_sc_hd__xnor2_1
XFILLER_96_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19848_ _25732_/Q vssd1 vssd1 vccd1 vccd1 _20643_/A sky130_fd_sc_hd__buf_8
XFILLER_69_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19779_ _19779_/A vssd1 vssd1 vccd1 vccd1 _20015_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21810_ _26035_/Q _20891_/X _21816_/S vssd1 vssd1 vccd1 vccd1 _21811_/A sky130_fd_sc_hd__mux2_1
XFILLER_260_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22790_ _22790_/A vssd1 vssd1 vccd1 vccd1 _26379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21741_ _20525_/X _26005_/Q _21743_/S vssd1 vssd1 vccd1 vccd1 _21742_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24460_ _24464_/A _24948_/A vssd1 vssd1 vccd1 vccd1 _24460_/Y sky130_fd_sc_hd__nand2_1
XFILLER_269_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21672_ _25976_/Q input211/X _21674_/S vssd1 vssd1 vccd1 vccd1 _21673_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23411_ _26640_/Q _23101_/X _23419_/S vssd1 vssd1 vccd1 vccd1 _23412_/A sky130_fd_sc_hd__mux2_1
X_20623_ _20623_/A vssd1 vssd1 vccd1 vccd1 _25723_/D sky130_fd_sc_hd__clkbuf_1
X_24391_ _24506_/A vssd1 vssd1 vccd1 vccd1 _24391_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26130_ _26240_/CLK _26130_/D vssd1 vssd1 vccd1 vccd1 _26130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20554_ _23734_/A vssd1 vssd1 vccd1 vccd1 _20554_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23342_ _20584_/X _26610_/Q _23346_/S vssd1 vssd1 vccd1 vccd1 _23343_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26061_ _27164_/CLK _26061_/D vssd1 vssd1 vccd1 vccd1 _26061_/Q sky130_fd_sc_hd__dfxtp_1
X_20485_ _20485_/A vssd1 vssd1 vccd1 vccd1 _25249_/A sky130_fd_sc_hd__buf_4
X_23273_ _26579_/Q _23124_/X _23277_/S vssd1 vssd1 vccd1 vccd1 _23274_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25012_ _24645_/Y _25137_/A _25011_/Y _24773_/X vssd1 vssd1 vccd1 vccd1 _25012_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22224_ _26189_/Q _22222_/X _22206_/X _22223_/X _22155_/A vssd1 vssd1 vccd1 vccd1
+ _22224_/X sky130_fd_sc_hd__a221o_1
XFILLER_180_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22155_ _22155_/A vssd1 vssd1 vccd1 vccd1 _22155_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput460 _25743_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[19] sky130_fd_sc_hd__buf_2
XFILLER_279_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput471 _25753_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[29] sky130_fd_sc_hd__buf_2
X_21106_ _25910_/Q _21094_/X _21095_/X input40/X vssd1 vssd1 vccd1 vccd1 _21107_/B
+ sky130_fd_sc_hd__o22a_1
Xoutput482 _26940_/Q vssd1 vssd1 vccd1 vccd1 probe_state sky130_fd_sc_hd__buf_2
X_26963_ _26995_/CLK _26963_/D vssd1 vssd1 vccd1 vccd1 _26963_/Q sky130_fd_sc_hd__dfxtp_1
X_22086_ _26151_/Q _20945_/X _22088_/S vssd1 vssd1 vccd1 vccd1 _22087_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_182_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26580_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_154_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_111_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26974_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_25914_ _27117_/CLK _25914_/D vssd1 vssd1 vccd1 vccd1 _25914_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21037_ _25888_/Q _20932_/X _21037_/S vssd1 vssd1 vccd1 vccd1 _21038_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26894_ _26925_/CLK _26894_/D vssd1 vssd1 vccd1 vccd1 _26894_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_208_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25845_ _26796_/CLK _25845_/D vssd1 vssd1 vccd1 vccd1 _25845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_274_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12810_ _12810_/A _18076_/B _17133_/A _12810_/D vssd1 vssd1 vccd1 vccd1 _14443_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_216_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25776_ _27281_/CLK _25776_/D vssd1 vssd1 vccd1 vccd1 _25776_/Q sky130_fd_sc_hd__dfxtp_1
X_13790_ _13485_/X _13788_/X _13789_/X _12755_/A vssd1 vssd1 vccd1 vccd1 _13790_/X
+ sky130_fd_sc_hd__o211a_1
X_22988_ _22988_/A vssd1 vssd1 vccd1 vccd1 _26466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _25594_/Q vssd1 vssd1 vccd1 vccd1 _17443_/A sky130_fd_sc_hd__buf_4
X_24727_ _24742_/A _24727_/B vssd1 vssd1 vccd1 vccd1 _27088_/D sky130_fd_sc_hd__nor2_1
XFILLER_203_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21939_ _21939_/A vssd1 vssd1 vccd1 vccd1 _26085_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _15458_/X _15459_/X _15460_/S vssd1 vssd1 vccd1 vccd1 _15460_/X sky130_fd_sc_hd__mux2_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _25585_/Q vssd1 vssd1 vccd1 vccd1 _12673_/A sky130_fd_sc_hd__buf_2
X_24658_ _24749_/A vssd1 vssd1 vccd1 vccd1 _24682_/A sky130_fd_sc_hd__buf_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _14411_/A _15345_/A _13567_/B vssd1 vssd1 vccd1 vccd1 _14411_/X sky130_fd_sc_hd__or3b_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23609_ _23609_/A vssd1 vssd1 vccd1 vccd1 _23609_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15391_ _12674_/A _16368_/S _15244_/X _15390_/Y vssd1 vssd1 vccd1 vccd1 _17790_/A
+ sky130_fd_sc_hd__o22a_4
X_24589_ _24615_/A vssd1 vssd1 vccd1 vccd1 _24589_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_169_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17130_ _21300_/A _17114_/X hold4/X _17120_/X vssd1 vssd1 vccd1 vccd1 _25472_/D sky130_fd_sc_hd__o211a_1
X_26328_ _27266_/CLK _26328_/D vssd1 vssd1 vccd1 vccd1 _26328_/Q sky130_fd_sc_hd__dfxtp_2
X_14342_ _26622_/Q _26718_/Q _14344_/S vssd1 vssd1 vccd1 vccd1 _14342_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17061_ _17061_/A vssd1 vssd1 vccd1 vccd1 _17061_/X sky130_fd_sc_hd__clkbuf_2
X_26259_ _26974_/CLK _26259_/D vssd1 vssd1 vccd1 vccd1 _26259_/Q sky130_fd_sc_hd__dfxtp_1
X_14273_ _25695_/Q _14273_/B vssd1 vssd1 vccd1 vccd1 _14273_/X sky130_fd_sc_hd__or2_1
XFILLER_195_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16012_ _16000_/X _16003_/X _16011_/X vssd1 vssd1 vccd1 vccd1 _16012_/Y sky130_fd_sc_hd__o21ai_4
X_13224_ _14536_/S vssd1 vssd1 vccd1 vccd1 _14296_/S sky130_fd_sc_hd__buf_2
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13155_ _15453_/A vssd1 vssd1 vccd1 vccd1 _16067_/S sky130_fd_sc_hd__buf_4
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13086_ _13694_/A vssd1 vssd1 vccd1 vccd1 _13086_/X sky130_fd_sc_hd__clkbuf_2
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17963_ _18343_/A vssd1 vssd1 vccd1 vccd1 _18685_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_239_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19702_ _20630_/A _19698_/X _19701_/X _19604_/X vssd1 vssd1 vccd1 vccd1 _19704_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_16914_ _16924_/A _16914_/B vssd1 vssd1 vccd1 vccd1 _16915_/A sky130_fd_sc_hd__and2_1
XFILLER_266_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17894_ _17889_/X _17892_/X _18197_/S vssd1 vssd1 vccd1 vccd1 _17894_/X sky130_fd_sc_hd__mux2_1
XFILLER_254_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19633_ _19639_/A _19639_/B _19633_/C _19633_/D vssd1 vssd1 vccd1 vccd1 _19634_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_281_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16845_ _16845_/A vssd1 vssd1 vccd1 vccd1 _16845_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_225_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19564_ _19551_/X _19407_/X _19563_/X _19555_/X vssd1 vssd1 vccd1 vccd1 _25659_/D
+ sky130_fd_sc_hd__o211a_1
X_16776_ _16776_/A vssd1 vssd1 vccd1 vccd1 _19256_/B sky130_fd_sc_hd__buf_4
XFILLER_18_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13988_ _13986_/X _13987_/X _14246_/S vssd1 vssd1 vccd1 vccd1 _13988_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15727_ _15725_/X _15726_/X _15727_/S vssd1 vssd1 vccd1 vccd1 _15727_/X sky130_fd_sc_hd__mux2_1
X_18515_ _27140_/Q vssd1 vssd1 vccd1 vccd1 _19839_/A sky130_fd_sc_hd__clkbuf_4
X_12939_ _25913_/Q _12902_/A _12937_/Y _14404_/A vssd1 vssd1 vccd1 vccd1 _12940_/D
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19495_ _25633_/Q _19497_/B vssd1 vssd1 vccd1 vccd1 _19495_/X sky130_fd_sc_hd__or2_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18446_ _18813_/A vssd1 vssd1 vccd1 vccd1 _19364_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15658_ _15073_/A _23562_/A _15657_/X _15388_/A vssd1 vssd1 vccd1 vccd1 _16889_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14609_ _14609_/A vssd1 vssd1 vccd1 vccd1 _24351_/B sky130_fd_sc_hd__buf_2
XFILLER_21_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18377_ _18377_/A vssd1 vssd1 vccd1 vccd1 _18891_/A sky130_fd_sc_hd__clkbuf_2
X_15589_ _15589_/A vssd1 vssd1 vccd1 vccd1 _15676_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17328_ _17327_/X _17331_/C _17318_/X vssd1 vssd1 vccd1 vccd1 _17328_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17259_ _25508_/Q vssd1 vssd1 vccd1 vccd1 _17259_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_147_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20270_ _20268_/X _20269_/Y _20240_/Y _20242_/Y vssd1 vssd1 vccd1 vccd1 _20270_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23960_ _23960_/A vssd1 vssd1 vccd1 vccd1 _26855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22911_ _22911_/A vssd1 vssd1 vccd1 vccd1 _26432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_272_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23891_ _23728_/X _26825_/Q _23893_/S vssd1 vssd1 vccd1 vccd1 _23892_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25630_ _26813_/CLK _25630_/D vssd1 vssd1 vccd1 vccd1 _25630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22842_ _22888_/S vssd1 vssd1 vccd1 vccd1 _22851_/S sky130_fd_sc_hd__buf_2
XFILLER_84_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25561_ _27001_/CLK _25561_/D vssd1 vssd1 vccd1 vccd1 _25561_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_231_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22773_ _22773_/A vssd1 vssd1 vccd1 vccd1 _26371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27300_ _27301_/CLK _27300_/D vssd1 vssd1 vccd1 vccd1 _27300_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_25_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24512_ _24370_/S _25624_/Q _24511_/X vssd1 vssd1 vccd1 vccd1 _24974_/A sky130_fd_sc_hd__o21ai_4
XFILLER_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21724_ _20484_/X _25997_/Q _21732_/S vssd1 vssd1 vccd1 vccd1 _21725_/A sky130_fd_sc_hd__mux2_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25492_ _26683_/CLK _25492_/D vssd1 vssd1 vccd1 vccd1 _25492_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27231_ _27295_/CLK _27231_/D vssd1 vssd1 vccd1 vccd1 _27231_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24443_ _27018_/Q _24421_/X _24440_/Y _24442_/X vssd1 vssd1 vccd1 vccd1 _27018_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21655_ _21698_/A vssd1 vssd1 vccd1 vccd1 _21662_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27162_ _27164_/CLK _27162_/D vssd1 vssd1 vccd1 vccd1 _27162_/Q sky130_fd_sc_hd__dfxtp_1
X_20606_ _20605_/X _25719_/Q _20614_/S vssd1 vssd1 vccd1 vccd1 _20607_/A sky130_fd_sc_hd__mux2_1
X_24374_ _24390_/A vssd1 vssd1 vccd1 vccd1 _24494_/A sky130_fd_sc_hd__buf_2
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21586_ _21586_/A vssd1 vssd1 vccd1 vccd1 _21586_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26113_ _27280_/CLK _26113_/D vssd1 vssd1 vccd1 vccd1 _26113_/Q sky130_fd_sc_hd__dfxtp_1
X_23325_ _23325_/A vssd1 vssd1 vccd1 vccd1 _26602_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20537_ _23546_/A vssd1 vssd1 vccd1 vccd1 _23722_/A sky130_fd_sc_hd__buf_4
XFILLER_20_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27093_ _27093_/CLK _27093_/D vssd1 vssd1 vccd1 vccd1 _27093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26044_ _26531_/CLK _26044_/D vssd1 vssd1 vccd1 vccd1 _26044_/Q sky130_fd_sc_hd__dfxtp_1
X_20468_ _19472_/A _18019_/X _19477_/Y _20376_/Y vssd1 vssd1 vccd1 vccd1 _20468_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23256_ _23256_/A vssd1 vssd1 vccd1 vccd1 _26571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22207_ input3/X input269/X _22207_/S vssd1 vssd1 vccd1 vccd1 _22207_/X sky130_fd_sc_hd__mux2_1
X_20399_ _20399_/A _20399_/B _20379_/B vssd1 vssd1 vccd1 vccd1 _20400_/B sky130_fd_sc_hd__or3b_1
X_23187_ _23187_/A vssd1 vssd1 vccd1 vccd1 _26540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22138_ _26164_/Q _22122_/X _22124_/X input258/X _22137_/X vssd1 vssd1 vccd1 vccd1
+ _22138_/X sky130_fd_sc_hd__a221o_1
XFILLER_160_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput290 _17068_/X vssd1 vssd1 vccd1 vccd1 addr0[5] sky130_fd_sc_hd__buf_2
XFILLER_160_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26946_ _26980_/CLK _26946_/D vssd1 vssd1 vccd1 vccd1 _26946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14960_ _26936_/Q _14960_/B vssd1 vssd1 vccd1 vccd1 _14960_/X sky130_fd_sc_hd__or2_1
X_22069_ _26143_/Q _20919_/X _22077_/S vssd1 vssd1 vccd1 vccd1 _22070_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13911_ _13911_/A vssd1 vssd1 vccd1 vccd1 _13911_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26877_ _26877_/CLK _26877_/D vssd1 vssd1 vccd1 vccd1 _26877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14891_ _14891_/A vssd1 vssd1 vccd1 vccd1 _15005_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16630_ _18855_/A _18851_/B vssd1 vssd1 vccd1 vccd1 _16636_/C sky130_fd_sc_hd__xnor2_4
XFILLER_47_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13842_ _26527_/Q _26135_/Q _15775_/S vssd1 vssd1 vccd1 vccd1 _13843_/B sky130_fd_sc_hd__mux2_1
X_25828_ _26881_/CLK _25828_/D vssd1 vssd1 vccd1 vccd1 _25828_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16561_ _16561_/A _16561_/B vssd1 vssd1 vccd1 vccd1 _19356_/A sky130_fd_sc_hd__nor2_4
XFILLER_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_307 _25903_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_25759_ _26909_/CLK _25759_/D vssd1 vssd1 vccd1 vccd1 _25759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13773_ _13773_/A vssd1 vssd1 vccd1 vccd1 _13966_/A sky130_fd_sc_hd__buf_2
XINSDIODE2_318 _19620_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_329 _19616_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18300_ _25537_/Q _18825_/A _18299_/X _18829_/A _18830_/A vssd1 vssd1 vccd1 vccd1
+ _18300_/X sky130_fd_sc_hd__a221o_1
X_15512_ _15491_/X _26114_/Q _26015_/Q _15850_/S _15852_/A vssd1 vssd1 vccd1 vccd1
+ _15512_/X sky130_fd_sc_hd__a221o_1
XFILLER_71_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19280_ _19078_/X _19256_/Y _19271_/X _19279_/Y _18716_/X vssd1 vssd1 vccd1 vccd1
+ _19280_/X sky130_fd_sc_hd__a32o_1
X_12724_ _17669_/A vssd1 vssd1 vccd1 vccd1 _16591_/A sky130_fd_sc_hd__buf_4
X_16492_ _16499_/S _16489_/X _16491_/X _14650_/X vssd1 vssd1 vccd1 vccd1 _16492_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_203_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18231_ _25504_/Q _18807_/A _18808_/A _25536_/Q vssd1 vssd1 vccd1 vccd1 _18231_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15443_ _25648_/Q _15443_/B vssd1 vssd1 vccd1 vccd1 _15443_/X sky130_fd_sc_hd__and2_1
XFILLER_31_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18162_ _27103_/Q _18232_/A vssd1 vssd1 vccd1 vccd1 _18162_/X sky130_fd_sc_hd__or2_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15374_ _26640_/Q _26736_/Q _15374_/S vssd1 vssd1 vccd1 vccd1 _15374_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17113_ _17612_/A vssd1 vssd1 vccd1 vccd1 _17224_/B sky130_fd_sc_hd__buf_2
X_14325_ _14322_/X _14324_/X _14325_/S vssd1 vssd1 vccd1 vccd1 _14325_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18093_ _18927_/A vssd1 vssd1 vccd1 vccd1 _19078_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17044_ _17042_/X _16959_/B _16959_/C _17013_/X input233/X vssd1 vssd1 vccd1 vccd1
+ _17044_/X sky130_fd_sc_hd__a32o_4
X_14256_ _27266_/Q _26459_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _14256_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13207_ _13207_/A vssd1 vssd1 vccd1 vccd1 _14789_/A sky130_fd_sc_hd__buf_6
X_14187_ _14187_/A _16823_/B vssd1 vssd1 vccd1 vccd1 _14187_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _25808_/Q _15255_/A _16059_/S _13137_/X vssd1 vssd1 vccd1 vccd1 _13138_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _18742_/X _18985_/X _18994_/X vssd1 vssd1 vccd1 vccd1 _18995_/X sky130_fd_sc_hd__a21o_4
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _14089_/S vssd1 vssd1 vccd1 vccd1 _13998_/S sky130_fd_sc_hd__buf_2
X_17946_ _17821_/B _16206_/B _17950_/S vssd1 vssd1 vccd1 vccd1 _17946_/X sky130_fd_sc_hd__mux2_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17877_ _18058_/S vssd1 vssd1 vccd1 vccd1 _17958_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_38_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19616_ _27067_/Q _19616_/B _19616_/C vssd1 vssd1 vccd1 vccd1 _19616_/X sky130_fd_sc_hd__and3_1
XFILLER_94_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16828_ _16828_/A _16895_/A _16873_/B vssd1 vssd1 vccd1 vccd1 _16829_/A sky130_fd_sc_hd__and3_2
XFILLER_65_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19547_ _25653_/Q _19549_/B vssd1 vssd1 vccd1 vccd1 _19547_/X sky130_fd_sc_hd__or2_1
XFILLER_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16759_ _25679_/Q vssd1 vssd1 vccd1 vccd1 _22511_/A sky130_fd_sc_hd__buf_2
XFILLER_81_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19478_ _18929_/X _19476_/X _19477_/Y _18782_/X vssd1 vssd1 vccd1 vccd1 _19478_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18429_ _18366_/X _18428_/X _14023_/B vssd1 vssd1 vccd1 vccd1 _18429_/X sky130_fd_sc_hd__a21o_1
XFILLER_222_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21440_ _21421_/X _25863_/Q _21439_/Y _21386_/X vssd1 vssd1 vccd1 vccd1 _21440_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21371_ _25866_/Q vssd1 vssd1 vccd1 vccd1 _21646_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_175_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23110_ _23110_/A vssd1 vssd1 vccd1 vccd1 _26510_/D sky130_fd_sc_hd__clkbuf_1
X_20322_ _20291_/Y _20293_/Y _20339_/A _20320_/Y vssd1 vssd1 vccd1 vccd1 _20339_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_190_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24090_ _26913_/Q _23526_/X _24098_/S vssd1 vssd1 vccd1 vccd1 _24091_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23041_ _23514_/A vssd1 vssd1 vccd1 vccd1 _23041_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20253_ _20280_/B _20251_/Y _19600_/X _20252_/Y vssd1 vssd1 vccd1 vccd1 _20253_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_89_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20184_ _20184_/A _20184_/B vssd1 vssd1 vccd1 vccd1 _20184_/Y sky130_fd_sc_hd__xnor2_1
XTAP_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26800_ _27283_/CLK _26800_/D vssd1 vssd1 vccd1 vccd1 _26800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_276_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24992_ _24988_/X _24994_/B _24991_/X vssd1 vssd1 vccd1 vccd1 _24992_/X sky130_fd_sc_hd__a21bo_1
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26731_ _27311_/CLK _26731_/D vssd1 vssd1 vccd1 vccd1 _26731_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_257_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23943_ _26848_/Q _23523_/X _23943_/S vssd1 vssd1 vccd1 vccd1 _23944_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26662_ _27309_/CLK _26662_/D vssd1 vssd1 vccd1 vccd1 _26662_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23874_ _23702_/X _26817_/Q _23882_/S vssd1 vssd1 vccd1 vccd1 _23875_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25613_ _25660_/CLK _25613_/D vssd1 vssd1 vccd1 vccd1 _25613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22825_ _26394_/Q _22650_/X _22829_/S vssd1 vssd1 vccd1 vccd1 _22826_/A sky130_fd_sc_hd__mux2_1
X_26593_ _26593_/CLK _26593_/D vssd1 vssd1 vccd1 vccd1 _26593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25544_ _25545_/CLK _25544_/D vssd1 vssd1 vccd1 vccd1 _25544_/Q sky130_fd_sc_hd__dfxtp_1
X_22756_ _26364_/Q _22656_/X _22756_/S vssd1 vssd1 vccd1 vccd1 _22757_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21707_ _25992_/Q _21259_/X _21707_/S vssd1 vssd1 vccd1 vccd1 _21708_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25475_ _25590_/CLK _25475_/D vssd1 vssd1 vccd1 vccd1 _25475_/Q sky130_fd_sc_hd__dfxtp_2
X_22687_ _22687_/A vssd1 vssd1 vccd1 vccd1 _26341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27214_ _27221_/CLK _27214_/D vssd1 vssd1 vccd1 vccd1 _27214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24426_ _27015_/Q _24421_/X _24425_/Y _24415_/X vssd1 vssd1 vccd1 vccd1 _27015_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_197_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21638_ _21634_/Y _21637_/X _21202_/A vssd1 vssd1 vccd1 vccd1 _21638_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27145_ _27160_/CLK _27145_/D vssd1 vssd1 vccd1 vccd1 _27145_/Q sky130_fd_sc_hd__dfxtp_4
X_24357_ _24538_/A vssd1 vssd1 vccd1 vccd1 _24357_/X sky130_fd_sc_hd__clkbuf_2
X_21569_ _21569_/A vssd1 vssd1 vccd1 vccd1 _21569_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14110_ _26333_/Q _14103_/X _14178_/S _14109_/X vssd1 vssd1 vccd1 vccd1 _14110_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23308_ _23308_/A vssd1 vssd1 vccd1 vccd1 _26594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15090_ _14754_/A _15088_/X _15089_/X _14794_/A vssd1 vssd1 vccd1 vccd1 _15090_/X
+ sky130_fd_sc_hd__a211o_1
X_27076_ _27176_/CLK _27076_/D vssd1 vssd1 vccd1 vccd1 _27076_/Q sky130_fd_sc_hd__dfxtp_1
X_24288_ _26986_/Q _24286_/B _24287_/Y vssd1 vssd1 vccd1 vccd1 _26986_/D sky130_fd_sc_hd__o21a_1
XFILLER_158_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14041_ _27268_/Q _26461_/Q _14307_/S vssd1 vssd1 vccd1 vccd1 _14041_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26027_ _27293_/CLK _26027_/D vssd1 vssd1 vccd1 vccd1 _26027_/Q sky130_fd_sc_hd__dfxtp_1
X_23239_ _23239_/A vssd1 vssd1 vccd1 vccd1 _26563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17800_ _17800_/A _17986_/A _17800_/C vssd1 vssd1 vccd1 vccd1 _17802_/A sky130_fd_sc_hd__and3_1
X_15992_ _13608_/X _15983_/X _15991_/X _14713_/C vssd1 vssd1 vccd1 vccd1 _15992_/X
+ sky130_fd_sc_hd__a211o_1
X_18780_ _18552_/X _18739_/X _18778_/X _18779_/X vssd1 vssd1 vccd1 vccd1 _18780_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17731_ _26941_/Q _18460_/A _18462_/A _26973_/Q vssd1 vssd1 vccd1 vccd1 _17731_/X
+ sky130_fd_sc_hd__a22o_1
X_14943_ _12776_/A _26904_/Q _26776_/Q _14960_/B _14688_/A vssd1 vssd1 vccd1 vccd1
+ _14943_/X sky130_fd_sc_hd__a221o_1
XFILLER_94_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26929_ _26929_/CLK _26929_/D vssd1 vssd1 vccd1 vccd1 _26929_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14874_ _14867_/X _14873_/X _16221_/S vssd1 vssd1 vccd1 vccd1 _14874_/X sky130_fd_sc_hd__mux2_1
X_17662_ _17662_/A _17662_/B vssd1 vssd1 vccd1 vccd1 _19914_/A sky130_fd_sc_hd__or2_2
XFILLER_263_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19401_ _27162_/Q _19465_/B vssd1 vssd1 vccd1 vccd1 _19401_/X sky130_fd_sc_hd__or2_1
XFILLER_91_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13825_ _15606_/A _13823_/X _13824_/X _14228_/A vssd1 vssd1 vccd1 vccd1 _13825_/X
+ sky130_fd_sc_hd__a31o_1
X_16613_ _16613_/A _16613_/B vssd1 vssd1 vccd1 vccd1 _16762_/A sky130_fd_sc_hd__and2_2
XINSDIODE2_104 _21530_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17593_ _25917_/Q _17554_/X _17592_/X vssd1 vssd1 vccd1 vccd1 _17593_/Y sky130_fd_sc_hd__o21ai_1
XINSDIODE2_115 _22815_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_126 _23821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_137 _14621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16544_ _14804_/X _16540_/X _16543_/X _14818_/X vssd1 vssd1 vccd1 vccd1 _16544_/X
+ sky130_fd_sc_hd__o211a_1
X_19332_ _27096_/Q _19058_/X _19059_/X _27194_/Q _19060_/X vssd1 vssd1 vccd1 vccd1
+ _19332_/X sky130_fd_sc_hd__a221o_1
XINSDIODE2_148 _13304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13756_ _19847_/A _13756_/B vssd1 vssd1 vccd1 vccd1 _13756_/X sky130_fd_sc_hd__or2_1
XFILLER_189_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_159 _14777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12707_ _25591_/Q vssd1 vssd1 vccd1 vccd1 _19798_/A sky130_fd_sc_hd__buf_8
XFILLER_231_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19263_ _27062_/Q _18503_/X _19260_/X _19262_/X _18519_/X vssd1 vssd1 vccd1 vccd1
+ _19263_/X sky130_fd_sc_hd__o221a_2
X_16475_ _16473_/X _16474_/X _16479_/A vssd1 vssd1 vccd1 vccd1 _16475_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13687_ _13689_/A _13688_/A vssd1 vssd1 vccd1 vccd1 _18604_/S sky130_fd_sc_hd__and2_1
XFILLER_231_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15426_ _16259_/S vssd1 vssd1 vccd1 vccd1 _16347_/S sky130_fd_sc_hd__buf_4
X_18214_ _18214_/A vssd1 vssd1 vccd1 vccd1 _18548_/A sky130_fd_sc_hd__buf_2
X_19194_ _18602_/X _18547_/X _18544_/B _19358_/A vssd1 vssd1 vccd1 vccd1 _19194_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_157_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18145_ _14481_/X _18013_/X _18144_/Y _18022_/X _14407_/X vssd1 vssd1 vccd1 vccd1
+ _18146_/B sky130_fd_sc_hd__a32o_1
X_15357_ _16151_/S vssd1 vssd1 vccd1 vccd1 _16240_/S sky130_fd_sc_hd__buf_4
XFILLER_157_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14308_ _27266_/Q _26459_/Q _14308_/S vssd1 vssd1 vccd1 vccd1 _14308_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18076_ _18076_/A _18076_/B vssd1 vssd1 vccd1 vccd1 _18369_/A sky130_fd_sc_hd__nand2_2
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15288_ _15270_/X _15287_/X _15071_/A vssd1 vssd1 vccd1 vccd1 _15288_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17027_ _17021_/X _16880_/B _17025_/X input220/X vssd1 vssd1 vccd1 vccd1 _17027_/X
+ sky130_fd_sc_hd__a22o_4
X_14239_ _14239_/A _14239_/B vssd1 vssd1 vccd1 vccd1 _14239_/Y sky130_fd_sc_hd__nand2_1
XFILLER_171_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18978_ _18978_/A _18978_/B vssd1 vssd1 vccd1 vccd1 _19575_/A sky130_fd_sc_hd__xnor2_2
XFILLER_86_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _17810_/B _17779_/Y _18681_/A vssd1 vssd1 vccd1 vccd1 _17929_/X sky130_fd_sc_hd__mux2_1
XFILLER_273_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20940_ _25850_/Q _20939_/X _20949_/S vssd1 vssd1 vccd1 vccd1 _20941_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20871_ _20952_/A vssd1 vssd1 vccd1 vccd1 _20971_/S sky130_fd_sc_hd__buf_8
X_22610_ _26319_/Q _22618_/B vssd1 vssd1 vccd1 vccd1 _22610_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23590_ _23590_/A vssd1 vssd1 vccd1 vccd1 _23590_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_241_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22541_ _26293_/Q _22551_/B vssd1 vssd1 vccd1 vccd1 _22541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25260_ _23699_/X _27235_/Q _25260_/S vssd1 vssd1 vccd1 vccd1 _25261_/A sky130_fd_sc_hd__mux2_1
XFILLER_277_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22472_ _25757_/Q _22472_/B vssd1 vssd1 vccd1 vccd1 _22473_/A sky130_fd_sc_hd__and2_1
X_24211_ _26960_/Q _24213_/C _24210_/Y vssd1 vssd1 vccd1 vccd1 _26960_/D sky130_fd_sc_hd__o21a_1
XFILLER_182_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21423_ _21423_/A vssd1 vssd1 vccd1 vccd1 _21423_/Y sky130_fd_sc_hd__inv_2
X_25191_ _25199_/A vssd1 vssd1 vccd1 vccd1 _25191_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24142_ _26937_/Q _23603_/X _24142_/S vssd1 vssd1 vccd1 vccd1 _24143_/A sky130_fd_sc_hd__mux2_1
X_21354_ _21354_/A vssd1 vssd1 vccd1 vccd1 _21354_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20305_ _20305_/A _20305_/B _20305_/C vssd1 vssd1 vccd1 vccd1 _20305_/X sky130_fd_sc_hd__or3_1
XFILLER_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24073_ _24073_/A vssd1 vssd1 vccd1 vccd1 _26906_/D sky130_fd_sc_hd__clkbuf_1
X_21285_ _21285_/A vssd1 vssd1 vccd1 vccd1 _21286_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23024_ _26483_/Q _22730_/X _23028_/S vssd1 vssd1 vccd1 vccd1 _23025_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20236_ _20236_/A vssd1 vssd1 vccd1 vccd1 _20707_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_104_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_89_wb_clk_i _25501_/CLK vssd1 vssd1 vccd1 vccd1 _26813_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20167_ _20670_/A _20091_/A _20142_/Y _20119_/B _20144_/A vssd1 vssd1 vccd1 vccd1
+ _20174_/A sky130_fd_sc_hd__o221a_1
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27311_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24975_ _27159_/Q _24923_/B _24974_/Y _24970_/X vssd1 vssd1 vccd1 vccd1 _27159_/D
+ sky130_fd_sc_hd__o211a_1
X_20098_ _25676_/Q _25675_/Q _20098_/C vssd1 vssd1 vccd1 vccd1 _20151_/C sky130_fd_sc_hd__and3_1
XFILLER_57_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23926_ _23779_/X _26841_/Q _23926_/S vssd1 vssd1 vccd1 vccd1 _23927_/A sky130_fd_sc_hd__mux2_1
X_26714_ _27259_/CLK _26714_/D vssd1 vssd1 vccd1 vccd1 _26714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_268_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26645_ _27257_/CLK _26645_/D vssd1 vssd1 vccd1 vccd1 _26645_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23857_ _23857_/A vssd1 vssd1 vccd1 vccd1 _26810_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13610_ _13610_/A vssd1 vssd1 vccd1 vccd1 _13611_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22808_ _22808_/A vssd1 vssd1 vccd1 vccd1 _26387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14590_ _14590_/A vssd1 vssd1 vccd1 vccd1 _14591_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26576_ _26739_/CLK _26576_/D vssd1 vssd1 vccd1 vccd1 _26576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23788_ _23788_/A _23788_/B vssd1 vssd1 vccd1 vccd1 _23845_/A sky130_fd_sc_hd__or2_4
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13541_ _15843_/A vssd1 vssd1 vccd1 vccd1 _15401_/A sky130_fd_sc_hd__clkbuf_2
X_25527_ _25992_/CLK _25527_/D vssd1 vssd1 vccd1 vccd1 _25527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22739_ _23782_/A vssd1 vssd1 vccd1 vccd1 _22739_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16260_ _27286_/Q _26479_/Q _16260_/S vssd1 vssd1 vccd1 vccd1 _16260_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13472_ _13472_/A vssd1 vssd1 vccd1 vccd1 _13472_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25458_ _25458_/A vssd1 vssd1 vccd1 vccd1 _27323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15211_ _14743_/A _26708_/Q _26836_/Q _15228_/S _15210_/X vssd1 vssd1 vccd1 vccd1
+ _15211_/X sky130_fd_sc_hd__a221o_1
X_24409_ _27012_/Q _24391_/X _24408_/Y _24379_/X vssd1 vssd1 vccd1 vccd1 _27012_/D
+ sky130_fd_sc_hd__o211a_1
X_16191_ _14742_/A _26413_/Q _15301_/S _16190_/X vssd1 vssd1 vccd1 vccd1 _16191_/X
+ sky130_fd_sc_hd__o211a_1
X_25389_ _27293_/Q _23782_/A _25391_/S vssd1 vssd1 vccd1 vccd1 _25390_/A sky130_fd_sc_hd__mux2_1
X_27128_ _27130_/CLK _27128_/D vssd1 vssd1 vccd1 vccd1 _27128_/Q sky130_fd_sc_hd__dfxtp_4
X_15142_ _15142_/A vssd1 vssd1 vccd1 vccd1 _15142_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_154_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27059_ _27062_/CLK _27059_/D vssd1 vssd1 vccd1 vccd1 _27059_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_154_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19950_ _19950_/A _19977_/B vssd1 vssd1 vccd1 vccd1 _19951_/C sky130_fd_sc_hd__xnor2_1
X_15073_ _15073_/A vssd1 vssd1 vccd1 vccd1 _16463_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_141_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18901_ _18686_/B _19192_/B _18901_/S vssd1 vssd1 vccd1 vccd1 _18901_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14024_ _17813_/B vssd1 vssd1 vccd1 vccd1 _18423_/A sky130_fd_sc_hd__inv_2
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19881_ _19881_/A vssd1 vssd1 vccd1 vccd1 _19920_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18832_ _18832_/A vssd1 vssd1 vccd1 vccd1 _18832_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18763_ _18825_/A vssd1 vssd1 vccd1 vccd1 _18763_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_209_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ _13126_/A _15970_/X _15974_/X _13163_/A vssd1 vssd1 vccd1 vccd1 _15975_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_212_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17714_ _17753_/A vssd1 vssd1 vccd1 vccd1 _18161_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14926_ _14755_/A _14924_/X _14925_/X _14794_/A vssd1 vssd1 vccd1 vccd1 _14926_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_236_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18694_ _27112_/Q _18504_/X _18692_/X _18693_/X vssd1 vssd1 vccd1 vccd1 _18694_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_282_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17645_ _17560_/X _17627_/X _14033_/X _17544_/X _25931_/Q vssd1 vssd1 vccd1 vccd1
+ _17645_/Y sky130_fd_sc_hd__o32ai_4
X_14857_ _27292_/Q _26485_/Q _14878_/S vssd1 vssd1 vccd1 vccd1 _14857_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13808_ _13808_/A vssd1 vssd1 vccd1 vccd1 _13827_/A sky130_fd_sc_hd__buf_2
XFILLER_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17576_ _17634_/A vssd1 vssd1 vccd1 vccd1 _17595_/A sky130_fd_sc_hd__clkbuf_2
X_14788_ _20119_/A _14782_/X _14785_/X _14787_/X vssd1 vssd1 vccd1 vccd1 _14788_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_17_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19315_ _19315_/A _19346_/C vssd1 vssd1 vccd1 vccd1 _19315_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_232_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13739_ _14834_/A _14834_/B _14485_/A vssd1 vssd1 vccd1 vccd1 _15134_/A sky130_fd_sc_hd__nor3_1
X_16527_ _16513_/X _26907_/Q _26779_/Q _16526_/S _14773_/X vssd1 vssd1 vccd1 vccd1
+ _16527_/X sky130_fd_sc_hd__a221o_1
XFILLER_32_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19246_ _19246_/A _25747_/Q _19246_/C vssd1 vssd1 vccd1 vccd1 _19283_/B sky130_fd_sc_hd__and3_1
X_16458_ _16458_/A _16458_/B vssd1 vssd1 vccd1 vccd1 _19393_/A sky130_fd_sc_hd__and2_1
XFILLER_192_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15409_ _16194_/S vssd1 vssd1 vccd1 vccd1 _16273_/S sky130_fd_sc_hd__buf_4
X_16389_ _26091_/Q _16235_/S _16241_/S _16388_/X vssd1 vssd1 vccd1 vccd1 _16389_/X
+ sky130_fd_sc_hd__o211a_1
X_19177_ _18220_/X _19161_/X _19176_/X _18779_/X vssd1 vssd1 vccd1 vccd1 _19177_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18128_ _18172_/A vssd1 vssd1 vccd1 vccd1 _19069_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_144_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18059_ _18059_/A _18059_/B _18059_/C vssd1 vssd1 vccd1 vccd1 _18059_/X sky130_fd_sc_hd__and3_1
XFILLER_99_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21070_ _21070_/A _21070_/B _21197_/A vssd1 vssd1 vccd1 vccd1 _25901_/D sky130_fd_sc_hd__nor3_1
XFILLER_104_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20021_ _27114_/Q _19877_/X _19967_/X _20020_/Y vssd1 vssd1 vccd1 vccd1 _20021_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24760_ _24764_/A _24760_/B vssd1 vssd1 vccd1 vccd1 _27096_/D sky130_fd_sc_hd__nor2_1
X_21972_ _26100_/Q _20884_/X _21972_/S vssd1 vssd1 vccd1 vccd1 _21973_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23711_ _23711_/A vssd1 vssd1 vccd1 vccd1 _26755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20923_ _23738_/A vssd1 vssd1 vccd1 vccd1 _20923_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24691_ _27080_/Q _24680_/X _24690_/Y _24676_/X vssd1 vssd1 vccd1 vccd1 _24692_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26430_ _26462_/CLK _26430_/D vssd1 vssd1 vccd1 vccd1 _26430_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_270_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23642_ _23642_/A vssd1 vssd1 vccd1 vccd1 _26728_/D sky130_fd_sc_hd__clkbuf_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_270_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20854_ _25823_/Q vssd1 vssd1 vccd1 vccd1 _20855_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_230_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26361_ _27266_/CLK _26361_/D vssd1 vssd1 vccd1 vccd1 _26361_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_136_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27133_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23573_ _23573_/A vssd1 vssd1 vccd1 vccd1 _26703_/D sky130_fd_sc_hd__clkbuf_1
X_20785_ _20617_/X _25788_/Q _20787_/S vssd1 vssd1 vccd1 vccd1 _20786_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_490 _23584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_25312_ _25312_/A vssd1 vssd1 vccd1 vccd1 _27258_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22524_ _22524_/A _22524_/B vssd1 vssd1 vccd1 vccd1 _22525_/A sky130_fd_sc_hd__and2_1
XFILLER_210_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26292_ _26292_/CLK _26292_/D vssd1 vssd1 vccd1 vccd1 _26292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25243_ _27066_/Q _21873_/A input175/X _25214_/X _25178_/A vssd1 vssd1 vccd1 vccd1
+ _25243_/X sky130_fd_sc_hd__a41o_1
XFILLER_41_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22455_ _24415_/A vssd1 vssd1 vccd1 vccd1 _22455_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21406_ _20654_/A _21343_/X _21350_/X _21405_/X vssd1 vssd1 vccd1 vccd1 _21406_/X
+ sky130_fd_sc_hd__o211a_1
X_25174_ _25225_/A vssd1 vssd1 vccd1 vccd1 _25217_/A sky130_fd_sc_hd__clkbuf_2
X_22386_ _26239_/Q _22361_/A vssd1 vssd1 vccd1 vccd1 _22387_/A sky130_fd_sc_hd__or2b_1
XFILLER_163_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24125_ _26929_/Q _23578_/X _24131_/S vssd1 vssd1 vccd1 vccd1 _24126_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21337_ _21276_/X _21335_/X _21336_/X vssd1 vssd1 vccd1 vccd1 _21337_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_136_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24056_ _24056_/A vssd1 vssd1 vccd1 vccd1 _26898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21268_ _20628_/A _21277_/A _21279_/A _21267_/X vssd1 vssd1 vccd1 vccd1 _21268_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_249_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23007_ _23007_/A vssd1 vssd1 vccd1 vccd1 _26475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20219_ _27153_/Q _20219_/B vssd1 vssd1 vccd1 vccd1 _20219_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21199_ _21198_/Y _17455_/X _16679_/X vssd1 vssd1 vccd1 vccd1 _21199_/X sky130_fd_sc_hd__a21bo_1
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15760_ _15760_/A _15760_/B vssd1 vssd1 vccd1 vccd1 _15760_/X sky130_fd_sc_hd__or2_1
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24958_ _24600_/A _24941_/X _24938_/X vssd1 vssd1 vccd1 vccd1 _24958_/Y sky130_fd_sc_hd__a21oi_1
X_12972_ _25473_/Q _12961_/A _12969_/Y _12971_/X vssd1 vssd1 vccd1 vccd1 _12973_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _12706_/A _14697_/X _14707_/X _17195_/A vssd1 vssd1 vccd1 vccd1 _14711_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23909_ _23754_/X _26833_/Q _23915_/S vssd1 vssd1 vccd1 vccd1 _23910_/A sky130_fd_sc_hd__mux2_1
X_15691_ _14741_/A _26924_/Q _26408_/Q _16259_/S _13330_/A vssd1 vssd1 vccd1 vccd1
+ _15691_/X sky130_fd_sc_hd__a221o_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24889_ _24887_/Y _24888_/X _21242_/X vssd1 vssd1 vccd1 vccd1 _27129_/D sky130_fd_sc_hd__a21oi_1
XFILLER_61_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _17430_/A _17430_/B vssd1 vssd1 vccd1 vccd1 _17430_/Y sky130_fd_sc_hd__nor2_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14642_ _14948_/S vssd1 vssd1 vccd1 vccd1 _14693_/S sky130_fd_sc_hd__buf_2
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26628_ _27303_/CLK _26628_/D vssd1 vssd1 vccd1 vccd1 _26628_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17361_ _17380_/A _17361_/B _17362_/B vssd1 vssd1 vccd1 vccd1 _25539_/D sky130_fd_sc_hd__nor3_1
XFILLER_220_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14573_ _18423_/A _16720_/B _18428_/S vssd1 vssd1 vccd1 vccd1 _16723_/B sky130_fd_sc_hd__a21o_2
X_26559_ _27238_/CLK _26559_/D vssd1 vssd1 vccd1 vccd1 _26559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19100_ _19100_/A _19231_/B vssd1 vssd1 vccd1 vccd1 _19100_/Y sky130_fd_sc_hd__nor2_1
X_13524_ _14552_/S vssd1 vssd1 vccd1 vccd1 _13653_/S sky130_fd_sc_hd__buf_2
X_16312_ _16397_/S _16309_/X _16311_/X _15040_/A vssd1 vssd1 vccd1 vccd1 _16312_/X
+ sky130_fd_sc_hd__a211o_1
X_17292_ _17287_/X _17293_/C _25518_/Q vssd1 vssd1 vccd1 vccd1 _17294_/B sky130_fd_sc_hd__a21oi_1
XFILLER_40_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16243_ _25892_/Q _16243_/B vssd1 vssd1 vccd1 vccd1 _16243_/X sky130_fd_sc_hd__or2_1
X_19031_ _19031_/A _19374_/B vssd1 vssd1 vccd1 vccd1 _19031_/Y sky130_fd_sc_hd__nor2_1
XFILLER_186_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13455_ _13011_/A _23542_/A _13454_/X _13028_/A vssd1 vssd1 vccd1 vccd1 _16852_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_185_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16174_ _16336_/A _16172_/X _16173_/X vssd1 vssd1 vccd1 vccd1 _16174_/X sky130_fd_sc_hd__o21a_1
X_13386_ _12892_/A _13561_/A _13385_/X _12915_/A _25928_/Q vssd1 vssd1 vccd1 vccd1
+ _14323_/A sky130_fd_sc_hd__o32a_1
XFILLER_63_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15125_ _14787_/X _15117_/X _15124_/X _14724_/A vssd1 vssd1 vccd1 vccd1 _15125_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15056_ _15050_/X _15055_/X _16221_/S vssd1 vssd1 vccd1 vccd1 _15056_/X sky130_fd_sc_hd__mux2_1
X_19933_ _19933_/A _19933_/B _19933_/C vssd1 vssd1 vccd1 vccd1 _19935_/B sky130_fd_sc_hd__and3_1
XFILLER_123_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14007_ _13431_/X _14004_/X _14006_/X _13142_/A vssd1 vssd1 vccd1 vccd1 _14007_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_141_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19864_ _19870_/A _27075_/Q vssd1 vssd1 vccd1 vccd1 _19864_/X sky130_fd_sc_hd__or2_1
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18815_ _18815_/A vssd1 vssd1 vccd1 vccd1 _18815_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_268_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19795_ _20236_/A vssd1 vssd1 vccd1 vccd1 _20067_/A sky130_fd_sc_hd__buf_2
XFILLER_110_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18746_ _18810_/A vssd1 vssd1 vccd1 vccd1 _18746_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15958_ _25610_/Q _14594_/A _15957_/Y _12977_/A vssd1 vssd1 vccd1 vccd1 _15959_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput190 localMemory_wb_adr_i[0] vssd1 vssd1 vccd1 vccd1 input190/X sky130_fd_sc_hd__clkbuf_1
XFILLER_224_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14909_ _14746_/A _26125_/Q _26026_/Q _14981_/S _14772_/A vssd1 vssd1 vccd1 vccd1
+ _14909_/X sky130_fd_sc_hd__a221o_1
X_18677_ _18724_/B _18677_/B vssd1 vssd1 vccd1 vccd1 _19574_/B sky130_fd_sc_hd__and2b_1
XFILLER_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15889_ _15979_/S _15889_/B vssd1 vssd1 vccd1 vccd1 _15889_/X sky130_fd_sc_hd__or2_1
XFILLER_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17628_ _17560_/X _17627_/X _13736_/X _17554_/X _25926_/Q vssd1 vssd1 vccd1 vccd1
+ _17628_/Y sky130_fd_sc_hd__o32ai_2
XFILLER_252_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17559_ _17575_/A _17559_/B vssd1 vssd1 vccd1 vccd1 _25571_/D sky130_fd_sc_hd__nor2_1
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20570_ _23571_/A vssd1 vssd1 vccd1 vccd1 _23747_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19229_ _25525_/Q _18444_/A _19226_/X _19228_/X _18469_/A vssd1 vssd1 vccd1 vccd1
+ _19229_/X sky130_fd_sc_hd__o221a_1
XFILLER_176_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22240_ _22317_/A vssd1 vssd1 vccd1 vccd1 _22271_/A sky130_fd_sc_hd__buf_2
XFILLER_118_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22171_ _22249_/A vssd1 vssd1 vccd1 vccd1 _22171_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21122_ _21136_/A _21122_/B vssd1 vssd1 vccd1 vccd1 _21123_/A sky130_fd_sc_hd__or2_1
XFILLER_99_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25930_ _27221_/CLK _25930_/D vssd1 vssd1 vccd1 vccd1 _25930_/Q sky130_fd_sc_hd__dfxtp_4
X_21053_ _25895_/Q _20955_/X _21059_/S vssd1 vssd1 vccd1 vccd1 _21054_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20004_ _19991_/X _20002_/X _20003_/X vssd1 vssd1 vccd1 vccd1 _20004_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_59_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25861_ _27203_/CLK _25861_/D vssd1 vssd1 vccd1 vccd1 _25861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_275_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24812_ _20641_/A _24810_/X _24671_/Y _24811_/X vssd1 vssd1 vccd1 vccd1 _24812_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_25792_ _25796_/CLK _25792_/D vssd1 vssd1 vccd1 vccd1 _25792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24743_ _25466_/A vssd1 vssd1 vccd1 vccd1 _24764_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21955_ _20613_/X _26093_/Q _21955_/S vssd1 vssd1 vccd1 vccd1 _21956_/A sky130_fd_sc_hd__mux2_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20906_ _20906_/A vssd1 vssd1 vccd1 vccd1 _25839_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24674_ _24682_/A _24674_/B vssd1 vssd1 vccd1 vccd1 _24674_/Y sky130_fd_sc_hd__nand2_2
X_21886_ _21867_/Y _21884_/X _21885_/X _21878_/X vssd1 vssd1 vccd1 vccd1 _26063_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23625_ _23682_/S vssd1 vssd1 vccd1 vccd1 _23634_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_42_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26413_ _26609_/CLK _26413_/D vssd1 vssd1 vccd1 vccd1 _26413_/Q sky130_fd_sc_hd__dfxtp_1
X_20837_ _20837_/A vssd1 vssd1 vccd1 vccd1 _25814_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26344_ _26604_/CLK _26344_/D vssd1 vssd1 vccd1 vccd1 _26344_/Q sky130_fd_sc_hd__dfxtp_1
X_23556_ _26698_/Q _23555_/X _23556_/S vssd1 vssd1 vccd1 vccd1 _23557_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20768_ _20584_/X _25780_/Q _20772_/S vssd1 vssd1 vccd1 vccd1 _20769_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22507_ _22507_/A _22513_/B vssd1 vssd1 vccd1 vccd1 _22508_/A sky130_fd_sc_hd__and2_1
XFILLER_122_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26275_ _26282_/CLK _26275_/D vssd1 vssd1 vccd1 vccd1 _26275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23487_ _26674_/Q _23108_/X _23491_/S vssd1 vssd1 vccd1 vccd1 _23488_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20699_ _20699_/A _20707_/C vssd1 vssd1 vccd1 vccd1 _20699_/X sky130_fd_sc_hd__or2_1
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13240_ _13832_/A vssd1 vssd1 vccd1 vccd1 _13241_/A sky130_fd_sc_hd__clkbuf_4
X_25226_ _19617_/X _25209_/X _25179_/A vssd1 vssd1 vccd1 vccd1 _25226_/X sky130_fd_sc_hd__a21o_1
X_22438_ _26248_/Q _22444_/B vssd1 vssd1 vccd1 vccd1 _22438_/X sky130_fd_sc_hd__or2_1
XFILLER_182_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13171_ _13171_/A vssd1 vssd1 vccd1 vccd1 _13172_/A sky130_fd_sc_hd__buf_2
X_25157_ _22531_/A _25015_/X _25139_/X _17055_/B _25005_/X vssd1 vssd1 vccd1 vccd1
+ _25157_/X sky130_fd_sc_hd__a221o_1
XFILLER_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22369_ _22369_/A vssd1 vssd1 vccd1 vccd1 _26233_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24108_ _24108_/A vssd1 vssd1 vccd1 vccd1 _26921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26916_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_25088_ _22502_/A _25065_/X _25087_/X _18932_/B _25079_/X vssd1 vssd1 vccd1 vccd1
+ _25088_/X sky130_fd_sc_hd__a221o_1
XFILLER_151_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24039_ _24061_/A vssd1 vssd1 vccd1 vccd1 _24048_/S sky130_fd_sc_hd__buf_2
X_16930_ _16986_/A _16930_/B vssd1 vssd1 vccd1 vccd1 _16931_/A sky130_fd_sc_hd__and2_1
XFILLER_2_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16861_ _16906_/A vssd1 vssd1 vccd1 vccd1 _16868_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18600_ _18426_/Y _18599_/Y _18685_/S vssd1 vssd1 vccd1 vccd1 _18600_/X sky130_fd_sc_hd__mux2_1
X_15812_ _13114_/A _15799_/X _15803_/X _15811_/X _13168_/A vssd1 vssd1 vccd1 vccd1
+ _15812_/X sky130_fd_sc_hd__a311o_1
XFILLER_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19580_ _18905_/B _18855_/Y _19189_/Y _19579_/Y _18795_/Y vssd1 vssd1 vccd1 vccd1
+ _19581_/C sky130_fd_sc_hd__a2111o_1
X_16792_ _16973_/B _16794_/B _19639_/B _16955_/B _16982_/B vssd1 vssd1 vccd1 vccd1
+ _16792_/X sky130_fd_sc_hd__o2111a_4
XFILLER_237_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18531_ _18588_/C _18531_/B vssd1 vssd1 vccd1 vccd1 _18531_/X sky130_fd_sc_hd__or2_1
X_15743_ _26079_/Q _15961_/B _14107_/X _15742_/X vssd1 vssd1 vccd1 vccd1 _15743_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_206_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12955_ _12959_/A _25477_/Q vssd1 vssd1 vccd1 vccd1 _13197_/A sky130_fd_sc_hd__or2b_2
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18462_ _18462_/A vssd1 vssd1 vccd1 vccd1 _18463_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_261_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _12860_/B _12878_/Y _12941_/A _14407_/A vssd1 vssd1 vccd1 vccd1 _15706_/B
+ sky130_fd_sc_hd__a31oi_2
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _16193_/S vssd1 vssd1 vccd1 vccd1 _15674_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _25556_/Q vssd1 vssd1 vccd1 vccd1 _17418_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14625_ _16144_/S vssd1 vssd1 vccd1 vccd1 _15263_/S sky130_fd_sc_hd__buf_4
XFILLER_260_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18393_ _18817_/A vssd1 vssd1 vccd1 vccd1 _18510_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_199_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _25534_/Q _17344_/B vssd1 vssd1 vccd1 vccd1 _17351_/C sky130_fd_sc_hd__and2_1
X_14556_ _13278_/A _14552_/X _14555_/X _13310_/A vssd1 vssd1 vccd1 vccd1 _14556_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13507_ _12982_/A _13577_/A _13204_/B _13204_/C vssd1 vssd1 vccd1 vccd1 _13508_/A
+ sky130_fd_sc_hd__o211a_2
X_17275_ _25513_/Q _17275_/B vssd1 vssd1 vccd1 vccd1 _17282_/C sky130_fd_sc_hd__and2_1
X_14487_ _14484_/X _14486_/X _14401_/A vssd1 vssd1 vccd1 vccd1 _14528_/A sky130_fd_sc_hd__a21o_1
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19014_ _18040_/X _18211_/X _18191_/X _18321_/A vssd1 vssd1 vccd1 vccd1 _19018_/B
+ sky130_fd_sc_hd__o211a_1
X_13438_ _26106_/Q _26007_/Q _15964_/S vssd1 vssd1 vccd1 vccd1 _13438_/X sky130_fd_sc_hd__mux2_1
X_16226_ _12774_/A _26707_/Q _26835_/Q _16385_/S _15048_/X vssd1 vssd1 vccd1 vccd1
+ _16226_/X sky130_fd_sc_hd__a221o_1
XFILLER_127_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16157_ _16154_/X _16155_/X _16156_/X _15376_/S _15647_/S vssd1 vssd1 vccd1 vccd1
+ _16157_/X sky130_fd_sc_hd__a221o_1
X_13369_ _13369_/A _13369_/B vssd1 vssd1 vccd1 vccd1 _13369_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ _26646_/Q _26742_/Q _15119_/S vssd1 vssd1 vccd1 vccd1 _15108_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16088_ _16088_/A _16088_/B vssd1 vssd1 vccd1 vccd1 _16088_/X sky130_fd_sc_hd__or2_1
XFILLER_142_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19916_ _19916_/A _20249_/B vssd1 vssd1 vccd1 vccd1 _19978_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15039_ _15039_/A vssd1 vssd1 vccd1 vccd1 _15040_/A sky130_fd_sc_hd__buf_4
XFILLER_130_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19847_ _19847_/A _20249_/B vssd1 vssd1 vccd1 vccd1 _19852_/A sky130_fd_sc_hd__nand2_1
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19778_ _19853_/B _19778_/B vssd1 vssd1 vccd1 vccd1 _19778_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_271_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18729_ _18729_/A _18729_/B vssd1 vssd1 vccd1 vccd1 _18729_/X sky130_fd_sc_hd__or2_1
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21740_ _21740_/A vssd1 vssd1 vccd1 vccd1 _26004_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21671_ _21671_/A vssd1 vssd1 vccd1 vccd1 _25975_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23410_ _23421_/A vssd1 vssd1 vccd1 vccd1 _23419_/S sky130_fd_sc_hd__buf_4
X_20622_ _20621_/X _25723_/Q _20622_/S vssd1 vssd1 vccd1 vccd1 _20623_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24390_ _24390_/A vssd1 vssd1 vccd1 vccd1 _24506_/A sky130_fd_sc_hd__buf_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23341_ _23341_/A vssd1 vssd1 vccd1 vccd1 _26609_/D sky130_fd_sc_hd__clkbuf_1
X_20553_ _23558_/A vssd1 vssd1 vccd1 vccd1 _23734_/A sky130_fd_sc_hd__buf_2
XFILLER_138_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26060_ _26683_/CLK _26060_/D vssd1 vssd1 vccd1 vccd1 _26060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23272_ _23272_/A vssd1 vssd1 vccd1 vccd1 _26578_/D sky130_fd_sc_hd__clkbuf_1
X_20484_ _23684_/A vssd1 vssd1 vccd1 vccd1 _20484_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25011_ _20626_/A _25003_/X _25010_/X vssd1 vssd1 vccd1 vccd1 _25011_/Y sky130_fd_sc_hd__o21ai_1
X_22223_ input7/X input282/X _22226_/S vssd1 vssd1 vccd1 vccd1 _22223_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_1_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _26681_/CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_180_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22154_ _22154_/A vssd1 vssd1 vccd1 vccd1 _22154_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput450 _25724_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[0] sky130_fd_sc_hd__buf_2
Xoutput461 _25725_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[1] sky130_fd_sc_hd__buf_2
XFILLER_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21105_ _21105_/A vssd1 vssd1 vccd1 vccd1 _25909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput472 _25726_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[2] sky130_fd_sc_hd__buf_2
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26962_ _26992_/CLK _26962_/D vssd1 vssd1 vccd1 vccd1 _26962_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput483 _16678_/Y vssd1 vssd1 vccd1 vccd1 web0 sky130_fd_sc_hd__buf_2
X_22085_ _22085_/A vssd1 vssd1 vccd1 vccd1 _26150_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21036_ _21036_/A vssd1 vssd1 vccd1 vccd1 _25887_/D sky130_fd_sc_hd__clkbuf_1
X_25913_ _27117_/CLK _25913_/D vssd1 vssd1 vccd1 vccd1 _25913_/Q sky130_fd_sc_hd__dfxtp_4
X_26893_ _27311_/CLK _26893_/D vssd1 vssd1 vccd1 vccd1 _26893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25844_ _26531_/CLK _25844_/D vssd1 vssd1 vccd1 vccd1 _25844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_274_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_151_wb_clk_i clkbuf_opt_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27221_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22987_ _26466_/Q _22675_/X _22995_/S vssd1 vssd1 vccd1 vccd1 _22988_/A sky130_fd_sc_hd__mux2_1
X_25775_ _27280_/CLK _25775_/D vssd1 vssd1 vccd1 vccd1 _25775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12740_ _17669_/C _12740_/B _12740_/C vssd1 vssd1 vccd1 vccd1 _19570_/B sky130_fd_sc_hd__or3_4
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21938_ _20580_/X _26085_/Q _21944_/S vssd1 vssd1 vccd1 vccd1 _21939_/A sky130_fd_sc_hd__mux2_1
X_24726_ _27088_/Q _24724_/X _24725_/Y _24720_/X vssd1 vssd1 vccd1 vccd1 _24727_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _16641_/A vssd1 vssd1 vccd1 vccd1 _12671_/Y sky130_fd_sc_hd__inv_2
X_24657_ _24701_/A vssd1 vssd1 vccd1 vccd1 _24657_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_242_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21869_ _24455_/A vssd1 vssd1 vccd1 vccd1 _21869_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14485_/B vssd1 vssd1 vccd1 vccd1 _14410_/Y sky130_fd_sc_hd__inv_2
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23608_ _23608_/A vssd1 vssd1 vccd1 vccd1 _26714_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _16170_/A _16916_/A vssd1 vssd1 vccd1 vccd1 _15390_/Y sky130_fd_sc_hd__nor2_1
X_24588_ _27051_/Q _24576_/X _24587_/Y _24580_/X vssd1 vssd1 vccd1 vccd1 _27051_/D
+ sky130_fd_sc_hd__o211a_1
X_14341_ _14440_/S _14330_/X _14334_/X _14340_/X vssd1 vssd1 vccd1 vccd1 _14341_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_211_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26327_ _26327_/CLK _26327_/D vssd1 vssd1 vccd1 vccd1 _26327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23539_ _23539_/A vssd1 vssd1 vccd1 vccd1 _23539_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17060_ _17060_/A vssd1 vssd1 vccd1 vccd1 _17061_/A sky130_fd_sc_hd__clkbuf_2
X_26258_ _26974_/CLK _26258_/D vssd1 vssd1 vccd1 vccd1 _26258_/Q sky130_fd_sc_hd__dfxtp_1
X_14272_ _14269_/X _14271_/X _14272_/S vssd1 vssd1 vccd1 vccd1 _14272_/X sky130_fd_sc_hd__mux2_2
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16011_ _16007_/X _16010_/X _13543_/A vssd1 vssd1 vccd1 vccd1 _16011_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13223_ _14472_/S vssd1 vssd1 vccd1 vccd1 _14536_/S sky130_fd_sc_hd__buf_2
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25209_ _25214_/A vssd1 vssd1 vccd1 vccd1 _25209_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26189_ _26222_/CLK _26189_/D vssd1 vssd1 vccd1 vccd1 _26189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13154_ _27274_/Q _26467_/Q _15467_/S vssd1 vssd1 vccd1 vccd1 _13154_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _13085_/A vssd1 vssd1 vccd1 vccd1 _13694_/A sky130_fd_sc_hd__buf_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _17986_/A vssd1 vssd1 vccd1 vccd1 _18343_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19701_ _20252_/B _18229_/X _19600_/X _19700_/Y vssd1 vssd1 vccd1 vccd1 _19701_/X
+ sky130_fd_sc_hd__o31a_1
X_16913_ _16907_/X _16963_/C _16912_/X vssd1 vssd1 vccd1 vccd1 _16914_/B sky130_fd_sc_hd__o21a_2
XFILLER_78_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17893_ _17975_/A vssd1 vssd1 vccd1 vccd1 _18197_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_265_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19632_ _21195_/B _19639_/B _12778_/B vssd1 vssd1 vccd1 vccd1 _19634_/B sky130_fd_sc_hd__o21a_1
X_16844_ _16864_/A _16844_/B vssd1 vssd1 vccd1 vccd1 _16845_/A sky130_fd_sc_hd__and2_1
XFILLER_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19563_ _25659_/Q _19563_/B vssd1 vssd1 vccd1 vccd1 _19563_/X sky130_fd_sc_hd__or2_1
X_16775_ _25685_/Q vssd1 vssd1 vccd1 vccd1 _22524_/A sky130_fd_sc_hd__clkbuf_4
X_13987_ _26102_/Q _26003_/Q _14253_/S vssd1 vssd1 vccd1 vccd1 _13987_/X sky130_fd_sc_hd__mux2_1
XFILLER_280_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18514_ _18514_/A vssd1 vssd1 vccd1 vccd1 _18514_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15726_ _26111_/Q _26012_/Q _15726_/S vssd1 vssd1 vccd1 vccd1 _15726_/X sky130_fd_sc_hd__mux2_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19494_ _19484_/X _18177_/X _19493_/X _19489_/X vssd1 vssd1 vccd1 vccd1 _25632_/D
+ sky130_fd_sc_hd__o211a_1
X_12938_ _13748_/A vssd1 vssd1 vccd1 vccd1 _14404_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18445_ _27107_/Q _18812_/A vssd1 vssd1 vccd1 vccd1 _18445_/X sky130_fd_sc_hd__or2_1
XFILLER_209_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15657_ _15639_/X _15656_/X _14591_/A vssd1 vssd1 vccd1 vccd1 _15657_/X sky130_fd_sc_hd__a21o_2
X_12869_ _12869_/A vssd1 vssd1 vccd1 vccd1 _12869_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14608_ _16212_/B vssd1 vssd1 vccd1 vccd1 _14609_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_178_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18376_ _18352_/Y _18360_/X _18374_/Y _18375_/X vssd1 vssd1 vccd1 vccd1 _18376_/X
+ sky130_fd_sc_hd__o31a_1
X_15588_ _15588_/A vssd1 vssd1 vccd1 vccd1 _15589_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17327_ _25529_/Q vssd1 vssd1 vccd1 vccd1 _17327_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14539_ _26520_/Q _26128_/Q _14539_/S vssd1 vssd1 vccd1 vccd1 _14539_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17258_ _17263_/C _17258_/B vssd1 vssd1 vccd1 vccd1 _25507_/D sky130_fd_sc_hd__nor2_1
XFILLER_88_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16209_ _16206_/Y _19105_/S _16207_/A vssd1 vssd1 vccd1 vccd1 _16209_/X sky130_fd_sc_hd__a21o_1
XFILLER_162_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17189_ _16480_/S _17170_/X _17185_/X _17188_/X vssd1 vssd1 vccd1 vccd1 _25489_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_7_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22910_ _26432_/Q _22669_/X _22912_/S vssd1 vssd1 vccd1 vccd1 _22911_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23890_ _23890_/A vssd1 vssd1 vccd1 vccd1 _26824_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22841_ _22841_/A vssd1 vssd1 vccd1 vccd1 _26401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25560_ _27000_/CLK _25560_/D vssd1 vssd1 vccd1 vccd1 _25560_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22772_ _26371_/Q _22679_/X _22778_/S vssd1 vssd1 vccd1 vccd1 _22773_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24511_ _26319_/Q _21869_/X _21871_/X input233/X _24501_/X vssd1 vssd1 vccd1 vccd1
+ _24511_/X sky130_fd_sc_hd__a221o_1
X_21723_ _21791_/S vssd1 vssd1 vccd1 vccd1 _21732_/S sky130_fd_sc_hd__buf_2
XFILLER_25_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25491_ _26683_/CLK _25491_/D vssd1 vssd1 vccd1 vccd1 _25491_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_197_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24442_ _24551_/A vssd1 vssd1 vccd1 vccd1 _24442_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_27230_ _27230_/CLK _27230_/D vssd1 vssd1 vccd1 vccd1 _27230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21654_ _20487_/B _21349_/B _21654_/C _21654_/D vssd1 vssd1 vccd1 vccd1 _21698_/A
+ sky130_fd_sc_hd__and4bb_4
XFILLER_220_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27161_ _27164_/CLK _27161_/D vssd1 vssd1 vccd1 vccd1 _27161_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20605_ _23773_/A vssd1 vssd1 vccd1 vccd1 _20605_/X sky130_fd_sc_hd__clkbuf_2
X_24373_ _27007_/Q _24357_/X _24372_/Y _22468_/X vssd1 vssd1 vccd1 vccd1 _27007_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21585_ _25494_/Q _21620_/B vssd1 vssd1 vccd1 vccd1 _21585_/X sky130_fd_sc_hd__or2_1
X_26112_ _26673_/CLK _26112_/D vssd1 vssd1 vccd1 vccd1 _26112_/Q sky130_fd_sc_hd__dfxtp_1
X_23324_ _20550_/X _26602_/Q _23324_/S vssd1 vssd1 vccd1 vccd1 _23325_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20536_ _20536_/A vssd1 vssd1 vccd1 vccd1 _25702_/D sky130_fd_sc_hd__clkbuf_1
X_27092_ _27228_/CLK _27092_/D vssd1 vssd1 vccd1 vccd1 _27092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26043_ _26599_/CLK _26043_/D vssd1 vssd1 vccd1 vccd1 _26043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23255_ _26571_/Q _23098_/X _23255_/S vssd1 vssd1 vccd1 vccd1 _23256_/A sky130_fd_sc_hd__mux2_1
X_20467_ _25691_/Q _25690_/Q _20467_/C vssd1 vssd1 vccd1 vccd1 _20467_/X sky130_fd_sc_hd__and3_1
XFILLER_4_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22206_ _22206_/A vssd1 vssd1 vccd1 vccd1 _22206_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_279_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23186_ _26540_/Q _23101_/X _23194_/S vssd1 vssd1 vccd1 vccd1 _23187_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20398_ _20398_/A _20398_/B vssd1 vssd1 vccd1 vccd1 _20398_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22137_ _22155_/A vssd1 vssd1 vccd1 vccd1 _22137_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput291 _17069_/X vssd1 vssd1 vccd1 vccd1 addr0[6] sky130_fd_sc_hd__buf_2
X_26945_ _26980_/CLK _26945_/D vssd1 vssd1 vccd1 vccd1 _26945_/Q sky130_fd_sc_hd__dfxtp_1
X_22068_ _22090_/A vssd1 vssd1 vccd1 vccd1 _22077_/S sky130_fd_sc_hd__buf_4
XFILLER_121_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21019_ _21019_/A vssd1 vssd1 vccd1 vccd1 _25879_/D sky130_fd_sc_hd__clkbuf_1
X_13910_ _17813_/A vssd1 vssd1 vccd1 vccd1 _18482_/A sky130_fd_sc_hd__inv_2
X_26876_ _26877_/CLK _26876_/D vssd1 vssd1 vccd1 vccd1 _26876_/Q sky130_fd_sc_hd__dfxtp_1
X_14890_ _14890_/A vssd1 vssd1 vccd1 vccd1 _14890_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_247_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13841_ _13841_/A vssd1 vssd1 vccd1 vccd1 _15775_/S sky130_fd_sc_hd__buf_4
X_25827_ _26917_/CLK _25827_/D vssd1 vssd1 vccd1 vccd1 _25827_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13772_ _13488_/A _25766_/Q _15514_/S _26852_/Q _13512_/A vssd1 vssd1 vccd1 vccd1
+ _13772_/X sky130_fd_sc_hd__o221a_1
XINSDIODE2_308 _25927_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16560_ _16560_/A vssd1 vssd1 vccd1 vccd1 _16561_/A sky130_fd_sc_hd__inv_2
X_25758_ _26909_/CLK _25758_/D vssd1 vssd1 vccd1 vccd1 _25758_/Q sky130_fd_sc_hd__dfxtp_2
XINSDIODE2_319 _19616_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15511_ _15491_/X _25847_/Q _26047_/Q _15850_/S _13806_/X vssd1 vssd1 vccd1 vccd1
+ _15511_/X sky130_fd_sc_hd__a221o_1
X_12723_ _25578_/Q vssd1 vssd1 vccd1 vccd1 _17669_/A sky130_fd_sc_hd__clkbuf_2
X_24709_ _24722_/A _24709_/B vssd1 vssd1 vccd1 vccd1 _27084_/D sky130_fd_sc_hd__nor2_1
XFILLER_243_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16491_ _17712_/B _26423_/Q _16480_/S _16490_/X vssd1 vssd1 vccd1 vccd1 _16491_/X
+ sky130_fd_sc_hd__o211a_1
X_25689_ _25690_/CLK _25689_/D vssd1 vssd1 vccd1 vccd1 _25689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18230_ _19219_/A _18230_/B vssd1 vssd1 vccd1 vccd1 _18230_/Y sky130_fd_sc_hd__nand2_1
X_15442_ _12913_/A _13391_/X _14603_/A vssd1 vssd1 vccd1 vccd1 _15442_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_230_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18161_ _18161_/A _18161_/B _18161_/C vssd1 vssd1 vccd1 vccd1 _18232_/A sky130_fd_sc_hd__or3_1
XFILLER_8_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15373_ _15371_/X _15372_/X _15384_/S vssd1 vssd1 vccd1 vccd1 _15373_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17112_ _25465_/S vssd1 vssd1 vccd1 vccd1 _17612_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_129_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14324_ _14411_/A _13391_/X _13397_/X _14323_/Y vssd1 vssd1 vccd1 vccd1 _14324_/X
+ sky130_fd_sc_hd__o211a_1
X_18092_ _18092_/A _18552_/A vssd1 vssd1 vccd1 vccd1 _18927_/A sky130_fd_sc_hd__nor2_1
XFILLER_239_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14255_ _15903_/S vssd1 vssd1 vccd1 vccd1 _15990_/S sky130_fd_sc_hd__clkbuf_8
X_17043_ _17042_/X _16949_/B _17039_/X input232/X vssd1 vssd1 vccd1 vccd1 _17043_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_183_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ _13638_/A vssd1 vssd1 vccd1 vccd1 _13207_/A sky130_fd_sc_hd__buf_6
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14186_ _13008_/A _23523_/A _14185_/X vssd1 vssd1 vccd1 vccd1 _16823_/B sky130_fd_sc_hd__o21ai_4
XFILLER_124_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13137_ _27242_/Q _15635_/B vssd1 vssd1 vccd1 vccd1 _13137_/X sky130_fd_sc_hd__or2_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18994_ _25518_/Q _18746_/X _18991_/X _18993_/X _18770_/X vssd1 vssd1 vccd1 vccd1
+ _18994_/X sky130_fd_sc_hd__o221a_1
XFILLER_124_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _13068_/A vssd1 vssd1 vccd1 vccd1 _14089_/S sky130_fd_sc_hd__buf_2
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _18349_/S vssd1 vssd1 vccd1 vccd1 _18896_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_79_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17876_ _14022_/A _17784_/B _17909_/S vssd1 vssd1 vccd1 vccd1 _17876_/X sky130_fd_sc_hd__mux2_2
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19615_ _19617_/B vssd1 vssd1 vccd1 vccd1 _21264_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16827_ _16982_/B _16827_/B vssd1 vssd1 vccd1 vccd1 _16873_/B sky130_fd_sc_hd__and2_2
XFILLER_253_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19546_ _19538_/X _19172_/X _19545_/X _19541_/X vssd1 vssd1 vccd1 vccd1 _25652_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16758_ _22509_/A _16756_/X _16757_/X _16637_/B vssd1 vssd1 vccd1 vccd1 _16758_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_207_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15709_ _12871_/Y _15705_/X _15707_/X _12943_/Y _15708_/Y vssd1 vssd1 vccd1 vccd1
+ _15709_/X sky130_fd_sc_hd__a32o_1
XFILLER_234_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19477_ _25755_/Q _19477_/B vssd1 vssd1 vccd1 vccd1 _19477_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_222_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16689_ _16689_/A vssd1 vssd1 vccd1 vccd1 _16689_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_210_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18428_ _18368_/X _18371_/X _18428_/S vssd1 vssd1 vccd1 vccd1 _18428_/X sky130_fd_sc_hd__mux2_1
XFILLER_250_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18359_ _18636_/A vssd1 vssd1 vccd1 vccd1 _18359_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_222_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21370_ _21342_/X _21369_/X _21336_/X vssd1 vssd1 vccd1 vccd1 _21370_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_108_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20321_ _20339_/A _20320_/Y _20291_/Y _20293_/Y vssd1 vssd1 vccd1 vccd1 _20321_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_190_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23040_ _23040_/A vssd1 vssd1 vccd1 vccd1 _26488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20252_ _20252_/A _20252_/B vssd1 vssd1 vccd1 vccd1 _20252_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20183_ _20160_/A _20159_/A _20158_/Y vssd1 vssd1 vccd1 vccd1 _20184_/B sky130_fd_sc_hd__o21a_1
XFILLER_249_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24991_ _24989_/X _24544_/B _24654_/A _24986_/Y vssd1 vssd1 vccd1 vccd1 _24991_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26730_ _27309_/CLK _26730_/D vssd1 vssd1 vccd1 vccd1 _26730_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23942_ _23942_/A vssd1 vssd1 vccd1 vccd1 _26847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26661_ _27303_/CLK _26661_/D vssd1 vssd1 vccd1 vccd1 _26661_/Q sky130_fd_sc_hd__dfxtp_1
X_23873_ _23930_/S vssd1 vssd1 vccd1 vccd1 _23882_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_29_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22824_ _22824_/A vssd1 vssd1 vccd1 vccd1 _26393_/D sky130_fd_sc_hd__clkbuf_1
X_25612_ _25660_/CLK _25612_/D vssd1 vssd1 vccd1 vccd1 _25612_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_232_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26592_ _26592_/CLK _26592_/D vssd1 vssd1 vccd1 vccd1 _26592_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_204_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22755_ _22755_/A vssd1 vssd1 vccd1 vccd1 _26363_/D sky130_fd_sc_hd__clkbuf_1
X_25543_ _25545_/CLK _25543_/D vssd1 vssd1 vccd1 vccd1 _25543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21706_ _21706_/A vssd1 vssd1 vccd1 vccd1 _25991_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25474_ _25598_/CLK _25474_/D vssd1 vssd1 vccd1 vccd1 _25474_/Q sky130_fd_sc_hd__dfxtp_1
X_22686_ _26341_/Q _22685_/X _22689_/S vssd1 vssd1 vccd1 vccd1 _22687_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24425_ _24434_/A _24577_/A vssd1 vssd1 vccd1 vccd1 _24425_/Y sky130_fd_sc_hd__nand2_1
XFILLER_197_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27213_ _27213_/CLK _27213_/D vssd1 vssd1 vccd1 vccd1 _27213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21637_ _21354_/A _25865_/Q _21636_/Y _21237_/X vssd1 vssd1 vccd1 vccd1 _21637_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24356_ _24390_/A vssd1 vssd1 vccd1 vccd1 _24538_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_165_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27144_ _27164_/CLK _27144_/D vssd1 vssd1 vccd1 vccd1 _27144_/Q sky130_fd_sc_hd__dfxtp_2
X_21568_ input59/X input94/X _21615_/S vssd1 vssd1 vccd1 vccd1 _21569_/A sky130_fd_sc_hd__mux2_8
XFILLER_138_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23307_ _20517_/X _26594_/Q _23313_/S vssd1 vssd1 vccd1 vccd1 _23308_/A sky130_fd_sc_hd__mux2_1
X_20519_ _20519_/A vssd1 vssd1 vccd1 vccd1 _25698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27075_ _27203_/CLK _27075_/D vssd1 vssd1 vccd1 vccd1 _27075_/Q sky130_fd_sc_hd__dfxtp_1
X_24287_ _24312_/A _24293_/C vssd1 vssd1 vccd1 vccd1 _24287_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21499_ _21480_/X _21498_/X _21473_/X vssd1 vssd1 vccd1 vccd1 _21499_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_154_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14040_ _25635_/Q _13803_/B _13578_/A _25603_/Q _14039_/X vssd1 vssd1 vccd1 vccd1
+ _23526_/A sky130_fd_sc_hd__a221o_4
X_23238_ _26563_/Q _23073_/X _23244_/S vssd1 vssd1 vccd1 vccd1 _23239_/A sky130_fd_sc_hd__mux2_1
X_26026_ _27291_/CLK _26026_/D vssd1 vssd1 vccd1 vccd1 _26026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23169_ _23169_/A vssd1 vssd1 vccd1 vccd1 _26532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_279_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ _15985_/X _15987_/X _15990_/X _15819_/S _13630_/X vssd1 vssd1 vccd1 vccd1
+ _15991_/X sky130_fd_sc_hd__o221a_1
XTAP_5731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17730_ _17730_/A _17730_/B vssd1 vssd1 vccd1 vccd1 _18462_/A sky130_fd_sc_hd__and2_2
XTAP_5753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26928_ _27316_/CLK _26928_/D vssd1 vssd1 vccd1 vccd1 _26928_/Q sky130_fd_sc_hd__dfxtp_1
X_14942_ _26680_/Q _25720_/Q _14953_/S vssd1 vssd1 vccd1 vccd1 _14942_/X sky130_fd_sc_hd__mux2_1
XTAP_5764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17661_ _18785_/A vssd1 vssd1 vccd1 vccd1 _18005_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_236_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26859_ _27311_/CLK _26859_/D vssd1 vssd1 vccd1 vccd1 _26859_/Q sky130_fd_sc_hd__dfxtp_2
X_14873_ _14868_/X _14869_/X _14877_/S vssd1 vssd1 vccd1 vccd1 _14873_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19400_ _27130_/Q _19056_/X _19398_/X _19399_/X vssd1 vssd1 vccd1 vccd1 _19400_/X
+ sky130_fd_sc_hd__o22a_2
X_16612_ _16612_/A _16612_/B vssd1 vssd1 vccd1 vccd1 _16613_/B sky130_fd_sc_hd__nand2_1
XFILLER_75_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13824_ _13472_/A _26883_/Q _26755_/Q _15758_/S _13358_/A vssd1 vssd1 vccd1 vccd1
+ _13824_/X sky130_fd_sc_hd__a221o_1
XFILLER_251_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17592_ _17592_/A _17592_/B _17592_/C vssd1 vssd1 vccd1 vccd1 _17592_/X sky130_fd_sc_hd__or3_1
XFILLER_63_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_105 _21557_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_116 _22815_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19331_ _27226_/Q _19331_/B vssd1 vssd1 vccd1 vccd1 _19331_/X sky130_fd_sc_hd__and2_1
XINSDIODE2_127 _12674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_138 _13529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16543_ _14755_/X _16541_/X _16542_/X _14794_/X vssd1 vssd1 vccd1 vccd1 _16543_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13755_ _25593_/Q vssd1 vssd1 vccd1 vccd1 _19847_/A sky130_fd_sc_hd__buf_8
XFILLER_204_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_149 _13335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19262_ _27030_/Q _18514_/X _19261_/X _18455_/X vssd1 vssd1 vccd1 vccd1 _19262_/X
+ sky130_fd_sc_hd__a22o_1
X_12706_ _12706_/A vssd1 vssd1 vccd1 vccd1 _12722_/B sky130_fd_sc_hd__buf_6
XFILLER_93_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16474_ _26127_/Q _26028_/Q _16498_/S vssd1 vssd1 vccd1 vccd1 _16474_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13686_ _14566_/A _19882_/A _13685_/X vssd1 vssd1 vccd1 vccd1 _13688_/A sky130_fd_sc_hd__o21a_1
XFILLER_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18213_ _18603_/A vssd1 vssd1 vccd1 vccd1 _18213_/X sky130_fd_sc_hd__buf_2
XFILLER_54_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15425_ _15333_/X _15422_/X _15424_/X _13242_/X vssd1 vssd1 vccd1 vccd1 _15430_/A
+ sky130_fd_sc_hd__o211a_1
XPHY_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19193_ _16288_/B _18861_/X _19191_/Y _16788_/A _19192_/X vssd1 vssd1 vccd1 vccd1
+ _19193_/X sky130_fd_sc_hd__o221a_1
XFILLER_169_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18144_ _18144_/A _18144_/B vssd1 vssd1 vccd1 vccd1 _18144_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15356_ _15623_/B vssd1 vssd1 vccd1 vccd1 _16151_/S sky130_fd_sc_hd__buf_2
XFILLER_8_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14307_ _26067_/Q _25872_/Q _14307_/S vssd1 vssd1 vccd1 vccd1 _14307_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18075_ _18040_/X _18056_/X _18074_/X vssd1 vssd1 vccd1 vccd1 _18075_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_156_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15287_ _12704_/A _15278_/X _15286_/X _14709_/A vssd1 vssd1 vccd1 vccd1 _15287_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17026_ _17021_/X _16875_/B _17025_/X input219/X vssd1 vssd1 vccd1 vccd1 _17026_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_236_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14238_ _12904_/C _14485_/B _12869_/X vssd1 vssd1 vccd1 vccd1 _14239_/B sky130_fd_sc_hd__a21oi_1
X_14169_ _26912_/Q _14169_/B vssd1 vssd1 vccd1 vccd1 _14169_/X sky130_fd_sc_hd__or2_1
XFILLER_113_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18977_ _18941_/A _18941_/B _17837_/X vssd1 vssd1 vccd1 vccd1 _18978_/B sky130_fd_sc_hd__o21ai_2
XFILLER_140_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _17807_/A _17927_/Y _18681_/A vssd1 vssd1 vccd1 vccd1 _17928_/X sky130_fd_sc_hd__mux2_1
XFILLER_285_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17859_ _19455_/C _19584_/S _18076_/B vssd1 vssd1 vccd1 vccd1 _17859_/X sky130_fd_sc_hd__or3b_1
XFILLER_282_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20870_ _23788_/A _24004_/B vssd1 vssd1 vccd1 vccd1 _20952_/A sky130_fd_sc_hd__nor2_8
XFILLER_254_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19529_ _19525_/X _18923_/X _19527_/X _19528_/X vssd1 vssd1 vccd1 vccd1 _25645_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22540_ _22632_/B vssd1 vssd1 vccd1 vccd1 _22551_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_210_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22471_ _26212_/Q _22459_/X _22470_/X _22468_/X vssd1 vssd1 vccd1 vccd1 _26260_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24210_ _26960_/Q _24213_/C _24209_/X vssd1 vssd1 vccd1 vccd1 _24210_/Y sky130_fd_sc_hd__a21oi_1
X_21422_ input47/X input82/X _21422_/S vssd1 vssd1 vccd1 vccd1 _21423_/A sky130_fd_sc_hd__mux2_8
X_25190_ _25190_/A vssd1 vssd1 vccd1 vccd1 _25199_/A sky130_fd_sc_hd__clkbuf_2
X_24141_ _24141_/A vssd1 vssd1 vccd1 vccd1 _26936_/D sky130_fd_sc_hd__clkbuf_1
X_21353_ _21552_/A vssd1 vssd1 vccd1 vccd1 _21354_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20304_ _20379_/A _20283_/B _20303_/Y vssd1 vssd1 vccd1 vccd1 _20305_/C sky130_fd_sc_hd__a21o_1
XFILLER_162_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24072_ _26906_/Q _23606_/X _24074_/S vssd1 vssd1 vccd1 vccd1 _24073_/A sky130_fd_sc_hd__mux2_1
X_21284_ _21284_/A vssd1 vssd1 vccd1 vccd1 _21284_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23023_ _23023_/A vssd1 vssd1 vccd1 vccd1 _26482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20235_ _20286_/C _20234_/Y _19926_/X vssd1 vssd1 vccd1 vccd1 _20235_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20166_ _25742_/Q vssd1 vssd1 vccd1 vccd1 _20670_/A sky130_fd_sc_hd__buf_8
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24974_ _24974_/A _24978_/B vssd1 vssd1 vccd1 vccd1 _24974_/Y sky130_fd_sc_hd__nand2_1
X_20097_ _19725_/X _20096_/X _20015_/X vssd1 vssd1 vccd1 vccd1 _20102_/A sky130_fd_sc_hd__a21o_1
XFILLER_258_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26713_ _26905_/CLK _26713_/D vssd1 vssd1 vccd1 vccd1 _26713_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23925_ _23925_/A vssd1 vssd1 vccd1 vccd1 _26840_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_58_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27277_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26644_ _26739_/CLK _26644_/D vssd1 vssd1 vccd1 vccd1 _26644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23856_ _23782_/X _26810_/Q _23858_/S vssd1 vssd1 vccd1 vccd1 _23857_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22807_ _26387_/Q _22730_/X _22811_/S vssd1 vssd1 vccd1 vccd1 _22808_/A sky130_fd_sc_hd__mux2_1
X_26575_ _27317_/CLK _26575_/D vssd1 vssd1 vccd1 vccd1 _26575_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20999_ _20999_/A vssd1 vssd1 vccd1 vccd1 _25870_/D sky130_fd_sc_hd__clkbuf_1
X_23787_ _23787_/A vssd1 vssd1 vccd1 vccd1 _26779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13540_ _13540_/A vssd1 vssd1 vccd1 vccd1 _15843_/A sky130_fd_sc_hd__clkbuf_4
X_25526_ _25985_/CLK _25526_/D vssd1 vssd1 vccd1 vccd1 _25526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22738_ _22738_/A vssd1 vssd1 vccd1 vccd1 _26357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ _26790_/Q _26434_/Q _15408_/A vssd1 vssd1 vccd1 vccd1 _13471_/X sky130_fd_sc_hd__mux2_1
X_22669_ _23712_/A vssd1 vssd1 vccd1 vccd1 _22669_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_240_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25457_ _23776_/X _27323_/Q _25459_/S vssd1 vssd1 vccd1 vccd1 _25458_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15210_ _15210_/A vssd1 vssd1 vccd1 vccd1 _15210_/X sky130_fd_sc_hd__clkbuf_4
X_24408_ _24408_/A _24569_/A vssd1 vssd1 vccd1 vccd1 _24408_/Y sky130_fd_sc_hd__nand2_1
X_16190_ _26929_/Q _16262_/S vssd1 vssd1 vccd1 vccd1 _16190_/X sky130_fd_sc_hd__or2_1
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25388_ _25388_/A vssd1 vssd1 vccd1 vccd1 _27292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_275_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27127_ _27130_/CLK _27127_/D vssd1 vssd1 vccd1 vccd1 _27127_/Q sky130_fd_sc_hd__dfxtp_4
X_15141_ _15141_/A vssd1 vssd1 vccd1 vccd1 _15142_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_181_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24339_ _25489_/Q _21208_/B _24340_/S vssd1 vssd1 vccd1 vccd1 _24341_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15072_ _15043_/X _15070_/X _15071_/X vssd1 vssd1 vccd1 vccd1 _15079_/B sky130_fd_sc_hd__a21oi_4
X_27058_ _27058_/CLK _27058_/D vssd1 vssd1 vccd1 vccd1 _27058_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_126_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18900_ _17967_/X _17918_/X _18364_/X _18682_/A vssd1 vssd1 vccd1 vccd1 _18903_/A
+ sky130_fd_sc_hd__o211a_1
X_14023_ _18428_/S _14023_/B vssd1 vssd1 vccd1 vccd1 _17813_/B sky130_fd_sc_hd__or2_4
X_26009_ _27307_/CLK _26009_/D vssd1 vssd1 vccd1 vccd1 _26009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19880_ _17443_/B _19676_/A _19976_/B _19860_/B vssd1 vssd1 vccd1 vccd1 _19889_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_268_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18831_ _25546_/Q _18825_/X _18828_/X _18829_/X _18830_/X vssd1 vssd1 vccd1 vccd1
+ _18831_/X sky130_fd_sc_hd__a221o_1
XFILLER_45_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_14_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_14_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
X_18762_ _27049_/Q _18747_/X _18755_/X _18760_/X _18761_/X vssd1 vssd1 vccd1 vccd1
+ _18762_/X sky130_fd_sc_hd__o221a_2
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15974_ _13065_/A _15971_/X _15973_/X _13142_/A vssd1 vssd1 vccd1 vccd1 _15974_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_212_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17713_ _17738_/A _21208_/A _17712_/Y vssd1 vssd1 vccd1 vccd1 _17753_/A sky130_fd_sc_hd__o21ai_4
XTAP_5583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14925_ _14746_/A _26617_/Q _14905_/S _26357_/Q _14917_/X vssd1 vssd1 vccd1 vccd1
+ _14925_/X sky130_fd_sc_hd__o221a_1
XTAP_5594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18693_ _27080_/Q _18508_/X _18509_/X _27178_/Q _18510_/X vssd1 vssd1 vccd1 vccd1
+ _18693_/X sky130_fd_sc_hd__a221o_1
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ _17650_/A _17644_/B vssd1 vssd1 vccd1 vccd1 _25593_/D sky130_fd_sc_hd__nor2_1
XFILLER_263_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14856_ _14854_/X _14855_/X _14969_/S vssd1 vssd1 vccd1 vccd1 _14856_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13807_ _26071_/Q _25876_/Q _16013_/S vssd1 vssd1 vccd1 vccd1 _13807_/X sky130_fd_sc_hd__mux2_1
XFILLER_223_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17575_ _17575_/A _17575_/B vssd1 vssd1 vccd1 vccd1 _25575_/D sky130_fd_sc_hd__nor2_1
XFILLER_251_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14787_ _16280_/S vssd1 vssd1 vccd1 vccd1 _14787_/X sky130_fd_sc_hd__buf_4
XFILLER_220_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19314_ _25750_/Q vssd1 vssd1 vccd1 vccd1 _19315_/A sky130_fd_sc_hd__buf_8
XFILLER_91_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16526_ _26683_/Q _25723_/Q _16526_/S vssd1 vssd1 vccd1 vccd1 _16526_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13738_ _12892_/A _13561_/A _13736_/X _14029_/B _25926_/Q vssd1 vssd1 vccd1 vccd1
+ _14485_/A sky130_fd_sc_hd__o32a_1
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19245_ _25748_/Q vssd1 vssd1 vccd1 vccd1 _19246_/A sky130_fd_sc_hd__buf_8
XFILLER_32_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16457_ _19325_/A _16567_/B _19327_/A _16456_/X vssd1 vssd1 vccd1 vccd1 _16562_/A
+ sky130_fd_sc_hd__a31o_2
X_13669_ _12738_/D _26693_/Q _26821_/Q _15915_/S _12738_/C vssd1 vssd1 vccd1 vccd1
+ _13669_/X sky130_fd_sc_hd__a221o_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15408_ _15408_/A vssd1 vssd1 vccd1 vccd1 _16194_/S sky130_fd_sc_hd__clkbuf_4
X_19176_ _18740_/X _19174_/Y _19175_/X _19183_/B _18839_/X vssd1 vssd1 vccd1 vccd1
+ _19176_/X sky130_fd_sc_hd__o32a_2
X_16388_ _25896_/Q _16388_/B vssd1 vssd1 vccd1 vccd1 _16388_/X sky130_fd_sc_hd__or2_1
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18127_ _26942_/Q _18569_/A _18570_/A _26974_/Q vssd1 vssd1 vccd1 vccd1 _18127_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15339_ _20252_/A vssd1 vssd1 vccd1 vccd1 _15339_/Y sky130_fd_sc_hd__clkinv_2
X_18058_ _17947_/X _17956_/X _18058_/S vssd1 vssd1 vccd1 vccd1 _18059_/C sky130_fd_sc_hd__mux2_2
XFILLER_117_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17009_ _16784_/X _17008_/X _16862_/B _17006_/X input240/X vssd1 vssd1 vccd1 vccd1
+ _17009_/X sky130_fd_sc_hd__a32o_4
XFILLER_99_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20020_ _20020_/A _20020_/B vssd1 vssd1 vccd1 vccd1 _20020_/Y sky130_fd_sc_hd__nand2_1
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21971_ _21971_/A vssd1 vssd1 vccd1 vccd1 _26099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20922_ _20922_/A vssd1 vssd1 vccd1 vccd1 _25844_/D sky130_fd_sc_hd__clkbuf_1
X_23710_ _23709_/X _26755_/Q _23716_/S vssd1 vssd1 vccd1 vccd1 _23711_/A sky130_fd_sc_hd__mux2_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24690_ _24703_/A _24690_/B vssd1 vssd1 vccd1 vccd1 _24690_/Y sky130_fd_sc_hd__nand2_1
XFILLER_215_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23641_ _26728_/Q _23549_/X _23645_/S vssd1 vssd1 vccd1 vccd1 _23642_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20853_ _20853_/A vssd1 vssd1 vccd1 vccd1 _25822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26360_ _27265_/CLK _26360_/D vssd1 vssd1 vccd1 vccd1 _26360_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_168_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23572_ _26703_/Q _23571_/X _23572_/S vssd1 vssd1 vccd1 vccd1 _23573_/A sky130_fd_sc_hd__mux2_1
X_20784_ _20784_/A vssd1 vssd1 vccd1 vccd1 _25787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_480 _23536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_491 _19268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22523_ _22523_/A vssd1 vssd1 vccd1 vccd1 _26285_/D sky130_fd_sc_hd__clkbuf_1
X_25311_ _23773_/X _27258_/Q _25315_/S vssd1 vssd1 vccd1 vccd1 _25312_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26291_ _26292_/CLK _26291_/D vssd1 vssd1 vccd1 vccd1 _26291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22454_ _26254_/Q _22457_/B vssd1 vssd1 vccd1 vccd1 _22454_/X sky130_fd_sc_hd__or2_1
X_25242_ _27227_/Q _25217_/X _25241_/X _25221_/X vssd1 vssd1 vccd1 vccd1 _27227_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_176_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25596_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21405_ _21402_/X _21404_/X _21367_/X vssd1 vssd1 vccd1 vccd1 _21405_/X sky130_fd_sc_hd__a21o_1
X_25173_ _25173_/A _25198_/A vssd1 vssd1 vccd1 vccd1 _25225_/A sky130_fd_sc_hd__nand2_1
X_22385_ _22393_/A _22406_/A vssd1 vssd1 vccd1 vccd1 _22385_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_105_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26326_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_175_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24124_ _24124_/A vssd1 vssd1 vccd1 vccd1 _26928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21336_ _21407_/A vssd1 vssd1 vccd1 vccd1 _21336_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24055_ _26898_/Q _23581_/X _24059_/S vssd1 vssd1 vccd1 vccd1 _24056_/A sky130_fd_sc_hd__mux2_1
X_21267_ _21265_/X _21266_/X _21289_/A vssd1 vssd1 vccd1 vccd1 _21267_/X sky130_fd_sc_hd__a21o_1
XFILLER_1_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23006_ _26475_/Q _22704_/X _23006_/S vssd1 vssd1 vccd1 vccd1 _23007_/A sky130_fd_sc_hd__mux2_1
XFILLER_277_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20218_ _20218_/A _20218_/B _20218_/C vssd1 vssd1 vccd1 vccd1 _20218_/Y sky130_fd_sc_hd__nor3_2
XFILLER_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21198_ _21198_/A _21870_/B vssd1 vssd1 vccd1 vccd1 _21198_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20149_ _20174_/B _20148_/Y vssd1 vssd1 vccd1 vccd1 _20149_/X sky130_fd_sc_hd__or2b_1
XFILLER_49_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_264_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24957_ _24957_/A vssd1 vssd1 vccd1 vccd1 _24957_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _25499_/Q _25497_/Q _12971_/C vssd1 vssd1 vccd1 vccd1 _12971_/X sky130_fd_sc_hd__or3_2
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14710_ _14710_/A vssd1 vssd1 vccd1 vccd1 _17195_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_261_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23908_ _23908_/A vssd1 vssd1 vccd1 vccd1 _26832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15690_ _15333_/A _15687_/X _15689_/X _14751_/A vssd1 vssd1 vccd1 vccd1 _15694_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24888_ _20696_/A _19724_/X _25155_/A _24782_/X vssd1 vssd1 vccd1 vccd1 _24888_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26627_ _27303_/CLK _26627_/D vssd1 vssd1 vccd1 vccd1 _26627_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _16378_/S vssd1 vssd1 vccd1 vccd1 _14948_/S sky130_fd_sc_hd__buf_2
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23839_ _23757_/X _26802_/Q _23843_/S vssd1 vssd1 vccd1 vccd1 _23840_/A sky130_fd_sc_hd__mux2_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17360_ _25538_/Q _25539_/Q _17360_/C vssd1 vssd1 vccd1 vccd1 _17362_/B sky130_fd_sc_hd__and3_1
X_26558_ _27238_/CLK _26558_/D vssd1 vssd1 vccd1 vccd1 _26558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14572_ _16717_/A _16717_/B _18372_/S vssd1 vssd1 vccd1 vccd1 _16720_/B sky130_fd_sc_hd__o21bai_4
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16311_ _26089_/Q _16399_/S _16144_/S _16310_/X vssd1 vssd1 vccd1 vccd1 _16311_/X
+ sky130_fd_sc_hd__o211a_1
X_13523_ _14047_/A vssd1 vssd1 vccd1 vccd1 _14552_/S sky130_fd_sc_hd__buf_2
X_25509_ _27049_/CLK _25509_/D vssd1 vssd1 vccd1 vccd1 _25509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17291_ _17339_/A vssd1 vssd1 vccd1 vccd1 _17332_/A sky130_fd_sc_hd__buf_2
X_26489_ _27297_/CLK _26489_/D vssd1 vssd1 vccd1 vccd1 _26489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19030_ _18806_/X _19020_/X _19029_/X vssd1 vssd1 vccd1 vccd1 _19030_/X sky130_fd_sc_hd__a21o_4
XFILLER_186_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16242_ _27286_/Q _26479_/Q _16242_/S vssd1 vssd1 vccd1 vccd1 _16242_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13454_ _13436_/X _13453_/X _14590_/A vssd1 vssd1 vccd1 vccd1 _13454_/X sky130_fd_sc_hd__a21o_4
XFILLER_186_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13385_ input125/X input160/X _14132_/S vssd1 vssd1 vccd1 vccd1 _13385_/X sky130_fd_sc_hd__mux2_8
X_16173_ _13255_/A _26897_/Q _26769_/Q _16260_/S _15210_/A vssd1 vssd1 vccd1 vccd1
+ _16173_/X sky130_fd_sc_hd__a221o_1
XFILLER_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15124_ _14759_/A _15120_/X _15123_/X _14779_/A vssd1 vssd1 vccd1 vccd1 _15124_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_182_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15055_ _15053_/X _15054_/X _16224_/S vssd1 vssd1 vccd1 vccd1 _15055_/X sky130_fd_sc_hd__mux2_1
X_19932_ _27142_/Q _19896_/B _19931_/X vssd1 vssd1 vccd1 vccd1 _19933_/C sky130_fd_sc_hd__o21ai_2
XFILLER_126_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14006_ _25803_/Q _13043_/A _14254_/S _14005_/X vssd1 vssd1 vccd1 vccd1 _14006_/X
+ sky130_fd_sc_hd__o211a_1
X_19863_ _27109_/Q _19722_/X _19761_/X _19862_/Y vssd1 vssd1 vccd1 vccd1 _19863_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_268_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18814_ _27212_/Q _19299_/B vssd1 vssd1 vccd1 vccd1 _18814_/X sky130_fd_sc_hd__and2_1
X_19794_ _25666_/Q _19834_/C _20452_/A vssd1 vssd1 vccd1 vccd1 _19794_/X sky130_fd_sc_hd__o21a_1
XFILLER_268_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18745_ _25513_/Q _18743_/X _18744_/X _25545_/Q vssd1 vssd1 vccd1 vccd1 _18745_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15957_ _13558_/A _15955_/X _15956_/Y vssd1 vssd1 vccd1 vccd1 _15957_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput180 irq[3] vssd1 vssd1 vccd1 vccd1 _19624_/C sky130_fd_sc_hd__buf_6
XFILLER_49_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput191 localMemory_wb_adr_i[10] vssd1 vssd1 vccd1 vccd1 input191/X sky130_fd_sc_hd__clkbuf_1
XFILLER_252_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14908_ _26549_/Q _26157_/Q _14991_/S vssd1 vssd1 vccd1 vccd1 _14908_/X sky130_fd_sc_hd__mux2_1
X_18676_ _18686_/A _18676_/B _18635_/A vssd1 vssd1 vccd1 vccd1 _18677_/B sky130_fd_sc_hd__or3b_1
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15888_ _25842_/Q _26042_/Q _15888_/S vssd1 vssd1 vccd1 vccd1 _15889_/B sky130_fd_sc_hd__mux2_1
XFILLER_263_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17627_ _17653_/B vssd1 vssd1 vccd1 vccd1 _17627_/X sky130_fd_sc_hd__buf_2
XFILLER_64_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14839_ _23603_/A vssd1 vssd1 vccd1 vccd1 _14839_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17558_ _17504_/A _17551_/X _17553_/X _17557_/Y vssd1 vssd1 vccd1 vccd1 _17559_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_108_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_3_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26610_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_108_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16509_ _25755_/Q vssd1 vssd1 vccd1 vccd1 _20703_/A sky130_fd_sc_hd__inv_4
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17489_ _26247_/Q _17454_/A _17461_/A _25975_/Q _17488_/X vssd1 vssd1 vccd1 vccd1
+ _17691_/B sky130_fd_sc_hd__a221o_4
XFILLER_60_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19228_ _25557_/Q _18459_/A _19227_/X _17688_/A _18466_/A vssd1 vssd1 vccd1 vccd1
+ _19228_/X sky130_fd_sc_hd__a221o_1
XFILLER_176_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19159_ _18733_/X _19158_/X _15343_/B vssd1 vssd1 vccd1 vccd1 _19159_/X sky130_fd_sc_hd__a21o_1
XFILLER_117_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22170_ _22170_/A vssd1 vssd1 vccd1 vccd1 _22249_/A sky130_fd_sc_hd__buf_2
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21121_ _25914_/Q _21112_/X _21113_/X input13/X vssd1 vssd1 vccd1 vccd1 _21122_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_132_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21052_ _21052_/A vssd1 vssd1 vccd1 vccd1 _25894_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20003_ _20052_/A vssd1 vssd1 vccd1 vccd1 _20003_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_219_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25860_ _26683_/CLK _25860_/D vssd1 vssd1 vccd1 vccd1 _25860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_274_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24811_ _24874_/A vssd1 vssd1 vccd1 vccd1 _24811_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25791_ _25796_/CLK _25791_/D vssd1 vssd1 vccd1 vccd1 _25791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_255_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24742_ _24742_/A _24742_/B vssd1 vssd1 vccd1 vccd1 _27092_/D sky130_fd_sc_hd__nor2_1
X_21954_ _21954_/A vssd1 vssd1 vccd1 vccd1 _26092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20905_ _25839_/Q _20903_/X _20917_/S vssd1 vssd1 vccd1 vccd1 _20906_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21885_ _21885_/A _21885_/B vssd1 vssd1 vccd1 vccd1 _21885_/X sky130_fd_sc_hd__or2_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24673_ _24678_/A _24673_/B vssd1 vssd1 vccd1 vccd1 _27076_/D sky130_fd_sc_hd__nor2_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26412_ _26609_/CLK _26412_/D vssd1 vssd1 vccd1 vccd1 _26412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_270_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23624_ _23624_/A vssd1 vssd1 vccd1 vccd1 _26720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20836_ _25814_/Q vssd1 vssd1 vccd1 vccd1 _20837_/A sky130_fd_sc_hd__clkbuf_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26343_ _27278_/CLK _26343_/D vssd1 vssd1 vccd1 vccd1 _26343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23555_ _23555_/A vssd1 vssd1 vccd1 vccd1 _23555_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20767_ _20767_/A vssd1 vssd1 vccd1 vccd1 _25779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22506_ _22506_/A vssd1 vssd1 vccd1 vccd1 _26277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26274_ _26286_/CLK _26274_/D vssd1 vssd1 vccd1 vccd1 _26274_/Q sky130_fd_sc_hd__dfxtp_1
X_23486_ _23486_/A vssd1 vssd1 vccd1 vccd1 _26673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20698_ _26289_/Q _20686_/X _20696_/Y _20697_/X vssd1 vssd1 vccd1 vccd1 _25752_/D
+ sky130_fd_sc_hd__o211a_1
X_22437_ _26199_/Q _22432_/X _22436_/X _22428_/X vssd1 vssd1 vccd1 vccd1 _26247_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_202_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25225_ _25225_/A vssd1 vssd1 vccd1 vccd1 _25225_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13170_ _12982_/A _13577_/A _13006_/B vssd1 vssd1 vccd1 vccd1 _13171_/A sky130_fd_sc_hd__o21ba_1
XFILLER_164_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22368_ _22368_/A _22368_/B vssd1 vssd1 vccd1 vccd1 _22369_/A sky130_fd_sc_hd__and2_1
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25156_ _27195_/Q _25151_/B _25154_/X _25155_/Y _22380_/X vssd1 vssd1 vccd1 vccd1
+ _27195_/D sky130_fd_sc_hd__o221a_1
XFILLER_272_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21319_ _25941_/Q _21310_/X _21318_/Y _21262_/X vssd1 vssd1 vccd1 vccd1 _25941_/D
+ sky130_fd_sc_hd__a211o_1
X_24107_ _26921_/Q _23552_/X _24109_/S vssd1 vssd1 vccd1 vccd1 _24108_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25087_ _25114_/A vssd1 vssd1 vccd1 vccd1 _25087_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22299_ _22315_/A vssd1 vssd1 vccd1 vccd1 _22299_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_24038_ _24038_/A vssd1 vssd1 vccd1 vccd1 _26890_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27267_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_266_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16860_ _16860_/A _16860_/B vssd1 vssd1 vccd1 vccd1 _16860_/X sky130_fd_sc_hd__and2_2
XFILLER_42_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15811_ _13433_/X _15806_/X _15810_/X _13164_/A vssd1 vssd1 vccd1 vccd1 _15811_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16791_ _16833_/A vssd1 vssd1 vccd1 vccd1 _16982_/B sky130_fd_sc_hd__buf_2
XFILLER_281_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25989_ _27000_/CLK _25989_/D vssd1 vssd1 vccd1 vccd1 _25989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18530_ _25731_/Q _18530_/B vssd1 vssd1 vccd1 vccd1 _18531_/B sky130_fd_sc_hd__nor2_1
XFILLER_246_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15742_ _25884_/Q _15972_/B vssd1 vssd1 vccd1 vccd1 _15742_/X sky130_fd_sc_hd__or2_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12954_ _12953_/A _25479_/Q vssd1 vssd1 vccd1 vccd1 _20485_/A sky130_fd_sc_hd__and2b_2
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _18461_/A vssd1 vssd1 vccd1 vccd1 _18461_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15673_ _15394_/A _15669_/X _15672_/X _13291_/X vssd1 vssd1 vccd1 vccd1 _15673_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_73_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12885_ _13569_/B vssd1 vssd1 vccd1 vccd1 _12941_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _25555_/Q _17410_/B _17411_/Y vssd1 vssd1 vccd1 vccd1 _25555_/D sky130_fd_sc_hd__o21a_1
XFILLER_233_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14624_ _16059_/S vssd1 vssd1 vccd1 vccd1 _16144_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18392_ _18816_/A vssd1 vssd1 vccd1 vccd1 _18509_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_199_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _24966_/A vssd1 vssd1 vccd1 vccd1 _17382_/A sky130_fd_sc_hd__clkbuf_2
X_14555_ _13644_/A _14553_/X _14554_/X _13955_/A vssd1 vssd1 vccd1 vccd1 _14555_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_187_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13506_ _14777_/A _13506_/B _13506_/C vssd1 vssd1 vccd1 vccd1 _13506_/X sky130_fd_sc_hd__or3_1
XFILLER_119_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17274_ _17283_/A _17274_/B _17275_/B vssd1 vssd1 vccd1 vccd1 _25512_/D sky130_fd_sc_hd__nor3_1
XFILLER_186_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14486_ _14486_/A _14486_/B _14486_/C _14485_/Y vssd1 vssd1 vccd1 vccd1 _14486_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_186_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19013_ _19575_/B _16637_/B _19328_/S vssd1 vssd1 vccd1 vccd1 _19013_/X sky130_fd_sc_hd__mux2_1
X_16225_ _26643_/Q _26739_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _16225_/X sky130_fd_sc_hd__mux2_1
X_13437_ _26530_/Q _26138_/Q _13616_/S vssd1 vssd1 vccd1 vccd1 _13437_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16156_ _12773_/A _25850_/Q _26050_/Q _16135_/B vssd1 vssd1 vccd1 vccd1 _16156_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13368_ _15308_/S _13360_/X _13364_/X _13367_/X vssd1 vssd1 vccd1 vccd1 _13369_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_154_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15107_ _16433_/S vssd1 vssd1 vccd1 vccd1 _15119_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_114_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16087_ _26639_/Q _26735_/Q _16087_/S vssd1 vssd1 vccd1 vccd1 _16088_/B sky130_fd_sc_hd__mux2_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13299_ _16193_/S vssd1 vssd1 vccd1 vccd1 _16267_/S sky130_fd_sc_hd__buf_6
XFILLER_138_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19915_ _20650_/A _19698_/X _19913_/X _19914_/X vssd1 vssd1 vccd1 vccd1 _19978_/A
+ sky130_fd_sc_hd__a22oi_4
X_15038_ _26090_/Q _16385_/S _15263_/S _15037_/X vssd1 vssd1 vccd1 vccd1 _15038_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_268_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_256_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19846_ _22487_/A _19845_/B _19738_/X vssd1 vssd1 vccd1 vccd1 _19846_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19777_ _19777_/A _19777_/B vssd1 vssd1 vccd1 vccd1 _19778_/B sky130_fd_sc_hd__nor2_1
X_16989_ _16989_/A vssd1 vssd1 vccd1 vccd1 _16990_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_249_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18728_ _19579_/A _18787_/B _19453_/S vssd1 vssd1 vccd1 vccd1 _18728_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18659_ _27047_/Q _18503_/X _18655_/X _18658_/X _18519_/X vssd1 vssd1 vccd1 vccd1
+ _18659_/X sky130_fd_sc_hd__o221a_1
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21670_ _25975_/Q input210/X _21674_/S vssd1 vssd1 vccd1 vccd1 _21671_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20621_ _23785_/A vssd1 vssd1 vccd1 vccd1 _20621_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23340_ _20580_/X _26609_/Q _23346_/S vssd1 vssd1 vccd1 vccd1 _23341_/A sky130_fd_sc_hd__mux2_1
X_20552_ _20552_/A vssd1 vssd1 vccd1 vccd1 _25706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23271_ _26578_/Q _23121_/X _23277_/S vssd1 vssd1 vccd1 vccd1 _23272_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20483_ _23508_/A vssd1 vssd1 vccd1 vccd1 _23684_/A sky130_fd_sc_hd__buf_2
XFILLER_285_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22222_ _22249_/A vssd1 vssd1 vccd1 vccd1 _22222_/X sky130_fd_sc_hd__buf_2
X_25010_ _16589_/B _25004_/X _25757_/Q _25005_/X vssd1 vssd1 vccd1 vccd1 _25010_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_192_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22153_ _22170_/A vssd1 vssd1 vccd1 vccd1 _22154_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput440 _25944_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[8] sky130_fd_sc_hd__buf_2
XFILLER_133_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput451 _25734_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[10] sky130_fd_sc_hd__buf_2
X_21104_ _21118_/A _21104_/B vssd1 vssd1 vccd1 vccd1 _21105_/A sky130_fd_sc_hd__or2_1
XFILLER_121_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput462 _25744_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[20] sky130_fd_sc_hd__buf_2
X_26961_ _26995_/CLK _26961_/D vssd1 vssd1 vccd1 vccd1 _26961_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput473 _25754_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[30] sky130_fd_sc_hd__buf_2
X_22084_ _26150_/Q _20942_/X _22088_/S vssd1 vssd1 vccd1 vccd1 _22085_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput484 _17052_/X vssd1 vssd1 vccd1 vccd1 wmask0[0] sky130_fd_sc_hd__buf_2
XFILLER_87_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21035_ _25887_/Q _20929_/X _21037_/S vssd1 vssd1 vccd1 vccd1 _21036_/A sky130_fd_sc_hd__mux2_1
X_25912_ _27117_/CLK _25912_/D vssd1 vssd1 vccd1 vccd1 _25912_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_247_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26892_ _27314_/CLK _26892_/D vssd1 vssd1 vccd1 vccd1 _26892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25843_ _26599_/CLK _25843_/D vssd1 vssd1 vccd1 vccd1 _25843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25774_ _26604_/CLK _25774_/D vssd1 vssd1 vccd1 vccd1 _25774_/Q sky130_fd_sc_hd__dfxtp_1
X_22986_ _23032_/S vssd1 vssd1 vccd1 vccd1 _22995_/S sky130_fd_sc_hd__buf_2
XFILLER_170_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24725_ _24725_/A _24725_/B vssd1 vssd1 vccd1 vccd1 _24725_/Y sky130_fd_sc_hd__nand2_4
X_21937_ _21937_/A vssd1 vssd1 vccd1 vccd1 _26084_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _25935_/Q _25934_/Q vssd1 vssd1 vccd1 vccd1 _16641_/A sky130_fd_sc_hd__or2b_2
Xclkbuf_leaf_191_wb_clk_i _26681_/CLK vssd1 vssd1 vccd1 vccd1 _27321_/CLK sky130_fd_sc_hd__clkbuf_16
X_24656_ _24723_/A vssd1 vssd1 vccd1 vccd1 _24678_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_230_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21868_ _21868_/A vssd1 vssd1 vccd1 vccd1 _24455_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23607_ _26714_/Q _23606_/X _23610_/S vssd1 vssd1 vccd1 vccd1 _23608_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_120_wb_clk_i clkbuf_opt_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25985_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20819_ _20819_/A vssd1 vssd1 vccd1 vccd1 _25805_/D sky130_fd_sc_hd__clkbuf_1
X_21799_ _26030_/Q _20875_/X _21805_/S vssd1 vssd1 vccd1 vccd1 _21800_/A sky130_fd_sc_hd__mux2_1
X_24587_ _24944_/A _24595_/B vssd1 vssd1 vccd1 vccd1 _24587_/Y sky130_fd_sc_hd__nand2_1
XFILLER_169_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26326_ _26326_/CLK _26326_/D vssd1 vssd1 vccd1 vccd1 _26326_/Q sky130_fd_sc_hd__dfxtp_1
X_14340_ _14330_/A _14335_/X _14336_/X _14339_/X _13012_/A vssd1 vssd1 vccd1 vccd1
+ _14340_/X sky130_fd_sc_hd__o311a_1
XFILLER_196_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23538_ _23538_/A vssd1 vssd1 vccd1 vccd1 _26692_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26257_ _26257_/CLK _26257_/D vssd1 vssd1 vccd1 vccd1 _26257_/Q sky130_fd_sc_hd__dfxtp_1
X_14271_ _26099_/Q _26000_/Q _14332_/S vssd1 vssd1 vccd1 vccd1 _14271_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23469_ _26666_/Q _23082_/X _23469_/S vssd1 vssd1 vccd1 vccd1 _23470_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16010_ _13834_/A _16008_/X _16009_/X _14077_/A vssd1 vssd1 vccd1 vccd1 _16010_/X
+ sky130_fd_sc_hd__a31o_1
X_13222_ _14060_/A vssd1 vssd1 vccd1 vccd1 _14472_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_183_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25208_ _25208_/A _25208_/B vssd1 vssd1 vccd1 vccd1 _25214_/A sky130_fd_sc_hd__and2_1
X_26188_ _26222_/CLK _26188_/D vssd1 vssd1 vccd1 vccd1 _26188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13153_ _13151_/X _13152_/X _15546_/S vssd1 vssd1 vccd1 vccd1 _13153_/X sky130_fd_sc_hd__mux2_1
X_25139_ _25139_/A vssd1 vssd1 vccd1 vccd1 _25139_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13084_ _13084_/A vssd1 vssd1 vccd1 vccd1 _13085_/A sky130_fd_sc_hd__clkbuf_4
X_17961_ _18896_/A _17961_/B vssd1 vssd1 vccd1 vccd1 _17961_/X sky130_fd_sc_hd__or2_1
XFILLER_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19700_ _19700_/A _19882_/B vssd1 vssd1 vccd1 vccd1 _19700_/Y sky130_fd_sc_hd__nand2_1
X_16912_ _16909_/X _16862_/B _16860_/X _16910_/X _16911_/X vssd1 vssd1 vccd1 vccd1
+ _16912_/X sky130_fd_sc_hd__o221a_1
XFILLER_278_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17892_ _17890_/X _17891_/X _18044_/S vssd1 vssd1 vccd1 vccd1 _17892_/X sky130_fd_sc_hd__mux2_1
XFILLER_239_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16843_ _16836_/X _16840_/Y _16940_/A _16842_/X vssd1 vssd1 vccd1 vccd1 _16844_/B
+ sky130_fd_sc_hd__o211a_4
X_19631_ _25119_/A _19633_/D vssd1 vssd1 vccd1 vccd1 _19640_/A sky130_fd_sc_hd__or2_1
XFILLER_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19562_ _19551_/X _19373_/X _19561_/X _19555_/X vssd1 vssd1 vccd1 vccd1 _25658_/D
+ sky130_fd_sc_hd__o211a_1
X_16774_ _22522_/A _16769_/X _16770_/X _19252_/B vssd1 vssd1 vccd1 vccd1 _16774_/X
+ sky130_fd_sc_hd__a22o_2
X_13986_ _26526_/Q _26134_/Q _14252_/S vssd1 vssd1 vccd1 vccd1 _13986_/X sky130_fd_sc_hd__mux2_1
XFILLER_280_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18513_ _18756_/A vssd1 vssd1 vccd1 vccd1 _18514_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15725_ _26535_/Q _26143_/Q _15725_/S vssd1 vssd1 vccd1 vccd1 _15725_/X sky130_fd_sc_hd__mux2_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19493_ _25632_/Q _19497_/B vssd1 vssd1 vccd1 vccd1 _19493_/X sky130_fd_sc_hd__or2_1
X_12937_ _17592_/B _12937_/B vssd1 vssd1 vccd1 vccd1 _12937_/Y sky130_fd_sc_hd__nor2_1
XFILLER_209_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18444_ _18444_/A vssd1 vssd1 vccd1 vccd1 _18444_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15656_ _14706_/A _15647_/X _15655_/X _14709_/A vssd1 vssd1 vccd1 vccd1 _15656_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_233_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12868_ _12911_/A _12911_/B vssd1 vssd1 vccd1 vccd1 _12868_/Y sky130_fd_sc_hd__nor2_2
XFILLER_61_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _16409_/B _15791_/C vssd1 vssd1 vccd1 vccd1 _14607_/Y sky130_fd_sc_hd__nor2_1
X_18375_ _18552_/A vssd1 vssd1 vccd1 vccd1 _18375_/X sky130_fd_sc_hd__clkbuf_2
X_15587_ _13532_/X _15583_/X _15586_/X _13291_/A vssd1 vssd1 vccd1 vccd1 _15587_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _12799_/A _17129_/A _17133_/A vssd1 vssd1 vccd1 vccd1 _17971_/B sky130_fd_sc_hd__or3_2
X_17326_ _25528_/Q _17324_/B _17325_/Y vssd1 vssd1 vccd1 vccd1 _25528_/D sky130_fd_sc_hd__o21a_1
XFILLER_187_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14538_ _13941_/A _14536_/X _14537_/X _13945_/A vssd1 vssd1 vccd1 vccd1 _14542_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17257_ _25507_/Q _17256_/B _20973_/A vssd1 vssd1 vccd1 vccd1 _17258_/B sky130_fd_sc_hd__o21ai_1
X_14469_ _14453_/X _26685_/Q _26813_/Q _13841_/A _14384_/X vssd1 vssd1 vccd1 vccd1
+ _14469_/X sky130_fd_sc_hd__a221o_1
XFILLER_175_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16208_ _19121_/B vssd1 vssd1 vccd1 vccd1 _19123_/A sky130_fd_sc_hd__clkinv_4
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17188_ _19352_/A vssd1 vssd1 vccd1 vccd1 _17188_/X sky130_fd_sc_hd__buf_2
XFILLER_255_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16139_ _27252_/Q _16243_/B vssd1 vssd1 vccd1 vccd1 _16139_/X sky130_fd_sc_hd__or2_1
XFILLER_89_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19829_ _19829_/A _19855_/A vssd1 vssd1 vccd1 vccd1 _19830_/C sky130_fd_sc_hd__xnor2_2
XFILLER_57_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22840_ _26401_/Q _22672_/X _22840_/S vssd1 vssd1 vccd1 vccd1 _22841_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22771_ _22771_/A vssd1 vssd1 vccd1 vccd1 _26370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24510_ _27030_/Q _24506_/X _24509_/Y _24499_/X vssd1 vssd1 vccd1 vccd1 _27030_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21722_ _21778_/A vssd1 vssd1 vccd1 vccd1 _21791_/S sky130_fd_sc_hd__buf_8
XFILLER_197_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25490_ _25624_/CLK _25490_/D vssd1 vssd1 vccd1 vccd1 _25490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24441_ _24441_/A vssd1 vssd1 vccd1 vccd1 _24551_/A sky130_fd_sc_hd__buf_2
X_21653_ _21651_/Y _21652_/X _21198_/A _17235_/X vssd1 vssd1 vccd1 vccd1 _25968_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_71_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27160_ _27160_/CLK _27160_/D vssd1 vssd1 vccd1 vccd1 _27160_/Q sky130_fd_sc_hd__dfxtp_2
X_20604_ _23597_/A vssd1 vssd1 vccd1 vccd1 _23773_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_21584_ _25961_/Q _21573_/X _21583_/Y _21531_/X vssd1 vssd1 vccd1 vccd1 _25961_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_221_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24372_ _24372_/A _24553_/A vssd1 vssd1 vccd1 vccd1 _24372_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26111_ _26531_/CLK _26111_/D vssd1 vssd1 vccd1 vccd1 _26111_/Q sky130_fd_sc_hd__dfxtp_1
X_23323_ _23323_/A vssd1 vssd1 vccd1 vccd1 _26601_/D sky130_fd_sc_hd__clkbuf_1
X_20535_ _20533_/X _25702_/Q _20551_/S vssd1 vssd1 vccd1 vccd1 _20536_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27091_ _27093_/CLK _27091_/D vssd1 vssd1 vccd1 vccd1 _27091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26042_ _26468_/CLK _26042_/D vssd1 vssd1 vccd1 vccd1 _26042_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_229_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23254_ _23254_/A vssd1 vssd1 vccd1 vccd1 _26570_/D sky130_fd_sc_hd__clkbuf_1
X_20466_ _22533_/A _20467_/C _25691_/Q vssd1 vssd1 vccd1 vccd1 _20466_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22205_ _26185_/Q _22200_/X _22204_/X _22195_/X vssd1 vssd1 vccd1 vccd1 _26185_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23185_ _23196_/A vssd1 vssd1 vccd1 vccd1 _23194_/S sky130_fd_sc_hd__buf_4
X_20397_ _20420_/B _20420_/C _19738_/X vssd1 vssd1 vccd1 vccd1 _20397_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_279_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22136_ _22152_/A vssd1 vssd1 vccd1 vccd1 _22136_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput292 _17070_/X vssd1 vssd1 vccd1 vccd1 addr0[7] sky130_fd_sc_hd__buf_2
XFILLER_88_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26944_ _26980_/CLK _26944_/D vssd1 vssd1 vccd1 vccd1 _26944_/Q sky130_fd_sc_hd__dfxtp_1
X_22067_ _22067_/A vssd1 vssd1 vccd1 vccd1 _26142_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21018_ _25879_/Q _20903_/X _21026_/S vssd1 vssd1 vccd1 vccd1 _21019_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26875_ _26938_/CLK _26875_/D vssd1 vssd1 vccd1 vccd1 _26875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13840_ _26787_/Q _26431_/Q _16013_/S vssd1 vssd1 vccd1 vccd1 _13840_/X sky130_fd_sc_hd__mux2_1
X_25826_ _26744_/CLK _25826_/D vssd1 vssd1 vccd1 vccd1 _25826_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_262_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13771_ _15515_/S vssd1 vssd1 vccd1 vccd1 _15514_/S sky130_fd_sc_hd__clkbuf_4
X_25757_ _26264_/CLK _25757_/D vssd1 vssd1 vccd1 vccd1 _25757_/Q sky130_fd_sc_hd__dfxtp_1
X_22969_ _26458_/Q _22650_/X _22973_/S vssd1 vssd1 vccd1 vccd1 _22970_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_309 _19620_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15510_ _15317_/A _15507_/X _15509_/X _13340_/A vssd1 vssd1 vccd1 vccd1 _15510_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24708_ _27084_/Q _24701_/X _24707_/Y _24697_/X vssd1 vssd1 vccd1 vccd1 _24709_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_12722_ _17738_/B _12722_/B _12722_/C vssd1 vssd1 vccd1 vccd1 _12740_/B sky130_fd_sc_hd__or3_1
X_16490_ _26939_/Q _16490_/B vssd1 vssd1 vccd1 vccd1 _16490_/X sky130_fd_sc_hd__or2_1
X_25688_ _25690_/CLK _25688_/D vssd1 vssd1 vccd1 vccd1 _25688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15441_ _25583_/Q vssd1 vssd1 vccd1 vccd1 _15441_/X sky130_fd_sc_hd__buf_6
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24639_ _24639_/A _12778_/B vssd1 vssd1 vccd1 vccd1 _24639_/X sky130_fd_sc_hd__or2b_1
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18160_ _27201_/Q _18234_/A _18159_/X vssd1 vssd1 vccd1 vccd1 _18160_/X sky130_fd_sc_hd__a21o_1
X_15372_ _25849_/Q _26049_/Q _15374_/S vssd1 vssd1 vccd1 vccd1 _15372_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17111_ _16639_/Y _16645_/X _16647_/X _16648_/X _24986_/A vssd1 vssd1 vccd1 vccd1
+ _25465_/S sky130_fd_sc_hd__o2111a_4
XFILLER_128_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26309_ _26327_/CLK _26309_/D vssd1 vssd1 vccd1 vccd1 _26309_/Q sky130_fd_sc_hd__dfxtp_2
X_14323_ _14323_/A _14323_/B vssd1 vssd1 vccd1 vccd1 _14323_/Y sky130_fd_sc_hd__nand2_1
XFILLER_184_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18091_ _20092_/A vssd1 vssd1 vccd1 vccd1 _18092_/A sky130_fd_sc_hd__buf_2
XFILLER_128_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27289_ _27292_/CLK _27289_/D vssd1 vssd1 vccd1 vccd1 _27289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17042_ _17042_/A vssd1 vssd1 vccd1 vccd1 _17042_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14254_ _14252_/X _14253_/X _14254_/S vssd1 vssd1 vccd1 vccd1 _14254_/X sky130_fd_sc_hd__mux2_1
X_13205_ _13464_/A vssd1 vssd1 vccd1 vccd1 _13638_/A sky130_fd_sc_hd__clkbuf_8
X_14185_ _13172_/A _14184_/X _13026_/A vssd1 vssd1 vccd1 vccd1 _14185_/X sky130_fd_sc_hd__o21a_1
XFILLER_152_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13136_ _13723_/A vssd1 vssd1 vccd1 vccd1 _16059_/S sky130_fd_sc_hd__buf_4
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ _17395_/X _18763_/X _18992_/X _18767_/X _18768_/X vssd1 vssd1 vccd1 vccd1
+ _18993_/X sky130_fd_sc_hd__a221o_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _13053_/X _13061_/X _15567_/S vssd1 vssd1 vccd1 vccd1 _13067_/X sky130_fd_sc_hd__mux2_1
X_17944_ _17932_/X _17940_/X _18489_/S vssd1 vssd1 vccd1 vccd1 _17944_/X sky130_fd_sc_hd__mux2_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17875_ _17797_/B _17782_/B _17954_/S vssd1 vssd1 vccd1 vccd1 _17875_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19614_ _19614_/A _19614_/B _19614_/C _19614_/D vssd1 vssd1 vccd1 vccd1 _19628_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_38_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16826_ _16826_/A vssd1 vssd1 vccd1 vccd1 _16895_/A sky130_fd_sc_hd__buf_2
XFILLER_171_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19545_ _25652_/Q _19549_/B vssd1 vssd1 vccd1 vccd1 _19545_/X sky130_fd_sc_hd__or2_1
X_16757_ _16770_/A vssd1 vssd1 vccd1 vccd1 _16757_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_281_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13969_ _13967_/X _13968_/X _14309_/S vssd1 vssd1 vccd1 vccd1 _13969_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15708_ _15708_/A _15708_/B vssd1 vssd1 vccd1 vccd1 _15708_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19476_ _18895_/X _19460_/X _19475_/X _18927_/X vssd1 vssd1 vccd1 vccd1 _19476_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16688_ _25756_/Q _20800_/B vssd1 vssd1 vccd1 vccd1 _16689_/A sky130_fd_sc_hd__and2_2
XFILLER_250_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18427_ _18898_/A _18426_/Y _17988_/X vssd1 vssd1 vccd1 vccd1 _18427_/X sky130_fd_sc_hd__a21bo_1
X_15639_ _14621_/A _15625_/X _15629_/X _15638_/X _14682_/A vssd1 vssd1 vccd1 vccd1
+ _15639_/X sky130_fd_sc_hd__a311o_1
XFILLER_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18358_ _18358_/A vssd1 vssd1 vccd1 vccd1 _18636_/A sky130_fd_sc_hd__clkbuf_2
X_17309_ _17308_/X _17312_/C _17269_/X vssd1 vssd1 vccd1 vccd1 _17309_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18289_ _18339_/A _18329_/A vssd1 vssd1 vccd1 vccd1 _18289_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20320_ _27157_/Q _27091_/Q vssd1 vssd1 vccd1 vccd1 _20320_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20251_ _20251_/A vssd1 vssd1 vccd1 vccd1 _20251_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20182_ _20180_/Y _20182_/B vssd1 vssd1 vccd1 vccd1 _20184_/A sky130_fd_sc_hd__and2b_1
XFILLER_115_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24990_ _24989_/X _24544_/B _20276_/A vssd1 vssd1 vccd1 vccd1 _24994_/B sky130_fd_sc_hd__o21a_1
XFILLER_229_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23941_ _26847_/Q _23520_/X _23943_/S vssd1 vssd1 vccd1 vccd1 _23942_/A sky130_fd_sc_hd__mux2_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26660_ _26916_/CLK _26660_/D vssd1 vssd1 vccd1 vccd1 _26660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23872_ _23872_/A vssd1 vssd1 vccd1 vccd1 _26816_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25611_ _25660_/CLK _25611_/D vssd1 vssd1 vccd1 vccd1 _25611_/Q sky130_fd_sc_hd__dfxtp_2
X_22823_ _26393_/Q _22647_/X _22829_/S vssd1 vssd1 vccd1 vccd1 _22824_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26591_ _26592_/CLK _26591_/D vssd1 vssd1 vccd1 vccd1 _26591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25542_ _25545_/CLK _25542_/D vssd1 vssd1 vccd1 vccd1 _25542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22754_ _26363_/Q _22653_/X _22756_/S vssd1 vssd1 vccd1 vccd1 _22755_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21705_ _25991_/Q _17456_/C _21707_/S vssd1 vssd1 vccd1 vccd1 _21706_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25473_ _25598_/CLK _25473_/D vssd1 vssd1 vccd1 vccd1 _25473_/Q sky130_fd_sc_hd__dfxtp_2
X_22685_ _23728_/A vssd1 vssd1 vccd1 vccd1 _22685_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_241_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27212_ _27213_/CLK _27212_/D vssd1 vssd1 vccd1 vccd1 _27212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24424_ _24686_/B vssd1 vssd1 vccd1 vccd1 _24577_/A sky130_fd_sc_hd__clkinv_2
XFILLER_185_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21636_ _21636_/A vssd1 vssd1 vccd1 vccd1 _21636_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27143_ _27166_/CLK _27143_/D vssd1 vssd1 vccd1 vccd1 _27143_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_139_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24355_ _25206_/B _24776_/C vssd1 vssd1 vccd1 vccd1 _24390_/A sky130_fd_sc_hd__nor2b_2
XFILLER_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21567_ _25866_/Q vssd1 vssd1 vccd1 vccd1 _21615_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_154_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23306_ _23306_/A vssd1 vssd1 vccd1 vccd1 _26593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20518_ _20517_/X _25698_/Q _20530_/S vssd1 vssd1 vccd1 vccd1 _20519_/A sky130_fd_sc_hd__mux2_1
X_27074_ _27203_/CLK _27074_/D vssd1 vssd1 vccd1 vccd1 _27074_/Q sky130_fd_sc_hd__dfxtp_2
X_24286_ _26986_/Q _24286_/B vssd1 vssd1 vccd1 vccd1 _24293_/C sky130_fd_sc_hd__and2_1
XFILLER_197_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21498_ _20675_/A _21481_/X _21459_/X _21497_/X vssd1 vssd1 vccd1 vccd1 _21498_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26025_ _26580_/CLK _26025_/D vssd1 vssd1 vccd1 vccd1 _26025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23237_ _23237_/A vssd1 vssd1 vccd1 vccd1 _26562_/D sky130_fd_sc_hd__clkbuf_1
X_20449_ _20471_/A _20449_/B vssd1 vssd1 vccd1 vccd1 _20450_/C sky130_fd_sc_hd__nand2_1
XFILLER_107_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23168_ _26532_/Q _23076_/X _23172_/S vssd1 vssd1 vccd1 vccd1 _23169_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22119_ input188/X _22113_/X _22115_/X _17085_/A _22118_/X vssd1 vssd1 vccd1 vccd1
+ _22119_/X sky130_fd_sc_hd__a221o_1
XFILLER_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15990_ _15988_/X _15989_/X _15990_/S vssd1 vssd1 vccd1 vccd1 _15990_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23099_ _26507_/Q _23098_/X _23099_/S vssd1 vssd1 vccd1 vccd1 _23100_/A sky130_fd_sc_hd__mux2_1
XFILLER_279_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14941_ _23600_/A vssd1 vssd1 vccd1 vccd1 _14941_/Y sky130_fd_sc_hd__inv_2
X_26927_ _27311_/CLK _26927_/D vssd1 vssd1 vccd1 vccd1 _26927_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17660_ _18338_/A vssd1 vssd1 vccd1 vccd1 _18336_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26858_ _27278_/CLK _26858_/D vssd1 vssd1 vccd1 vccd1 _26858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14872_ _16224_/S vssd1 vssd1 vccd1 vccd1 _14877_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_275_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16611_ _19121_/A _19123_/A vssd1 vssd1 vccd1 vccd1 _16638_/B sky130_fd_sc_hd__xnor2_4
X_13823_ _13472_/A _26691_/Q _26819_/Q _15758_/S _13821_/A vssd1 vssd1 vccd1 vccd1
+ _13823_/X sky130_fd_sc_hd__a221o_1
X_25809_ _26917_/CLK _25809_/D vssd1 vssd1 vccd1 vccd1 _25809_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_63_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17591_ _17595_/A _17591_/B vssd1 vssd1 vccd1 vccd1 _25579_/D sky130_fd_sc_hd__nor2_1
X_26789_ _27304_/CLK _26789_/D vssd1 vssd1 vccd1 vccd1 _26789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_106 _21616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_117 _23032_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19330_ _25528_/Q _18556_/X _18557_/X _25560_/Q vssd1 vssd1 vccd1 vccd1 _19330_/X
+ sky130_fd_sc_hd__a22o_1
X_16542_ _16513_/X _26619_/Q _16523_/S _26359_/Q _16540_/S vssd1 vssd1 vccd1 vccd1
+ _16542_/X sky130_fd_sc_hd__o221a_1
X_13754_ _13011_/A _13735_/Y _13753_/Y vssd1 vssd1 vccd1 vccd1 _16839_/A sky130_fd_sc_hd__a21oi_4
XINSDIODE2_128 _20189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_139 _13808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19261_ _27158_/Q _19261_/B vssd1 vssd1 vccd1 vccd1 _19261_/X sky130_fd_sc_hd__or2_1
X_12705_ _12705_/A vssd1 vssd1 vccd1 vccd1 _12706_/A sky130_fd_sc_hd__buf_4
XFILLER_232_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16473_ _26551_/Q _26159_/Q _16498_/S vssd1 vssd1 vccd1 vccd1 _16473_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13685_ _25733_/Q _16031_/S vssd1 vssd1 vccd1 vccd1 _13685_/X sky130_fd_sc_hd__or2_2
X_18212_ _18205_/X _18211_/X _18799_/A vssd1 vssd1 vccd1 vccd1 _18212_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15424_ _15424_/A _15424_/B vssd1 vssd1 vccd1 vccd1 _15424_/X sky130_fd_sc_hd__or2_1
XPHY_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19192_ _19192_/A _19192_/B vssd1 vssd1 vccd1 vccd1 _19192_/X sky130_fd_sc_hd__or2_1
XPHY_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18143_ _18027_/X _18032_/Y _18142_/X _18976_/A vssd1 vssd1 vccd1 vccd1 _18144_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_15355_ _15555_/S vssd1 vssd1 vccd1 vccd1 _15623_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_12_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14306_ _15760_/A _14302_/X _14305_/X _13529_/A vssd1 vssd1 vccd1 vccd1 _14306_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18074_ _18896_/A _18065_/X _18073_/X _18343_/A vssd1 vssd1 vccd1 vccd1 _18074_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15286_ _15285_/A _15281_/X _15285_/Y _15187_/X vssd1 vssd1 vccd1 vccd1 _15286_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17025_ _17039_/A vssd1 vssd1 vccd1 vccd1 _17025_/X sky130_fd_sc_hd__clkbuf_2
X_14237_ _14237_/A _14237_/B _14237_/C _14237_/D vssd1 vssd1 vccd1 vccd1 _14237_/Y
+ sky130_fd_sc_hd__nor4_1
XFILLER_153_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14168_ _27299_/Q _26556_/Q _15714_/A vssd1 vssd1 vccd1 vccd1 _14168_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13119_ _26919_/Q _15561_/B vssd1 vssd1 vccd1 vccd1 _13119_/X sky130_fd_sc_hd__or2_1
XFILLER_285_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14099_ _14165_/A _14098_/Y _13630_/A vssd1 vssd1 vccd1 vccd1 _14099_/Y sky130_fd_sc_hd__a21oi_1
X_18976_ _18976_/A vssd1 vssd1 vccd1 vccd1 _18976_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_252_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _17927_/A vssd1 vssd1 vccd1 vccd1 _17927_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17858_ _17857_/Y _19452_/B _16551_/B vssd1 vssd1 vccd1 vccd1 _19584_/S sky130_fd_sc_hd__a21o_1
XFILLER_226_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16809_ _16982_/B _16809_/B _16809_/C vssd1 vssd1 vccd1 vccd1 _16841_/B sky130_fd_sc_hd__and3_4
X_17789_ _19327_/A _17789_/B vssd1 vssd1 vccd1 vccd1 _19355_/B sky130_fd_sc_hd__or2_1
XFILLER_53_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19528_ _19541_/A vssd1 vssd1 vccd1 vccd1 _19528_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_207_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19459_ _18342_/A _17989_/Y _19458_/X _18738_/A vssd1 vssd1 vccd1 vccd1 _19459_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22470_ _26260_/Q _22470_/B vssd1 vssd1 vccd1 vccd1 _22470_/X sky130_fd_sc_hd__or2_1
XFILLER_195_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21421_ _21552_/A vssd1 vssd1 vccd1 vccd1 _21421_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21352_ _21342_/X _21351_/X _21336_/X vssd1 vssd1 vccd1 vccd1 _21352_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_148_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24140_ _26936_/Q _23600_/X _24142_/S vssd1 vssd1 vccd1 vccd1 _24141_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20303_ _20359_/A _20303_/B vssd1 vssd1 vccd1 vccd1 _20303_/Y sky130_fd_sc_hd__nor2_1
XFILLER_163_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21283_ _21283_/A vssd1 vssd1 vccd1 vccd1 _21284_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_24071_ _24071_/A vssd1 vssd1 vccd1 vccd1 _26905_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20234_ _25680_/Q _20233_/C _22516_/A vssd1 vssd1 vccd1 vccd1 _20234_/Y sky130_fd_sc_hd__a21oi_1
X_23022_ _26482_/Q _22727_/X _23028_/S vssd1 vssd1 vccd1 vccd1 _23023_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20165_ _22511_/A _20164_/B _19738_/X vssd1 vssd1 vccd1 vccd1 _20165_/Y sky130_fd_sc_hd__o21ai_1
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24973_ _27158_/Q _24953_/X _24972_/Y _24970_/X vssd1 vssd1 vccd1 vccd1 _27158_/D
+ sky130_fd_sc_hd__o211a_1
X_20096_ _20205_/B _20204_/A vssd1 vssd1 vccd1 vccd1 _20096_/X sky130_fd_sc_hd__xor2_1
XFILLER_58_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26712_ _26904_/CLK _26712_/D vssd1 vssd1 vccd1 vccd1 _26712_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23924_ _23776_/X _26840_/Q _23926_/S vssd1 vssd1 vccd1 vccd1 _23925_/A sky130_fd_sc_hd__mux2_1
XFILLER_273_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26643_ _26739_/CLK _26643_/D vssd1 vssd1 vccd1 vccd1 _26643_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23855_ _23855_/A vssd1 vssd1 vccd1 vccd1 _26809_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22806_ _22806_/A vssd1 vssd1 vccd1 vccd1 _26386_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26574_ _27317_/CLK _26574_/D vssd1 vssd1 vccd1 vccd1 _26574_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23786_ _23785_/X _26779_/Q _23786_/S vssd1 vssd1 vccd1 vccd1 _23787_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20998_ _25870_/Q _20875_/X _21004_/S vssd1 vssd1 vccd1 vccd1 _20999_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25525_ _25985_/CLK _25525_/D vssd1 vssd1 vccd1 vccd1 _25525_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_98_wb_clk_i clkbuf_4_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26240_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_164_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22737_ _26357_/Q _22736_/X _22737_/S vssd1 vssd1 vccd1 vccd1 _22738_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13470_ _15768_/S vssd1 vssd1 vccd1 vccd1 _15408_/A sky130_fd_sc_hd__buf_4
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25456_ _25456_/A vssd1 vssd1 vccd1 vccd1 _27322_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_27_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26939_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22668_ _22668_/A vssd1 vssd1 vccd1 vccd1 _26335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24407_ _24671_/B vssd1 vssd1 vccd1 vccd1 _24569_/A sky130_fd_sc_hd__clkinv_2
XFILLER_139_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21619_ _25964_/Q _21573_/X _21618_/Y _21597_/X vssd1 vssd1 vccd1 vccd1 _25964_/D
+ sky130_fd_sc_hd__a211o_1
X_25387_ _27292_/Q _23779_/A _25387_/S vssd1 vssd1 vccd1 vccd1 _25388_/A sky130_fd_sc_hd__mux2_1
X_22599_ _26315_/Q _22604_/B vssd1 vssd1 vccd1 vccd1 _22599_/Y sky130_fd_sc_hd__nand2_1
XFILLER_194_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15140_ _27319_/Q _26576_/Q _16387_/S vssd1 vssd1 vccd1 vccd1 _15140_/X sky130_fd_sc_hd__mux2_1
X_27126_ _27130_/CLK _27126_/D vssd1 vssd1 vccd1 vccd1 _27126_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24338_ _27004_/Q _24335_/B _24337_/Y vssd1 vssd1 vccd1 vccd1 _27004_/D sky130_fd_sc_hd__o21a_1
XFILLER_166_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27057_ _27062_/CLK _27057_/D vssd1 vssd1 vccd1 vccd1 _27057_/Q sky130_fd_sc_hd__dfxtp_2
X_15071_ _15071_/A vssd1 vssd1 vccd1 vccd1 _15071_/X sky130_fd_sc_hd__buf_4
X_24269_ _24269_/A _24275_/C vssd1 vssd1 vccd1 vccd1 _24269_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26008_ _26599_/CLK _26008_/D vssd1 vssd1 vccd1 vccd1 _26008_/Q sky130_fd_sc_hd__dfxtp_2
X_14022_ _14022_/A _17798_/A vssd1 vssd1 vccd1 vccd1 _14023_/B sky130_fd_sc_hd__nor2_1
XFILLER_106_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18830_ _18830_/A vssd1 vssd1 vccd1 vccd1 _18830_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15973_ _26076_/Q _15961_/B _14010_/S _15972_/X vssd1 vssd1 vccd1 vccd1 _15973_/X
+ sky130_fd_sc_hd__o211a_1
X_18761_ _18823_/A vssd1 vssd1 vccd1 vccd1 _18761_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_283_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17712_ _17738_/A _17712_/B vssd1 vssd1 vccd1 vccd1 _17712_/Y sky130_fd_sc_hd__nand2_1
X_14924_ _26517_/Q _26389_/Q _15005_/S vssd1 vssd1 vccd1 vccd1 _14924_/X sky130_fd_sc_hd__mux2_1
XTAP_5584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18692_ _27210_/Q _19258_/B vssd1 vssd1 vccd1 vccd1 _18692_/X sky130_fd_sc_hd__and2_1
XTAP_5595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14855_ _26517_/Q _26389_/Q _14876_/S vssd1 vssd1 vccd1 vccd1 _14855_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17643_ _17443_/B _17635_/X _17608_/A _17642_/Y vssd1 vssd1 vccd1 vccd1 _17644_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13806_ _15999_/A vssd1 vssd1 vccd1 vccd1 _13806_/X sky130_fd_sc_hd__buf_4
XFILLER_205_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17574_ _25575_/Q _17564_/X _17572_/X _17573_/X vssd1 vssd1 vccd1 vccd1 _17575_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_205_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14786_ _14786_/A vssd1 vssd1 vccd1 vccd1 _16280_/S sky130_fd_sc_hd__buf_2
XFILLER_223_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19313_ _18220_/X _19297_/X _19312_/X _18841_/X vssd1 vssd1 vccd1 vccd1 _19313_/X
+ sky130_fd_sc_hd__a22o_1
X_16525_ _16522_/X _16523_/X _16540_/S vssd1 vssd1 vccd1 vccd1 _16525_/X sky130_fd_sc_hd__mux2_1
X_13737_ _13737_/A vssd1 vssd1 vccd1 vccd1 _14029_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16456_ _19322_/A _19294_/S _16454_/B vssd1 vssd1 vccd1 vccd1 _16456_/X sky130_fd_sc_hd__o21ba_1
X_19244_ _18841_/X _19219_/Y _19234_/X _19243_/X _18375_/X vssd1 vssd1 vccd1 vccd1
+ _19244_/X sky130_fd_sc_hd__a32o_1
X_13668_ _26629_/Q _26725_/Q _15842_/S vssd1 vssd1 vccd1 vccd1 _13668_/X sky130_fd_sc_hd__mux2_1
X_15407_ _15406_/X _26348_/Q _26608_/Q _16443_/S _15417_/A vssd1 vssd1 vccd1 vccd1
+ _15407_/X sky130_fd_sc_hd__a221o_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19175_ _18947_/A _19173_/Y _18998_/X vssd1 vssd1 vccd1 vccd1 _19175_/X sky130_fd_sc_hd__o21a_1
X_16387_ _27290_/Q _26483_/Q _16387_/S vssd1 vssd1 vccd1 vccd1 _16387_/X sky130_fd_sc_hd__mux2_1
X_13599_ _14169_/B vssd1 vssd1 vccd1 vccd1 _14008_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_118_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18126_ _18462_/A vssd1 vssd1 vccd1 vccd1 _18570_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_247_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15338_ _14723_/A _15250_/Y _15337_/Y _14827_/A vssd1 vssd1 vccd1 vccd1 _20252_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_8_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18057_ _17950_/X _17946_/X _18063_/S vssd1 vssd1 vccd1 vccd1 _18057_/X sky130_fd_sc_hd__mux2_1
X_15269_ _14649_/A _15263_/X _15268_/X _14679_/A vssd1 vssd1 vccd1 vccd1 _15269_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_160_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17008_ _17042_/A vssd1 vssd1 vccd1 vccd1 _17008_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18959_ _18435_/A _18958_/X _18947_/B vssd1 vssd1 vccd1 vccd1 _18959_/X sky130_fd_sc_hd__a21o_1
XFILLER_239_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21970_ _26099_/Q _20881_/X _21972_/S vssd1 vssd1 vccd1 vccd1 _21971_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20921_ _25844_/Q _20919_/X _20933_/S vssd1 vssd1 vccd1 vccd1 _20922_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23640_ _23640_/A vssd1 vssd1 vccd1 vccd1 _26727_/D sky130_fd_sc_hd__clkbuf_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20852_ _25822_/Q vssd1 vssd1 vccd1 vccd1 _20853_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23571_ _23571_/A vssd1 vssd1 vccd1 vccd1 _23571_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_211_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20783_ _20613_/X _25787_/Q _20783_/S vssd1 vssd1 vccd1 vccd1 _20784_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_470 _23702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25310_ _25310_/A vssd1 vssd1 vccd1 vccd1 _27257_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_481 _19849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22522_ _22522_/A _22524_/B vssd1 vssd1 vccd1 vccd1 _22523_/A sky130_fd_sc_hd__and2_1
XFILLER_50_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26290_ _26292_/CLK _26290_/D vssd1 vssd1 vccd1 vccd1 _26290_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_492 _16414_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25241_ _25208_/A _19614_/B _24771_/A _24762_/B _25219_/X vssd1 vssd1 vccd1 vccd1
+ _25241_/X sky130_fd_sc_hd__a221o_1
X_22453_ _26205_/Q _22446_/X _22452_/X _22442_/X vssd1 vssd1 vccd1 vccd1 _26253_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21404_ _21364_/X _18772_/X _21365_/X _25809_/Q _21403_/X vssd1 vssd1 vccd1 vccd1
+ _21404_/X sky130_fd_sc_hd__a221o_1
X_25172_ _25198_/A vssd1 vssd1 vccd1 vccd1 _25172_/X sky130_fd_sc_hd__clkbuf_2
X_22384_ _26237_/Q vssd1 vssd1 vccd1 vccd1 _22406_/A sky130_fd_sc_hd__inv_2
XFILLER_175_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24123_ _26928_/Q _23574_/X _24131_/S vssd1 vssd1 vccd1 vccd1 _24124_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21335_ _20641_/A _21278_/X _21279_/X _21334_/X vssd1 vssd1 vccd1 vccd1 _21335_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24054_ _24054_/A vssd1 vssd1 vccd1 vccd1 _26897_/D sky130_fd_sc_hd__clkbuf_1
X_21266_ _21283_/A _18177_/X _21285_/A _25799_/Q _21346_/A vssd1 vssd1 vccd1 vccd1
+ _21266_/X sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_145_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25624_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_235_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23005_ _23005_/A vssd1 vssd1 vccd1 vccd1 _26474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20217_ _20218_/A _20218_/B _20218_/C vssd1 vssd1 vccd1 vccd1 _20217_/X sky130_fd_sc_hd__o21a_1
XFILLER_235_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21197_ _21197_/A _21197_/B vssd1 vssd1 vccd1 vccd1 _25935_/D sky130_fd_sc_hd__nor2_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20148_ _20200_/A _20148_/B vssd1 vssd1 vccd1 vccd1 _20148_/Y sky130_fd_sc_hd__nand2_1
XFILLER_265_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_253_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24956_ _27151_/Q _24953_/X _24955_/Y _24949_/X vssd1 vssd1 vccd1 vccd1 _27151_/D
+ sky130_fd_sc_hd__o211a_1
X_12970_ _25496_/Q _25495_/Q _25494_/Q _25493_/Q vssd1 vssd1 vccd1 vccd1 _12971_/C
+ sky130_fd_sc_hd__or4_1
X_20079_ _20079_/A vssd1 vssd1 vccd1 vccd1 _20079_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_218_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23907_ _23750_/X _26832_/Q _23915_/S vssd1 vssd1 vccd1 vccd1 _23908_/A sky130_fd_sc_hd__mux2_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24887_ _27129_/Q _24890_/B vssd1 vssd1 vccd1 vccd1 _24887_/Y sky130_fd_sc_hd__nand2_1
XFILLER_261_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26626_ _27301_/CLK _26626_/D vssd1 vssd1 vccd1 vccd1 _26626_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _16324_/S vssd1 vssd1 vccd1 vccd1 _16378_/S sky130_fd_sc_hd__buf_2
XFILLER_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23838_ _23838_/A vssd1 vssd1 vccd1 vccd1 _26801_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26557_ _26877_/CLK _26557_/D vssd1 vssd1 vccd1 vccd1 _26557_/Q sky130_fd_sc_hd__dfxtp_1
X_14571_ _18324_/B _16713_/A _16713_/B _14570_/Y vssd1 vssd1 vccd1 vccd1 _16717_/B
+ sky130_fd_sc_hd__o31a_2
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23769_ _23769_/A vssd1 vssd1 vccd1 vccd1 _26773_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16310_ _25894_/Q _16310_/B vssd1 vssd1 vccd1 vccd1 _16310_/X sky130_fd_sc_hd__or2_1
XFILLER_241_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13522_ _15490_/A vssd1 vssd1 vccd1 vccd1 _15488_/A sky130_fd_sc_hd__buf_2
X_25508_ _27049_/CLK _25508_/D vssd1 vssd1 vccd1 vccd1 _25508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17290_ _25109_/A vssd1 vssd1 vccd1 vccd1 _17339_/A sky130_fd_sc_hd__buf_6
X_26488_ _26520_/CLK _26488_/D vssd1 vssd1 vccd1 vccd1 _26488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16241_ _16239_/X _16240_/X _16241_/S vssd1 vssd1 vccd1 vccd1 _16241_/X sky130_fd_sc_hd__mux2_1
X_13453_ _12702_/A _13444_/X _13452_/X _13717_/A vssd1 vssd1 vccd1 vccd1 _13453_/X
+ sky130_fd_sc_hd__a211o_1
X_25439_ _25450_/A vssd1 vssd1 vccd1 vccd1 _25448_/S sky130_fd_sc_hd__buf_4
XFILLER_40_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16172_ _26673_/Q _25713_/Q _16194_/S vssd1 vssd1 vccd1 vccd1 _16172_/X sky130_fd_sc_hd__mux2_1
X_13384_ _14033_/S vssd1 vssd1 vccd1 vccd1 _14132_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_154_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15123_ _14765_/A _15121_/X _15122_/X _12756_/A vssd1 vssd1 vccd1 vccd1 _15123_/X
+ sky130_fd_sc_hd__o211a_1
X_27109_ _27110_/CLK _27109_/D vssd1 vssd1 vccd1 vccd1 _27109_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15054_ _26122_/Q _26023_/Q _16380_/B vssd1 vssd1 vccd1 vccd1 _15054_/X sky130_fd_sc_hd__mux2_1
X_19931_ _27142_/Q _27076_/Q _19898_/Y vssd1 vssd1 vccd1 vccd1 _19931_/X sky130_fd_sc_hd__a21o_1
XFILLER_126_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14005_ _27237_/Q _15808_/B vssd1 vssd1 vccd1 vccd1 _14005_/X sky130_fd_sc_hd__or2_1
X_19862_ _19906_/C _19846_/Y _19765_/X _19861_/X vssd1 vssd1 vccd1 vccd1 _19862_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_68_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_269_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18813_ _18813_/A vssd1 vssd1 vccd1 vccd1 _19299_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_233_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19793_ _22483_/A _19834_/C vssd1 vssd1 vccd1 vccd1 _19793_/Y sky130_fd_sc_hd__nand2_1
XFILLER_284_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18744_ _18808_/A vssd1 vssd1 vccd1 vccd1 _18744_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_209_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15956_ _25642_/Q _13803_/B _14611_/A vssd1 vssd1 vccd1 vccd1 _15956_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput170 dout1[9] vssd1 vssd1 vccd1 vccd1 input170/X sky130_fd_sc_hd__clkbuf_1
XTAP_5392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput181 irq[4] vssd1 vssd1 vccd1 vccd1 _19609_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_76_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput192 localMemory_wb_adr_i[11] vssd1 vssd1 vccd1 vccd1 input192/X sky130_fd_sc_hd__clkbuf_1
X_14907_ _14765_/A _14905_/X _14906_/X _12757_/A vssd1 vssd1 vccd1 vccd1 _14907_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_236_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15887_ _15990_/S _15887_/B vssd1 vssd1 vccd1 vccd1 _15887_/X sky130_fd_sc_hd__or2_1
X_18675_ _17822_/Y _18635_/A _18686_/A vssd1 vssd1 vccd1 vccd1 _18724_/B sky130_fd_sc_hd__a21boi_1
XFILLER_270_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17626_ _17633_/A _17626_/B vssd1 vssd1 vccd1 vccd1 _25588_/D sky130_fd_sc_hd__nor2_1
XFILLER_24_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14838_ _25627_/Q _14597_/X _14837_/X _14618_/X vssd1 vssd1 vccd1 vccd1 _23603_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_17_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17557_ _25908_/Q _17554_/X _17556_/X vssd1 vssd1 vccd1 vccd1 _17557_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14769_ _15210_/A vssd1 vssd1 vccd1 vccd1 _14770_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_251_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16508_ _20189_/A _16982_/C _16508_/S vssd1 vssd1 vccd1 vccd1 _16550_/A sky130_fd_sc_hd__mux2_1
X_17488_ _26248_/Q _17453_/A _17460_/A _25976_/Q vssd1 vssd1 vccd1 vccd1 _17488_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19227_ _26965_/Q _18461_/A _18463_/A _26997_/Q vssd1 vssd1 vccd1 vccd1 _19227_/X
+ sky130_fd_sc_hd__a22o_1
X_16439_ _16439_/A _16439_/B _16439_/C vssd1 vssd1 vccd1 vccd1 _16439_/X sky130_fd_sc_hd__or3_1
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19158_ _18213_/X _18734_/X _19158_/S vssd1 vssd1 vccd1 vccd1 _19158_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18109_ _18292_/A vssd1 vssd1 vccd1 vccd1 _19059_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_258_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19089_ _25521_/Q _18439_/A _18441_/A _17408_/A vssd1 vssd1 vccd1 vccd1 _19089_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_160_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21120_ _21138_/A vssd1 vssd1 vccd1 vccd1 _21136_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21051_ _25894_/Q _20951_/X _21059_/S vssd1 vssd1 vccd1 vccd1 _21052_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20002_ _19993_/X _19998_/X _19999_/Y _20001_/Y vssd1 vssd1 vccd1 vccd1 _20002_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_141_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24810_ _24810_/A vssd1 vssd1 vccd1 vccd1 _24810_/X sky130_fd_sc_hd__clkbuf_1
X_25790_ _25796_/CLK _25790_/D vssd1 vssd1 vccd1 vccd1 _25790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24741_ _27092_/Q _24724_/X _24739_/Y _24740_/X vssd1 vssd1 vccd1 vccd1 _24742_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_55_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21953_ _20609_/X _26092_/Q _21955_/S vssd1 vssd1 vccd1 vccd1 _21954_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20904_ _20971_/S vssd1 vssd1 vccd1 vccd1 _20917_/S sky130_fd_sc_hd__clkbuf_4
X_24672_ _19896_/B _24657_/X _24671_/Y _24660_/X vssd1 vssd1 vccd1 vccd1 _24673_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_215_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21884_ _26293_/Q _21881_/X _21883_/X input215/X vssd1 vssd1 vccd1 vccd1 _21884_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26411_ _26796_/CLK _26411_/D vssd1 vssd1 vccd1 vccd1 _26411_/Q sky130_fd_sc_hd__dfxtp_1
X_23623_ _26720_/Q _23523_/X _23623_/S vssd1 vssd1 vccd1 vccd1 _23624_/A sky130_fd_sc_hd__mux2_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20835_ _20835_/A vssd1 vssd1 vccd1 vccd1 _25813_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26342_ _26467_/CLK _26342_/D vssd1 vssd1 vccd1 vccd1 _26342_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_23_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23554_ _23554_/A vssd1 vssd1 vccd1 vccd1 _26697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20766_ _20580_/X _25779_/Q _20772_/S vssd1 vssd1 vccd1 vccd1 _20767_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22505_ _22505_/A _22513_/B vssd1 vssd1 vccd1 vccd1 _22506_/A sky130_fd_sc_hd__and2_1
XFILLER_10_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26273_ _26292_/CLK _26273_/D vssd1 vssd1 vccd1 vccd1 _26273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23485_ _26673_/Q _23105_/X _23491_/S vssd1 vssd1 vccd1 vccd1 _23486_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20697_ _21878_/A vssd1 vssd1 vccd1 vccd1 _20697_/X sky130_fd_sc_hd__buf_6
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25224_ _27219_/Q _25204_/X _25207_/X _24729_/B _25223_/X vssd1 vssd1 vccd1 vccd1
+ _27219_/D sky130_fd_sc_hd__o221a_1
X_22436_ _26247_/Q _22444_/B vssd1 vssd1 vccd1 vccd1 _22436_/X sky130_fd_sc_hd__or2_1
XFILLER_164_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25155_ _25155_/A _25159_/B vssd1 vssd1 vccd1 vccd1 _25155_/Y sky130_fd_sc_hd__nand2_1
X_22367_ _17087_/C _26226_/Q _22376_/S vssd1 vssd1 vccd1 vccd1 _22368_/B sky130_fd_sc_hd__mux2_1
XFILLER_184_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24106_ _24106_/A vssd1 vssd1 vccd1 vccd1 _26920_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21318_ _21315_/Y _21317_/Y _21297_/X vssd1 vssd1 vccd1 vccd1 _21318_/Y sky130_fd_sc_hd__a21oi_4
X_25086_ _25113_/A vssd1 vssd1 vccd1 vccd1 _25086_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22298_ _26212_/Q _22284_/X _22297_/X _22288_/X vssd1 vssd1 vccd1 vccd1 _26212_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24037_ _26890_/Q _23555_/X _24037_/S vssd1 vssd1 vccd1 vccd1 _24038_/A sky130_fd_sc_hd__mux2_1
X_21249_ _21283_/A vssd1 vssd1 vccd1 vccd1 _21586_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15810_ _13431_/X _15807_/X _15809_/X _13863_/X vssd1 vssd1 vccd1 vccd1 _15810_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_77_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16790_ _16938_/B vssd1 vssd1 vccd1 vccd1 _16955_/B sky130_fd_sc_hd__clkbuf_2
X_25988_ _25992_/CLK _25988_/D vssd1 vssd1 vccd1 vccd1 _25988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15741_ _27278_/Q _26471_/Q _15971_/S vssd1 vssd1 vccd1 vccd1 _15741_/X sky130_fd_sc_hd__mux2_1
X_24939_ _24582_/A _24917_/X _24938_/X vssd1 vssd1 vccd1 vccd1 _24939_/Y sky130_fd_sc_hd__a21oi_1
X_12953_ _12953_/A _25481_/Q _25480_/Q vssd1 vssd1 vccd1 vccd1 _12961_/A sky130_fd_sc_hd__nor3b_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18460_ _18460_/A vssd1 vssd1 vccd1 vccd1 _18461_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_42_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27306_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15672_ _15672_/A _15672_/B vssd1 vssd1 vccd1 vccd1 _15672_/X sky130_fd_sc_hd__or2_1
XFILLER_245_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12884_ _12946_/A _13916_/C _13916_/D vssd1 vssd1 vccd1 vccd1 _13569_/B sky130_fd_sc_hd__and3_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17411_ _17430_/A _17418_/C vssd1 vssd1 vccd1 vccd1 _17411_/Y sky130_fd_sc_hd__nor2_1
XFILLER_234_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14623_ _14623_/A vssd1 vssd1 vccd1 vccd1 _17197_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26609_ _26609_/CLK _26609_/D vssd1 vssd1 vccd1 vccd1 _26609_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18391_ _18391_/A vssd1 vssd1 vccd1 vccd1 _18508_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_233_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17380_/A _17342_/B _17344_/B vssd1 vssd1 vccd1 vccd1 _25533_/D sky130_fd_sc_hd__nor3_1
XFILLER_42_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _13520_/A _26588_/Q _14375_/S _26328_/Q _14458_/S vssd1 vssd1 vccd1 vccd1
+ _14554_/X sky130_fd_sc_hd__o221a_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _13485_/X _13503_/X _13504_/X _14757_/A vssd1 vssd1 vccd1 vccd1 _13506_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17273_ _25511_/Q _25512_/Q _17273_/C vssd1 vssd1 vccd1 vccd1 _17275_/B sky130_fd_sc_hd__and3_1
X_14485_ _14485_/A _14485_/B vssd1 vssd1 vccd1 vccd1 _14485_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16224_ _16222_/X _16223_/X _16224_/S vssd1 vssd1 vccd1 vccd1 _16224_/X sky130_fd_sc_hd__mux2_1
X_19012_ _19157_/S vssd1 vssd1 vccd1 vccd1 _19328_/S sky130_fd_sc_hd__buf_2
X_13436_ _13114_/A _13415_/X _13419_/X _13168_/A _13435_/X vssd1 vssd1 vccd1 vccd1
+ _13436_/X sky130_fd_sc_hd__a311o_1
XFILLER_174_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16155_ _26801_/Q _16135_/B _15169_/A vssd1 vssd1 vccd1 vccd1 _16155_/X sky130_fd_sc_hd__o21a_1
XFILLER_127_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13367_ _13367_/A vssd1 vssd1 vccd1 vccd1 _13367_/X sky130_fd_sc_hd__buf_6
XFILLER_127_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ _16271_/S vssd1 vssd1 vccd1 vccd1 _16433_/S sky130_fd_sc_hd__buf_4
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16086_ _26671_/Q _25711_/Q _16086_/S vssd1 vssd1 vccd1 vccd1 _16086_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13298_ _15930_/S vssd1 vssd1 vccd1 vccd1 _16193_/S sky130_fd_sc_hd__buf_4
XFILLER_114_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15037_ _25895_/Q _16243_/B vssd1 vssd1 vccd1 vccd1 _15037_/X sky130_fd_sc_hd__or2_1
X_19914_ _19914_/A vssd1 vssd1 vccd1 vccd1 _19914_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19845_ _25668_/Q _19845_/B vssd1 vssd1 vccd1 vccd1 _19906_/C sky130_fd_sc_hd__and2_1
XFILLER_256_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19776_ _19776_/A _19776_/B vssd1 vssd1 vccd1 vccd1 _19777_/A sky130_fd_sc_hd__nor2_1
XFILLER_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16988_ _16996_/A vssd1 vssd1 vccd1 vccd1 _16988_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18727_ _19157_/S vssd1 vssd1 vccd1 vccd1 _19453_/S sky130_fd_sc_hd__buf_2
X_15939_ _15939_/A _15939_/B vssd1 vssd1 vccd1 vccd1 _15939_/X sky130_fd_sc_hd__or2_1
XFILLER_271_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18658_ _27015_/Q _18514_/X _18657_/X _18455_/X vssd1 vssd1 vccd1 vccd1 _18658_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17609_ _25921_/Q _17597_/X _12922_/Y _17518_/X vssd1 vssd1 vccd1 vccd1 _17609_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18589_ _25732_/Q _18588_/C _25733_/Q vssd1 vssd1 vccd1 vccd1 _18590_/B sky130_fd_sc_hd__a21oi_1
XFILLER_212_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20620_ _23609_/A vssd1 vssd1 vccd1 vccd1 _23785_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_269_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20551_ _20550_/X _25706_/Q _20551_/S vssd1 vssd1 vccd1 vccd1 _20552_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23270_ _23270_/A vssd1 vssd1 vccd1 vccd1 _26577_/D sky130_fd_sc_hd__clkbuf_1
X_20482_ _22535_/A _19755_/X _20475_/X _20481_/Y _17235_/X vssd1 vssd1 vccd1 vccd1
+ _25691_/D sky130_fd_sc_hd__a221oi_1
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22221_ _26189_/Q _22200_/X _22220_/X _22217_/X vssd1 vssd1 vccd1 vccd1 _26189_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_285_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22152_ _22152_/A vssd1 vssd1 vccd1 vccd1 _22152_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_218_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput430 _25964_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[28] sky130_fd_sc_hd__buf_2
XFILLER_161_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput441 _25945_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[9] sky130_fd_sc_hd__buf_2
Xoutput452 _25735_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[11] sky130_fd_sc_hd__buf_2
X_21103_ _25909_/Q _21094_/X _21095_/X input39/X vssd1 vssd1 vccd1 vccd1 _21104_/B
+ sky130_fd_sc_hd__o22a_1
X_26960_ _26995_/CLK _26960_/D vssd1 vssd1 vccd1 vccd1 _26960_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput463 _25745_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[21] sky130_fd_sc_hd__buf_2
X_22083_ _22083_/A vssd1 vssd1 vccd1 vccd1 _26149_/D sky130_fd_sc_hd__clkbuf_1
Xoutput474 _25755_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[31] sky130_fd_sc_hd__buf_2
XFILLER_87_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput485 _17054_/X vssd1 vssd1 vccd1 vccd1 wmask0[1] sky130_fd_sc_hd__buf_2
XFILLER_232_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21034_ _21034_/A vssd1 vssd1 vccd1 vccd1 _25886_/D sky130_fd_sc_hd__clkbuf_1
X_25911_ _27122_/CLK _25911_/D vssd1 vssd1 vccd1 vccd1 _25911_/Q sky130_fd_sc_hd__dfxtp_4
X_26891_ _27311_/CLK _26891_/D vssd1 vssd1 vccd1 vccd1 _26891_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25842_ _26468_/CLK _25842_/D vssd1 vssd1 vccd1 vccd1 _25842_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_234_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25773_ _27281_/CLK _25773_/D vssd1 vssd1 vccd1 vccd1 _25773_/Q sky130_fd_sc_hd__dfxtp_1
X_22985_ _22985_/A vssd1 vssd1 vccd1 vccd1 _26465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24724_ _24744_/A vssd1 vssd1 vccd1 vccd1 _24724_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_21936_ _20575_/X _26084_/Q _21944_/S vssd1 vssd1 vccd1 vccd1 _21937_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24655_ _27072_/Q _24636_/X _24654_/Y _24631_/X vssd1 vssd1 vccd1 vccd1 _27072_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_203_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21867_ _21885_/B vssd1 vssd1 vccd1 vccd1 _21867_/Y sky130_fd_sc_hd__inv_2
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23606_ _23606_/A vssd1 vssd1 vccd1 vccd1 _23606_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_169_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20818_ _25805_/Q vssd1 vssd1 vccd1 vccd1 _20819_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24586_ _27050_/Q _24576_/X _24585_/Y _24580_/X vssd1 vssd1 vccd1 vccd1 _27050_/D
+ sky130_fd_sc_hd__o211a_1
X_21798_ _21798_/A vssd1 vssd1 vccd1 vccd1 _26029_/D sky130_fd_sc_hd__clkbuf_1
X_26325_ _26327_/CLK _26325_/D vssd1 vssd1 vccd1 vccd1 _26325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23537_ _26692_/Q _23536_/X _23540_/S vssd1 vssd1 vccd1 vccd1 _23538_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20749_ _20749_/A vssd1 vssd1 vccd1 vccd1 _25771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26256_ _26257_/CLK _26256_/D vssd1 vssd1 vccd1 vccd1 _26256_/Q sky130_fd_sc_hd__dfxtp_1
X_14270_ _14513_/S vssd1 vssd1 vccd1 vccd1 _14332_/S sky130_fd_sc_hd__buf_2
XFILLER_10_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23468_ _23468_/A vssd1 vssd1 vccd1 vccd1 _26665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_160_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27130_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_195_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25207_ _25228_/A vssd1 vssd1 vccd1 vccd1 _25207_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13221_ _13221_/A vssd1 vssd1 vccd1 vccd1 _14791_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_109_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22419_ _22638_/A _26219_/Q _22554_/A _22419_/D vssd1 vssd1 vccd1 vccd1 _22460_/A
+ sky130_fd_sc_hd__nor4_4
X_26187_ _26222_/CLK _26187_/D vssd1 vssd1 vccd1 vccd1 _26187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23399_ _23421_/A vssd1 vssd1 vccd1 vccd1 _23408_/S sky130_fd_sc_hd__buf_4
XFILLER_128_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13152_ _26499_/Q _26371_/Q _15555_/S vssd1 vssd1 vccd1 vccd1 _13152_/X sky130_fd_sc_hd__mux2_1
X_25138_ _25138_/A vssd1 vssd1 vccd1 vccd1 _25138_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13083_ _13083_/A vssd1 vssd1 vccd1 vccd1 _13084_/A sky130_fd_sc_hd__clkbuf_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17960_ _17952_/X _17959_/X _18347_/S vssd1 vssd1 vccd1 vccd1 _17961_/B sky130_fd_sc_hd__mux2_1
X_25069_ _27178_/Q _25058_/X _25068_/X vssd1 vssd1 vccd1 vccd1 _27178_/D sky130_fd_sc_hd__o21ba_1
XFILLER_266_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16911_ _16939_/B vssd1 vssd1 vccd1 vccd1 _16911_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_238_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17891_ _14562_/B _17852_/B _17990_/A vssd1 vssd1 vccd1 vccd1 _17891_/X sky130_fd_sc_hd__mux2_1
XFILLER_266_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19630_ _19676_/A _19606_/Y _19607_/X _25218_/A vssd1 vssd1 vccd1 vccd1 _19633_/D
+ sky130_fd_sc_hd__a31o_1
X_16842_ _16842_/A vssd1 vssd1 vccd1 vccd1 _16842_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19561_ _25658_/Q _19563_/B vssd1 vssd1 vccd1 vccd1 _19561_/X sky130_fd_sc_hd__or2_1
X_13985_ _15818_/S _13982_/X _13983_/X _13984_/X _15720_/S vssd1 vssd1 vccd1 vccd1
+ _13985_/X sky130_fd_sc_hd__a221o_1
X_16773_ _16773_/A vssd1 vssd1 vccd1 vccd1 _19252_/B sky130_fd_sc_hd__buf_4
XFILLER_93_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18512_ _27108_/Q _18504_/X _18506_/X _18511_/X vssd1 vssd1 vccd1 vccd1 _18512_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_248_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12936_ input109/X input144/X _14320_/S vssd1 vssd1 vccd1 vccd1 _12937_/B sky130_fd_sc_hd__mux2_8
X_15724_ _15818_/S _15723_/X _13998_/S vssd1 vssd1 vccd1 vccd1 _15724_/X sky130_fd_sc_hd__a21o_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19492_ _19484_/X _18133_/X _19491_/X _19489_/X vssd1 vssd1 vccd1 vccd1 _25631_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18443_ _18443_/A vssd1 vssd1 vccd1 vccd1 _18444_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12867_ _12863_/X _12865_/X _12866_/X vssd1 vssd1 vccd1 vccd1 _12911_/B sky130_fd_sc_hd__a21oi_2
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ _15649_/X _15651_/X _15654_/X _15647_/S _12703_/A vssd1 vssd1 vccd1 vccd1
+ _15655_/X sky130_fd_sc_hd__o221a_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14606_ _14834_/A _14834_/B _14606_/C vssd1 vssd1 vccd1 vccd1 _15791_/C sky130_fd_sc_hd__nor3_1
XFILLER_221_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15586_ _15670_/A _15586_/B vssd1 vssd1 vccd1 vccd1 _15586_/X sky130_fd_sc_hd__or2_1
X_18374_ _18544_/A _18365_/Y _18373_/X vssd1 vssd1 vccd1 vccd1 _18374_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_15_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ _13309_/A _17504_/A vssd1 vssd1 vccd1 vccd1 _17133_/A sky130_fd_sc_hd__nor2_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _17334_/A _17331_/C vssd1 vssd1 vccd1 vccd1 _17325_/Y sky130_fd_sc_hd__nor2_1
X_14537_ _12736_/A _26876_/Q _26748_/Q _13841_/A _14384_/X vssd1 vssd1 vccd1 vccd1
+ _14537_/X sky130_fd_sc_hd__a221o_1
XFILLER_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17256_ _25507_/Q _17256_/B vssd1 vssd1 vccd1 vccd1 _17263_/C sky130_fd_sc_hd__and2_1
X_14468_ _14468_/A _14468_/B vssd1 vssd1 vccd1 vccd1 _14468_/X sky130_fd_sc_hd__or2_1
XFILLER_147_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_14_0_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_14_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_13419_ _15567_/S _13416_/X _13418_/X _13144_/A vssd1 vssd1 vccd1 vccd1 _13419_/X
+ sky130_fd_sc_hd__a211o_1
X_16207_ _16207_/A _16206_/Y vssd1 vssd1 vccd1 vccd1 _19121_/B sky130_fd_sc_hd__nor2b_4
X_17187_ _20657_/A vssd1 vssd1 vccd1 vccd1 _19352_/A sky130_fd_sc_hd__clkbuf_4
X_14399_ _13180_/A _19665_/A _14398_/X vssd1 vssd1 vccd1 vccd1 _14562_/B sky130_fd_sc_hd__o21a_1
XFILLER_255_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16138_ _26865_/Q _25779_/Q _16399_/S vssd1 vssd1 vccd1 vccd1 _16138_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16069_ _26639_/Q _26735_/Q _16069_/S vssd1 vssd1 vccd1 vccd1 _16069_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19828_ _19828_/A _20249_/B vssd1 vssd1 vccd1 vccd1 _19855_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19759_ _22478_/A _19721_/X _19746_/X _19756_/X _19758_/X vssd1 vssd1 vccd1 vccd1
+ _25664_/D sky130_fd_sc_hd__o221a_1
XFILLER_110_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22770_ _26370_/Q _22675_/X _22778_/S vssd1 vssd1 vccd1 vccd1 _22771_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21721_ _23860_/A _23139_/A vssd1 vssd1 vccd1 vccd1 _21778_/A sky130_fd_sc_hd__or2_4
XFILLER_262_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24440_ _24464_/A _24585_/A vssd1 vssd1 vccd1 vccd1 _24440_/Y sky130_fd_sc_hd__nand2_1
XFILLER_220_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21652_ _17020_/A _20978_/B _21199_/X vssd1 vssd1 vccd1 vccd1 _21652_/X sky130_fd_sc_hd__a21o_2
XFILLER_240_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20603_ _20603_/A vssd1 vssd1 vccd1 vccd1 _25718_/D sky130_fd_sc_hd__clkbuf_1
X_24371_ _24649_/B vssd1 vssd1 vccd1 vccd1 _24553_/A sky130_fd_sc_hd__inv_2
X_21583_ _21578_/Y _21582_/X _21556_/X vssd1 vssd1 vccd1 vccd1 _21583_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_178_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26110_ _26599_/CLK _26110_/D vssd1 vssd1 vccd1 vccd1 _26110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23322_ _20546_/X _26601_/Q _23324_/S vssd1 vssd1 vccd1 vccd1 _23323_/A sky130_fd_sc_hd__mux2_1
X_20534_ _20622_/S vssd1 vssd1 vccd1 vccd1 _20551_/S sky130_fd_sc_hd__buf_2
X_27090_ _27213_/CLK _27090_/D vssd1 vssd1 vccd1 vccd1 _27090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26041_ _26468_/CLK _26041_/D vssd1 vssd1 vccd1 vccd1 _26041_/Q sky130_fd_sc_hd__dfxtp_1
X_23253_ _26570_/Q _23095_/X _23255_/S vssd1 vssd1 vccd1 vccd1 _23254_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20465_ _27132_/Q vssd1 vssd1 vccd1 vccd1 _20465_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22204_ _26184_/Q _22201_/X _22115_/X _22202_/X _22203_/X vssd1 vssd1 vccd1 vccd1
+ _22204_/X sky130_fd_sc_hd__a221o_1
XFILLER_134_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23184_ _23184_/A vssd1 vssd1 vccd1 vccd1 _26539_/D sky130_fd_sc_hd__clkbuf_1
X_20396_ _20420_/B _20420_/C vssd1 vssd1 vccd1 vccd1 _20396_/X sky130_fd_sc_hd__and2_1
XFILLER_3_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22135_ _26164_/Q _22110_/X _22134_/X _22132_/X vssd1 vssd1 vccd1 vccd1 _26164_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26943_ _26980_/CLK _26943_/D vssd1 vssd1 vccd1 vccd1 _26943_/Q sky130_fd_sc_hd__dfxtp_1
X_22066_ _26142_/Q _20916_/X _22066_/S vssd1 vssd1 vccd1 vccd1 _22067_/A sky130_fd_sc_hd__mux2_1
Xoutput293 _17071_/X vssd1 vssd1 vccd1 vccd1 addr0[8] sky130_fd_sc_hd__buf_2
XFILLER_0_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_0 wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21017_ _21063_/S vssd1 vssd1 vccd1 vccd1 _21026_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_248_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26874_ _26938_/CLK _26874_/D vssd1 vssd1 vccd1 vccd1 _26874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_275_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25825_ _26715_/CLK _25825_/D vssd1 vssd1 vccd1 vccd1 _25825_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_101_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13770_ _14310_/S vssd1 vssd1 vccd1 vccd1 _15515_/S sky130_fd_sc_hd__buf_2
X_25756_ _26264_/CLK _25756_/D vssd1 vssd1 vccd1 vccd1 _25756_/Q sky130_fd_sc_hd__dfxtp_1
X_22968_ _22968_/A vssd1 vssd1 vccd1 vccd1 _26457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_261_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12721_ _12721_/A _19774_/A _16481_/A _17995_/A vssd1 vssd1 vccd1 vccd1 _12722_/C
+ sky130_fd_sc_hd__or4_1
X_21919_ _21919_/A vssd1 vssd1 vccd1 vccd1 _26076_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24707_ _24725_/A _24707_/B vssd1 vssd1 vccd1 vccd1 _24707_/Y sky130_fd_sc_hd__nand2_2
XFILLER_216_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25687_ _26286_/CLK _25687_/D vssd1 vssd1 vccd1 vccd1 _25687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22899_ _26427_/Q _22653_/X _22901_/S vssd1 vssd1 vccd1 vccd1 _22900_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15440_ _19109_/A vssd1 vssd1 vccd1 vccd1 _16612_/A sky130_fd_sc_hd__inv_2
X_24638_ _25065_/A vssd1 vssd1 vccd1 vccd1 _24639_/A sky130_fd_sc_hd__buf_2
XFILLER_71_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15371_ _26800_/Q _26444_/Q _15374_/S vssd1 vssd1 vccd1 vccd1 _15371_/X sky130_fd_sc_hd__mux2_1
X_24569_ _24569_/A _24569_/B vssd1 vssd1 vccd1 vccd1 _24569_/Y sky130_fd_sc_hd__nand2_1
XFILLER_169_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14322_ _25904_/Q _13922_/B _14321_/Y _13928_/A vssd1 vssd1 vccd1 vccd1 _14322_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_17110_ _17110_/A vssd1 vssd1 vccd1 vccd1 _25468_/D sky130_fd_sc_hd__clkbuf_1
X_26308_ _26327_/CLK _26308_/D vssd1 vssd1 vccd1 vccd1 _26308_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_157_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18090_ _20280_/B vssd1 vssd1 vccd1 vccd1 _20092_/A sky130_fd_sc_hd__buf_2
XFILLER_156_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27288_ _27288_/CLK _27288_/D vssd1 vssd1 vccd1 vccd1 _27288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17041_ _17035_/X _16943_/B _17039_/X input231/X vssd1 vssd1 vccd1 vccd1 _17041_/X
+ sky130_fd_sc_hd__a22o_4
X_26239_ _26240_/CLK _26239_/D vssd1 vssd1 vccd1 vccd1 _26239_/Q sky130_fd_sc_hd__dfxtp_1
X_14253_ _26491_/Q _26363_/Q _14253_/S vssd1 vssd1 vccd1 vccd1 _14253_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13204_ _20487_/C _13204_/B _13204_/C vssd1 vssd1 vccd1 vccd1 _13464_/A sky130_fd_sc_hd__nand3b_2
XFILLER_171_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14184_ _13107_/A _14157_/X _14166_/X _14183_/X vssd1 vssd1 vccd1 vccd1 _14184_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_99_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13135_ _13135_/A vssd1 vssd1 vccd1 vccd1 _13723_/A sky130_fd_sc_hd__buf_2
XFILLER_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18992_ _26958_/Q _18764_/X _18765_/X _26990_/Q vssd1 vssd1 vccd1 vccd1 _18992_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _15460_/S vssd1 vssd1 vccd1 vccd1 _15567_/S sky130_fd_sc_hd__clkbuf_4
X_17943_ _18210_/S vssd1 vssd1 vccd1 vccd1 _18489_/S sky130_fd_sc_hd__clkbuf_2
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17874_ _17957_/S vssd1 vssd1 vccd1 vccd1 _17954_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19613_ _27063_/Q _19616_/B _19613_/C vssd1 vssd1 vccd1 vccd1 _19614_/D sky130_fd_sc_hd__and3_1
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16825_ _16825_/A vssd1 vssd1 vccd1 vccd1 _16825_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19544_ _19538_/X _19139_/X _19543_/X _19541_/X vssd1 vssd1 vccd1 vccd1 _25651_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16756_ _16769_/A vssd1 vssd1 vccd1 vccd1 _16756_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13968_ _27269_/Q _26462_/Q _16005_/S vssd1 vssd1 vccd1 vccd1 _13968_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15707_ _15954_/A _15954_/B _15706_/X vssd1 vssd1 vccd1 vccd1 _15707_/X sky130_fd_sc_hd__or3b_1
XFILLER_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12919_ _14033_/S vssd1 vssd1 vccd1 vccd1 _14320_/S sky130_fd_sc_hd__buf_4
X_19475_ _19196_/X _19473_/Y _19474_/X _25166_/A _18777_/X vssd1 vssd1 vccd1 vccd1
+ _19475_/X sky130_fd_sc_hd__o32a_1
XFILLER_222_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13899_ _13887_/X _13895_/X _13898_/X _15983_/S _13630_/X vssd1 vssd1 vccd1 vccd1
+ _13899_/X sky130_fd_sc_hd__o221a_1
X_16687_ _16769_/A vssd1 vssd1 vccd1 vccd1 _20800_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_250_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18426_ _18858_/S _18046_/X _18271_/X vssd1 vssd1 vccd1 vccd1 _18426_/Y sky130_fd_sc_hd__o21ai_1
X_15638_ _15538_/X _15633_/X _15637_/X _14678_/A vssd1 vssd1 vccd1 vccd1 _15638_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18357_ _18357_/A _19289_/B vssd1 vssd1 vccd1 vccd1 _18357_/X sky130_fd_sc_hd__or2_1
X_15569_ _15187_/A _15560_/X _15568_/X _14708_/A vssd1 vssd1 vccd1 vccd1 _15569_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17308_ _25523_/Q vssd1 vssd1 vccd1 vccd1 _17308_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18288_ _18432_/C _18288_/B vssd1 vssd1 vccd1 vccd1 _18288_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17239_ _25109_/A vssd1 vssd1 vccd1 vccd1 _24291_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20250_ _25746_/Q vssd1 vssd1 vccd1 vccd1 _20681_/A sky130_fd_sc_hd__buf_8
XFILLER_115_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20181_ _27152_/Q _27086_/Q vssd1 vssd1 vccd1 vccd1 _20182_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_276_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23940_ _23940_/A vssd1 vssd1 vccd1 vccd1 _26846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23871_ _23699_/X _26816_/Q _23871_/S vssd1 vssd1 vccd1 vccd1 _23872_/A sky130_fd_sc_hd__mux2_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25610_ _25660_/CLK _25610_/D vssd1 vssd1 vccd1 vccd1 _25610_/Q sky130_fd_sc_hd__dfxtp_2
X_22822_ _22822_/A vssd1 vssd1 vccd1 vccd1 _26392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26590_ _26909_/CLK _26590_/D vssd1 vssd1 vccd1 vccd1 _26590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_272_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25541_ _25545_/CLK _25541_/D vssd1 vssd1 vccd1 vccd1 _25541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22753_ _22753_/A vssd1 vssd1 vccd1 vccd1 _26362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21704_ _21704_/A vssd1 vssd1 vccd1 vccd1 _25990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25472_ _25598_/CLK _25472_/D vssd1 vssd1 vccd1 vccd1 _25472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22684_ _22684_/A vssd1 vssd1 vccd1 vccd1 _26340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24423_ _24381_/X _25608_/Q _24422_/X vssd1 vssd1 vccd1 vccd1 _24686_/B sky130_fd_sc_hd__o21a_4
X_27211_ _27228_/CLK _27211_/D vssd1 vssd1 vccd1 vccd1 _27211_/Q sky130_fd_sc_hd__dfxtp_1
X_21635_ input66/X input101/X _21646_/S vssd1 vssd1 vccd1 vccd1 _21636_/A sky130_fd_sc_hd__mux2_8
XFILLER_21_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27142_ _27166_/CLK _27142_/D vssd1 vssd1 vccd1 vccd1 _27142_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_139_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24354_ _25206_/C _24633_/C vssd1 vssd1 vccd1 vccd1 _24776_/C sky130_fd_sc_hd__nor2_1
X_21566_ _25865_/Q vssd1 vssd1 vccd1 vccd1 _21566_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_193_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23305_ _20512_/X _26593_/Q _23313_/S vssd1 vssd1 vccd1 vccd1 _23306_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20517_ _23706_/A vssd1 vssd1 vccd1 vccd1 _20517_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_27073_ _27203_/CLK _27073_/D vssd1 vssd1 vccd1 vccd1 _27073_/Q sky130_fd_sc_hd__dfxtp_1
X_24285_ _24285_/A _24285_/B _24286_/B vssd1 vssd1 vccd1 vccd1 _26985_/D sky130_fd_sc_hd__nor3_1
XFILLER_153_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21497_ _21495_/X _21496_/X _21433_/X vssd1 vssd1 vccd1 vccd1 _21497_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26024_ _26903_/CLK _26024_/D vssd1 vssd1 vccd1 vccd1 _26024_/Q sky130_fd_sc_hd__dfxtp_1
X_23236_ _26562_/Q _23069_/X _23244_/S vssd1 vssd1 vccd1 vccd1 _23237_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20448_ _20448_/A _20448_/B vssd1 vssd1 vccd1 vccd1 _20449_/B sky130_fd_sc_hd__or2_1
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23167_ _23167_/A vssd1 vssd1 vccd1 vccd1 _26531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20379_ _20379_/A _20379_/B vssd1 vssd1 vccd1 vccd1 _20398_/B sky130_fd_sc_hd__xnor2_1
XFILLER_122_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22118_ _22155_/A vssd1 vssd1 vccd1 vccd1 _22118_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_267_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23098_ _23571_/A vssd1 vssd1 vccd1 vccd1 _23098_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22049_ _26134_/Q _20891_/X _22055_/S vssd1 vssd1 vccd1 vccd1 _22050_/A sky130_fd_sc_hd__mux2_1
X_14940_ _25626_/Q _14597_/X _14939_/X _14618_/X vssd1 vssd1 vccd1 vccd1 _23600_/A
+ sky130_fd_sc_hd__o22a_4
X_26926_ _27308_/CLK _26926_/D vssd1 vssd1 vccd1 vccd1 _26926_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_134_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26857_ _27308_/CLK _26857_/D vssd1 vssd1 vccd1 vccd1 _26857_/Q sky130_fd_sc_hd__dfxtp_2
X_14871_ _16320_/S vssd1 vssd1 vccd1 vccd1 _16224_/S sky130_fd_sc_hd__buf_4
XTAP_5799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16610_ _19105_/S _16613_/A vssd1 vssd1 vccd1 vccd1 _19121_/A sky130_fd_sc_hd__nand2_4
X_13822_ _15769_/A _13819_/X _13821_/X _13762_/A vssd1 vssd1 vccd1 vccd1 _13822_/X
+ sky130_fd_sc_hd__o211a_1
X_25808_ _26917_/CLK _25808_/D vssd1 vssd1 vccd1 vccd1 _25808_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_235_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17590_ _19455_/C _17584_/X _17572_/X _17589_/X vssd1 vssd1 vccd1 vccd1 _17591_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_26788_ _26916_/CLK _26788_/D vssd1 vssd1 vccd1 vccd1 _26788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_107 _21618_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_118 _23032_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13753_ _13011_/A _23536_/A _13028_/A vssd1 vssd1 vccd1 vccd1 _13753_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16541_ _26519_/Q _26391_/Q _16541_/S vssd1 vssd1 vccd1 vccd1 _16541_/X sky130_fd_sc_hd__mux2_1
XFILLER_244_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25739_ _26282_/CLK _25739_/D vssd1 vssd1 vccd1 vccd1 _25739_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_129 _14362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12704_ _12704_/A vssd1 vssd1 vccd1 vccd1 _12705_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19260_ _27126_/Q _18504_/X _19258_/X _19259_/X vssd1 vssd1 vccd1 vccd1 _19260_/X
+ sky130_fd_sc_hd__o22a_2
X_13684_ _13638_/X _23539_/A _13682_/X _13683_/X vssd1 vssd1 vccd1 vccd1 _19882_/A
+ sky130_fd_sc_hd__o211a_4
X_16472_ _12760_/B _16469_/X _16471_/X vssd1 vssd1 vccd1 vccd1 _16472_/X sky130_fd_sc_hd__o21a_1
XFILLER_31_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18211_ _18207_/X _18210_/X _18684_/S vssd1 vssd1 vccd1 vccd1 _18211_/X sky130_fd_sc_hd__mux2_1
XPHY_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15423_ _25817_/Q _27251_/Q _15662_/S vssd1 vssd1 vccd1 vccd1 _15424_/B sky130_fd_sc_hd__mux2_1
X_19191_ _19392_/A _19191_/B vssd1 vssd1 vccd1 vccd1 _19191_/Y sky130_fd_sc_hd__nor2_1
XPHY_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18142_ _18895_/A _18087_/X _19078_/A _18141_/X vssd1 vssd1 vccd1 vccd1 _18142_/X
+ sky130_fd_sc_hd__a22o_1
X_15354_ _26864_/Q _25778_/Q _16395_/S vssd1 vssd1 vccd1 vccd1 _15354_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14305_ _13239_/A _14303_/X _14304_/X _13278_/A vssd1 vssd1 vccd1 vccd1 _14305_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18073_ _18729_/A _18073_/B vssd1 vssd1 vccd1 vccd1 _18073_/X sky130_fd_sc_hd__or2_1
X_15285_ _15285_/A _15285_/B vssd1 vssd1 vccd1 vccd1 _15285_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17024_ _17021_/X _16870_/B _17017_/X input218/X vssd1 vssd1 vccd1 vccd1 _17024_/X
+ sky130_fd_sc_hd__a22o_4
X_14236_ _18001_/A _17776_/A vssd1 vssd1 vccd1 vccd1 _14362_/B sky130_fd_sc_hd__or2_2
XFILLER_153_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14167_ _14354_/S vssd1 vssd1 vccd1 vccd1 _14440_/S sky130_fd_sc_hd__buf_2
XFILLER_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13118_ _15460_/S vssd1 vssd1 vccd1 vccd1 _15174_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_152_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14098_ _13889_/A _14096_/X _14097_/X vssd1 vssd1 vccd1 vccd1 _14098_/Y sky130_fd_sc_hd__o21ai_1
X_18975_ _18975_/A _18978_/A vssd1 vssd1 vccd1 vccd1 _18975_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_252_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13049_ _13049_/A vssd1 vssd1 vccd1 vccd1 _13050_/A sky130_fd_sc_hd__clkbuf_2
X_17926_ _17922_/X _17924_/X _18042_/S vssd1 vssd1 vccd1 vccd1 _17926_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17857_ _17857_/A vssd1 vssd1 vccd1 vccd1 _17857_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16808_ _16951_/A vssd1 vssd1 vccd1 vccd1 _16824_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_226_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17788_ _17846_/A _17785_/X _17787_/Y vssd1 vssd1 vccd1 vccd1 _17789_/B sky130_fd_sc_hd__o21a_1
XFILLER_82_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19527_ _25645_/Q _19536_/B vssd1 vssd1 vccd1 vccd1 _19527_/X sky130_fd_sc_hd__or2_1
XFILLER_207_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16739_ _25672_/Q vssd1 vssd1 vccd1 vccd1 _22496_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19458_ _19456_/X _19457_/X _19452_/A _16788_/A vssd1 vssd1 vccd1 vccd1 _19458_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_50_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18409_ _19253_/A vssd1 vssd1 vccd1 vccd1 _18409_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19389_ _19392_/B _19389_/B _19389_/C vssd1 vssd1 vccd1 vccd1 _19389_/X sky130_fd_sc_hd__and3_1
XFILLER_148_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21420_ _21414_/X _21419_/X _21407_/X vssd1 vssd1 vccd1 vccd1 _21420_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_277_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21351_ _20643_/A _21343_/X _21348_/X _21350_/X vssd1 vssd1 vccd1 vccd1 _21351_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20302_ _20302_/A vssd1 vssd1 vccd1 vccd1 _20302_/Y sky130_fd_sc_hd__inv_2
X_24070_ _26905_/Q _23603_/X _24070_/S vssd1 vssd1 vccd1 vccd1 _24071_/A sky130_fd_sc_hd__mux2_1
X_21282_ _25471_/Q _21332_/B vssd1 vssd1 vccd1 vccd1 _21282_/X sky130_fd_sc_hd__or2_1
XFILLER_190_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23021_ _23021_/A vssd1 vssd1 vccd1 vccd1 _26481_/D sky130_fd_sc_hd__clkbuf_1
X_20233_ _25681_/Q _25680_/Q _20233_/C vssd1 vssd1 vccd1 vccd1 _20286_/C sky130_fd_sc_hd__and3_1
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20164_ _25679_/Q _20164_/B vssd1 vssd1 vccd1 vccd1 _20233_/C sky130_fd_sc_hd__and2_1
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24972_ _24972_/A _24972_/B vssd1 vssd1 vccd1 vccd1 _24972_/Y sky130_fd_sc_hd__nand2_1
X_20095_ _20095_/A _20095_/B vssd1 vssd1 vccd1 vccd1 _20204_/A sky130_fd_sc_hd__xnor2_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26711_ _26903_/CLK _26711_/D vssd1 vssd1 vccd1 vccd1 _26711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23923_ _23923_/A vssd1 vssd1 vccd1 vccd1 _26839_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26642_ _27317_/CLK _26642_/D vssd1 vssd1 vccd1 vccd1 _26642_/Q sky130_fd_sc_hd__dfxtp_1
X_23854_ _23779_/X _26809_/Q _23854_/S vssd1 vssd1 vccd1 vccd1 _23855_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22805_ _26386_/Q _22727_/X _22811_/S vssd1 vssd1 vccd1 vccd1 _22806_/A sky130_fd_sc_hd__mux2_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23785_ _23785_/A vssd1 vssd1 vccd1 vccd1 _23785_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26573_ _27315_/CLK _26573_/D vssd1 vssd1 vccd1 vccd1 _26573_/Q sky130_fd_sc_hd__dfxtp_1
X_20997_ _20997_/A vssd1 vssd1 vccd1 vccd1 _25869_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25524_ _25985_/CLK _25524_/D vssd1 vssd1 vccd1 vccd1 _25524_/Q sky130_fd_sc_hd__dfxtp_1
X_22736_ _23779_/A vssd1 vssd1 vccd1 vccd1 _22736_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25455_ _23773_/X _27322_/Q _25459_/S vssd1 vssd1 vccd1 vccd1 _25456_/A sky130_fd_sc_hd__mux2_1
X_22667_ _26335_/Q _22666_/X _22673_/S vssd1 vssd1 vccd1 vccd1 _22668_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24406_ _24361_/S _25605_/Q _24405_/X vssd1 vssd1 vccd1 vccd1 _24671_/B sky130_fd_sc_hd__o21a_4
X_21618_ _21614_/Y _21617_/X _21202_/A vssd1 vssd1 vccd1 vccd1 _21618_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_166_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25386_ _25386_/A vssd1 vssd1 vccd1 vccd1 _27291_/D sky130_fd_sc_hd__clkbuf_1
X_22598_ _22593_/X _22597_/Y _22587_/X vssd1 vssd1 vccd1 vccd1 _26314_/D sky130_fd_sc_hd__a21oi_1
XFILLER_139_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24337_ _27004_/Q _24335_/B _24314_/X vssd1 vssd1 vccd1 vccd1 _24337_/Y sky130_fd_sc_hd__a21oi_1
X_27125_ _27130_/CLK _27125_/D vssd1 vssd1 vccd1 vccd1 _27125_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_67_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26594_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_193_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21549_ _21546_/X _21548_/X _21512_/X vssd1 vssd1 vccd1 vccd1 _21549_/X sky130_fd_sc_hd__a21o_1
XFILLER_126_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27056_ _27062_/CLK _27056_/D vssd1 vssd1 vccd1 vccd1 _27056_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15070_ _12705_/A _15056_/X _15069_/X _14710_/A vssd1 vssd1 vccd1 vccd1 _15070_/X
+ sky130_fd_sc_hd__a211o_1
X_24268_ _26980_/Q _24268_/B vssd1 vssd1 vccd1 vccd1 _24275_/C sky130_fd_sc_hd__and2_1
XFILLER_181_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26007_ _27277_/CLK _26007_/D vssd1 vssd1 vccd1 vccd1 _26007_/Q sky130_fd_sc_hd__dfxtp_2
X_14021_ _14022_/A _17798_/A vssd1 vssd1 vccd1 vccd1 _18428_/S sky130_fd_sc_hd__and2_1
X_23219_ _23219_/A vssd1 vssd1 vccd1 vccd1 _26554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24199_ _26956_/Q _24195_/B _24198_/Y vssd1 vssd1 vccd1 vccd1 _26956_/D sky130_fd_sc_hd__o21a_1
XFILLER_162_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18760_ _27017_/Q _18756_/X _18758_/X _18759_/X vssd1 vssd1 vccd1 vccd1 _18760_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_283_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15972_ _25881_/Q _15972_/B vssd1 vssd1 vccd1 vccd1 _15972_/X sky130_fd_sc_hd__or2_1
XFILLER_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17711_ _17736_/B _17736_/C _17711_/C vssd1 vssd1 vccd1 vccd1 _17725_/D sky130_fd_sc_hd__and3_1
XFILLER_276_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26909_ _26909_/CLK _26909_/D vssd1 vssd1 vccd1 vccd1 _26909_/Q sky130_fd_sc_hd__dfxtp_1
X_14923_ _14921_/X _14922_/X _15004_/S vssd1 vssd1 vccd1 vccd1 _14923_/X sky130_fd_sc_hd__mux2_1
XTAP_5574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18691_ _25512_/Q _18439_/X _18441_/X _17375_/X vssd1 vssd1 vccd1 vccd1 _18691_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17642_ _17592_/A _17627_/X _14139_/X _17597_/X _25930_/Q vssd1 vssd1 vccd1 vccd1
+ _17642_/Y sky130_fd_sc_hd__o32ai_2
XFILLER_36_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14854_ _26357_/Q _26617_/Q _14876_/S vssd1 vssd1 vccd1 vccd1 _14854_/X sky130_fd_sc_hd__mux2_1
XFILLER_264_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13805_ _13966_/A vssd1 vssd1 vccd1 vccd1 _15999_/A sky130_fd_sc_hd__clkbuf_2
X_17573_ _25912_/Q _17568_/X _13395_/Y _17525_/X vssd1 vssd1 vccd1 vccd1 _17573_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_263_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14785_ _16517_/A _14783_/X _14784_/X _14760_/X vssd1 vssd1 vccd1 vccd1 _14785_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19312_ _19234_/A _19310_/Y _19311_/X _19318_/B _18839_/X vssd1 vssd1 vccd1 vccd1
+ _19312_/X sky130_fd_sc_hd__o32a_1
XFILLER_205_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16524_ _16524_/A vssd1 vssd1 vccd1 vccd1 _16540_/S sky130_fd_sc_hd__buf_2
X_13736_ input123/X input158/X _14132_/S vssd1 vssd1 vccd1 vccd1 _13736_/X sky130_fd_sc_hd__mux2_8
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19243_ _19235_/Y _19239_/X _19242_/X _18738_/X vssd1 vssd1 vccd1 vccd1 _19243_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16455_ _17846_/D vssd1 vssd1 vccd1 vccd1 _19327_/A sky130_fd_sc_hd__buf_2
X_13667_ _13779_/A _13663_/X _13666_/X _13479_/A vssd1 vssd1 vccd1 vccd1 _13671_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_220_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ _15406_/A vssd1 vssd1 vccd1 vccd1 _15406_/X sky130_fd_sc_hd__buf_2
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19174_ _18741_/X _19172_/X _19173_/Y vssd1 vssd1 vccd1 vccd1 _19174_/Y sky130_fd_sc_hd__a21oi_1
X_13598_ _13596_/X _13597_/X _15727_/S vssd1 vssd1 vccd1 vccd1 _13598_/X sky130_fd_sc_hd__mux2_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16386_ _16384_/X _16385_/X _16386_/S vssd1 vssd1 vccd1 vccd1 _16386_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18125_ _18460_/A vssd1 vssd1 vccd1 vccd1 _18569_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_200_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15337_ _15310_/X _15336_/X _14723_/A vssd1 vssd1 vccd1 vccd1 _15337_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_184_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18056_ _18046_/X _18054_/X _18684_/S vssd1 vssd1 vccd1 vccd1 _18056_/X sky130_fd_sc_hd__mux2_2
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15268_ _15142_/X _15264_/X _15267_/X _14660_/A vssd1 vssd1 vccd1 vccd1 _15268_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17007_ _16784_/X _17001_/X _16818_/C _17006_/X input237/X vssd1 vssd1 vccd1 vccd1
+ _17007_/X sky130_fd_sc_hd__a32o_4
X_14219_ _13475_/A _14217_/X _14218_/X _13775_/A vssd1 vssd1 vccd1 vccd1 _14219_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15199_ _16255_/S vssd1 vssd1 vccd1 vccd1 _15228_/S sky130_fd_sc_hd__buf_2
XFILLER_153_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18958_ _18555_/A _18948_/X _18957_/X vssd1 vssd1 vccd1 vccd1 _18958_/X sky130_fd_sc_hd__a21o_4
XFILLER_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17909_ _17824_/B _15438_/B _17909_/S vssd1 vssd1 vccd1 vccd1 _17909_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18889_ _25612_/Q _18719_/X _18888_/X _18790_/X vssd1 vssd1 vccd1 vccd1 _25612_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_282_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20920_ _20952_/A vssd1 vssd1 vccd1 vccd1 _20933_/S sky130_fd_sc_hd__buf_4
XFILLER_254_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20851_ _20851_/A vssd1 vssd1 vccd1 vccd1 _25821_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_254_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23570_ _23570_/A vssd1 vssd1 vccd1 vccd1 _26702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20782_ _20782_/A vssd1 vssd1 vccd1 vccd1 _25786_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_460 _18663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_471 _22031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22521_ _22521_/A vssd1 vssd1 vccd1 vccd1 _26284_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_482 _17545_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_493 _17697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25240_ _27226_/Q _25217_/X _25239_/X _25221_/X vssd1 vssd1 vccd1 vccd1 _27226_/D
+ sky130_fd_sc_hd__o211a_1
X_22452_ _26253_/Q _22457_/B vssd1 vssd1 vccd1 vccd1 _22452_/X sky130_fd_sc_hd__or2_1
XFILLER_167_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21403_ _21547_/A vssd1 vssd1 vccd1 vccd1 _21403_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25171_ _25206_/B _25206_/C _25206_/D vssd1 vssd1 vccd1 vccd1 _25198_/A sky130_fd_sc_hd__or3_2
X_22383_ _22350_/S _22406_/B _22236_/C vssd1 vssd1 vccd1 vccd1 _22383_/X sky130_fd_sc_hd__o21ba_1
XFILLER_163_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24122_ _24133_/A vssd1 vssd1 vccd1 vccd1 _24131_/S sky130_fd_sc_hd__buf_4
XFILLER_194_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21334_ _21332_/X _21333_/X _21290_/X vssd1 vssd1 vccd1 vccd1 _21334_/X sky130_fd_sc_hd__a21o_1
XFILLER_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24053_ _26897_/Q _23578_/X _24059_/S vssd1 vssd1 vccd1 vccd1 _24054_/A sky130_fd_sc_hd__mux2_1
X_21265_ _25470_/Q _21507_/A vssd1 vssd1 vccd1 vccd1 _21265_/X sky130_fd_sc_hd__or2_1
XFILLER_237_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23004_ _26474_/Q _22701_/X _23006_/S vssd1 vssd1 vccd1 vccd1 _23005_/A sky130_fd_sc_hd__mux2_1
XFILLER_277_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20216_ _20180_/Y _20184_/B _20182_/B vssd1 vssd1 vccd1 vccd1 _20218_/C sky130_fd_sc_hd__o21a_1
XFILLER_116_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21196_ input9/X _21075_/B _21192_/X _21195_/Y vssd1 vssd1 vccd1 vccd1 _21197_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_249_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20147_ _20200_/A _20148_/B vssd1 vssd1 vccd1 vccd1 _20174_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24955_ hold2/X _24972_/B vssd1 vssd1 vccd1 vccd1 _24955_/Y sky130_fd_sc_hd__nand2_1
X_20078_ _20225_/A vssd1 vssd1 vccd1 vccd1 _20078_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_114_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27001_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23906_ _23917_/A vssd1 vssd1 vccd1 vccd1 _23915_/S sky130_fd_sc_hd__buf_4
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24886_ _24884_/Y _24885_/X _24871_/X vssd1 vssd1 vccd1 vccd1 _27128_/D sky130_fd_sc_hd__a21oi_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26625_ _26657_/CLK _26625_/D vssd1 vssd1 vccd1 vccd1 _26625_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23837_ _23754_/X _26801_/Q _23843_/S vssd1 vssd1 vccd1 vccd1 _23838_/A sky130_fd_sc_hd__mux2_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14570_ _17966_/A _14570_/B vssd1 vssd1 vccd1 vccd1 _14570_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26556_ _26657_/CLK _26556_/D vssd1 vssd1 vccd1 vccd1 _26556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23768_ _23766_/X _26773_/Q _23780_/S vssd1 vssd1 vccd1 vccd1 _23769_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13521_ _13521_/A vssd1 vssd1 vccd1 vccd1 _15490_/A sky130_fd_sc_hd__clkbuf_4
X_25507_ _27014_/CLK _25507_/D vssd1 vssd1 vccd1 vccd1 _25507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22719_ _22719_/A vssd1 vssd1 vccd1 vccd1 _26351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23699_ _23699_/A vssd1 vssd1 vccd1 vccd1 _23699_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26487_ _26913_/CLK _26487_/D vssd1 vssd1 vccd1 vccd1 _26487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13452_ _13711_/A _13447_/X _13451_/Y _13031_/A vssd1 vssd1 vccd1 vccd1 _13452_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_202_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16240_ _26511_/Q _26383_/Q _16240_/S vssd1 vssd1 vccd1 vccd1 _16240_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25438_ _25438_/A vssd1 vssd1 vccd1 vccd1 _27314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13383_ _17817_/D vssd1 vssd1 vccd1 vccd1 _18686_/A sky130_fd_sc_hd__buf_2
X_25369_ _25369_/A vssd1 vssd1 vccd1 vccd1 _27283_/D sky130_fd_sc_hd__clkbuf_1
X_16171_ _12751_/A _16368_/S _15244_/X _16170_/Y vssd1 vssd1 vccd1 vccd1 _17791_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_167_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15122_ _14744_/A _26902_/Q _26774_/Q _16422_/S _14771_/A vssd1 vssd1 vccd1 vccd1
+ _15122_/X sky130_fd_sc_hd__a221o_1
X_27108_ _27110_/CLK _27108_/D vssd1 vssd1 vccd1 vccd1 _27108_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_154_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15053_ _26546_/Q _26154_/Q _16380_/B vssd1 vssd1 vccd1 vccd1 _15053_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19930_ _19930_/A _27077_/Q vssd1 vssd1 vccd1 vccd1 _19933_/B sky130_fd_sc_hd__nand2_1
X_27039_ _27044_/CLK _27039_/D vssd1 vssd1 vccd1 vccd1 _27039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_269_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14004_ _26850_/Q _25764_/Q _14004_/S vssd1 vssd1 vccd1 vccd1 _14004_/X sky130_fd_sc_hd__mux2_1
X_19861_ _19766_/X _19860_/X _20208_/A vssd1 vssd1 vccd1 vccd1 _19861_/X sky130_fd_sc_hd__a21o_1
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18812_ _18812_/A vssd1 vssd1 vccd1 vccd1 _18812_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_284_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19792_ _22480_/A _19721_/X _19783_/X _19791_/X _19758_/X vssd1 vssd1 vccd1 vccd1
+ _25665_/D sky130_fd_sc_hd__o221a_1
XFILLER_95_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18743_ _18807_/A vssd1 vssd1 vccd1 vccd1 _18743_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15955_ _12871_/Y _15953_/X _15954_/X _12943_/Y _14138_/Y vssd1 vssd1 vccd1 vccd1
+ _15955_/X sky130_fd_sc_hd__a32o_1
XTAP_5371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput160 dout1[58] vssd1 vssd1 vccd1 vccd1 input160/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput171 irq[0] vssd1 vssd1 vccd1 vccd1 input171/X sky130_fd_sc_hd__buf_6
XFILLER_76_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput182 irq[5] vssd1 vssd1 vccd1 vccd1 _19617_/C sky130_fd_sc_hd__buf_4
XFILLER_36_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14906_ _14746_/A _26905_/Q _26777_/Q _14981_/S _14772_/A vssd1 vssd1 vccd1 vccd1
+ _14906_/X sky130_fd_sc_hd__a221o_1
Xinput193 localMemory_wb_adr_i[12] vssd1 vssd1 vccd1 vccd1 input193/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18674_ _18340_/A _18785_/A _18678_/A vssd1 vssd1 vccd1 vccd1 _18712_/A sky130_fd_sc_hd__o21a_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15886_ _26793_/Q _26437_/Q _15888_/S vssd1 vssd1 vccd1 vccd1 _15887_/B sky130_fd_sc_hd__mux2_1
XFILLER_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ _17738_/B _17584_/X _17604_/X _17624_/Y vssd1 vssd1 vccd1 vccd1 _17626_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14837_ _14601_/X _14835_/Y _14836_/X vssd1 vssd1 vccd1 vccd1 _14837_/X sky130_fd_sc_hd__o21a_1
XFILLER_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17556_ _17592_/A _17556_/B _17556_/C vssd1 vssd1 vccd1 vccd1 _17556_/X sky130_fd_sc_hd__or3_1
X_14768_ _14768_/A vssd1 vssd1 vccd1 vccd1 _15210_/A sky130_fd_sc_hd__clkbuf_4
X_16507_ _16463_/X _23609_/A _16506_/X _15388_/X vssd1 vssd1 vccd1 vccd1 _16982_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_189_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13719_ _13719_/A vssd1 vssd1 vccd1 vccd1 _15634_/S sky130_fd_sc_hd__buf_4
XFILLER_60_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17487_ _26255_/Q _17455_/A _17461_/A _25983_/Q vssd1 vssd1 vccd1 vccd1 _17683_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_108_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14699_ _26810_/Q _26454_/Q _14699_/S vssd1 vssd1 vccd1 vccd1 _14699_/X sky130_fd_sc_hd__mux2_1
XFILLER_258_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19226_ _27061_/Q _18503_/A _19223_/X _19225_/X _18519_/A vssd1 vssd1 vccd1 vccd1
+ _19226_/X sky130_fd_sc_hd__o221a_2
XFILLER_177_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16438_ _16336_/X _16436_/X _16437_/X _14758_/A vssd1 vssd1 vccd1 vccd1 _16439_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19157_ _19579_/D _19183_/B _19157_/S vssd1 vssd1 vccd1 vccd1 _19157_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16369_ _17784_/A _17783_/A vssd1 vssd1 vccd1 vccd1 _16370_/A sky130_fd_sc_hd__nand2_1
XFILLER_118_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18108_ _17753_/A _18108_/B vssd1 vssd1 vccd1 vccd1 _18292_/A sky130_fd_sc_hd__and2b_1
XFILLER_258_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19088_ _19219_/A _19118_/B vssd1 vssd1 vccd1 vccd1 _19088_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18039_ _19571_/A _18042_/S _17807_/Y _18038_/Y vssd1 vssd1 vccd1 vccd1 _18039_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_132_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21050_ _21050_/A vssd1 vssd1 vccd1 vccd1 _21059_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_98_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_259_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_259_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20001_ _27145_/Q _20219_/B vssd1 vssd1 vccd1 vccd1 _20001_/Y sky130_fd_sc_hd__nand2_1
XFILLER_275_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21952_ _21952_/A vssd1 vssd1 vccd1 vccd1 _26091_/D sky130_fd_sc_hd__clkbuf_1
X_24740_ _24740_/A vssd1 vssd1 vccd1 vccd1 _24740_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_223_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20903_ _23718_/A vssd1 vssd1 vccd1 vccd1 _20903_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24671_ _24765_/A _24671_/B vssd1 vssd1 vccd1 vccd1 _24671_/Y sky130_fd_sc_hd__nand2_4
X_21883_ _24474_/A vssd1 vssd1 vccd1 vccd1 _21883_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_270_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26410_ _27281_/CLK _26410_/D vssd1 vssd1 vccd1 vccd1 _26410_/Q sky130_fd_sc_hd__dfxtp_1
X_23622_ _23622_/A vssd1 vssd1 vccd1 vccd1 _26719_/D sky130_fd_sc_hd__clkbuf_1
X_20834_ _25813_/Q vssd1 vssd1 vccd1 vccd1 _20835_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26341_ _26601_/CLK _26341_/D vssd1 vssd1 vccd1 vccd1 _26341_/Q sky130_fd_sc_hd__dfxtp_2
X_23553_ _26697_/Q _23552_/X _23556_/S vssd1 vssd1 vccd1 vccd1 _23554_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20765_ _20765_/A vssd1 vssd1 vccd1 vccd1 _25778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_290 _25820_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22504_ _22515_/A vssd1 vssd1 vccd1 vccd1 _22513_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26272_ _26292_/CLK _26272_/D vssd1 vssd1 vccd1 vccd1 _26272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23484_ _23484_/A vssd1 vssd1 vccd1 vccd1 _26672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20696_ _20696_/A _20703_/B vssd1 vssd1 vccd1 vccd1 _20696_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25223_ _19614_/A _25209_/X _25179_/A vssd1 vssd1 vccd1 vccd1 _25223_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22435_ _26198_/Q _22432_/X _22434_/X _22428_/X vssd1 vssd1 vccd1 vccd1 _26246_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25154_ _19381_/A _25138_/X _25153_/X vssd1 vssd1 vccd1 vccd1 _25154_/X sky130_fd_sc_hd__o21a_1
X_22366_ _22366_/A vssd1 vssd1 vccd1 vccd1 _26232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24105_ _26920_/Q _23549_/X _24109_/S vssd1 vssd1 vccd1 vccd1 _24106_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21317_ _21231_/X _21316_/X _21259_/A vssd1 vssd1 vccd1 vccd1 _21317_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_2_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25085_ _25137_/A vssd1 vssd1 vccd1 vccd1 _25085_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22297_ _26211_/Q _22294_/X _22285_/X _26312_/Q _22286_/X vssd1 vssd1 vccd1 vccd1
+ _22297_/X sky130_fd_sc_hd__a221o_1
XFILLER_117_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24036_ _24036_/A vssd1 vssd1 vccd1 vccd1 _26889_/D sky130_fd_sc_hd__clkbuf_1
X_21248_ _25469_/Q _21507_/A vssd1 vssd1 vccd1 vccd1 _21248_/X sky130_fd_sc_hd__or2_1
XFILLER_116_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21179_ _21188_/A _21179_/B vssd1 vssd1 vccd1 vccd1 _21180_/A sky130_fd_sc_hd__or2_1
XFILLER_120_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25987_ _25992_/CLK _25987_/D vssd1 vssd1 vccd1 vccd1 _25987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15740_ _15738_/X _15739_/X _15979_/S vssd1 vssd1 vccd1 vccd1 _15740_/X sky130_fd_sc_hd__mux2_1
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12952_ _12871_/Y _12931_/X _14239_/A _12943_/Y _12951_/X vssd1 vssd1 vccd1 vccd1
+ _12952_/Y sky130_fd_sc_hd__a221oi_2
X_24938_ _24938_/A vssd1 vssd1 vccd1 vccd1 _24938_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _26504_/Q _26376_/Q _15671_/S vssd1 vssd1 vccd1 vccd1 _15672_/B sky130_fd_sc_hd__mux2_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _25482_/Q _12962_/C _12947_/B vssd1 vssd1 vccd1 vccd1 _13916_/D sky130_fd_sc_hd__a21oi_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24869_ _27124_/Q _24873_/B vssd1 vssd1 vccd1 vccd1 _24869_/Y sky130_fd_sc_hd__nand2_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _25555_/Q _17410_/B vssd1 vssd1 vccd1 vccd1 _17418_/C sky130_fd_sc_hd__and2_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _14622_/A vssd1 vssd1 vccd1 vccd1 _14623_/A sky130_fd_sc_hd__clkbuf_4
X_26608_ _27283_/CLK _26608_/D vssd1 vssd1 vccd1 vccd1 _26608_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _27204_/Q _18949_/B vssd1 vssd1 vccd1 vccd1 _18390_/X sky130_fd_sc_hd__and2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _25533_/Q _25532_/Q _17341_/C vssd1 vssd1 vccd1 vccd1 _17344_/B sky130_fd_sc_hd__and3_1
XFILLER_42_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14553_ _26488_/Q _26360_/Q _14553_/S vssd1 vssd1 vccd1 vccd1 _14553_/X sky130_fd_sc_hd__mux2_1
X_26539_ _26673_/CLK _26539_/D vssd1 vssd1 vccd1 vccd1 _26539_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_82_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26751_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_187_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _15109_/A _26106_/Q _26007_/Q _13492_/X _13494_/X vssd1 vssd1 vccd1 vccd1
+ _13504_/X sky130_fd_sc_hd__a221o_1
XFILLER_198_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17272_ _17268_/X _17273_/C _25512_/Q vssd1 vssd1 vccd1 vccd1 _17274_/B sky130_fd_sc_hd__a21oi_1
X_14484_ _25630_/Q _13933_/A _14401_/B _13557_/A vssd1 vssd1 vccd1 vccd1 _14484_/X
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_11_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27284_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_174_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19011_ _19011_/A _19011_/B vssd1 vssd1 vccd1 vccd1 _19575_/B sky130_fd_sc_hd__xnor2_2
X_16223_ _25852_/Q _26052_/Q _16223_/S vssd1 vssd1 vccd1 vccd1 _16223_/X sky130_fd_sc_hd__mux2_1
X_13435_ _13144_/A _13426_/X _13434_/X _13164_/A vssd1 vssd1 vccd1 vccd1 _13435_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_228_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13366_ _13366_/A vssd1 vssd1 vccd1 vccd1 _13367_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16154_ _26445_/Q _16154_/B vssd1 vssd1 vccd1 vccd1 _16154_/X sky130_fd_sc_hd__or2_1
XFILLER_177_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15105_ _16182_/S vssd1 vssd1 vccd1 vccd1 _16271_/S sky130_fd_sc_hd__buf_4
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13297_ _15768_/S vssd1 vssd1 vccd1 vccd1 _15930_/S sky130_fd_sc_hd__clkbuf_4
X_16085_ _12756_/A _16204_/S _15244_/X _16084_/Y vssd1 vssd1 vccd1 vccd1 _16124_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_6_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15036_ _27289_/Q _26482_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _15036_/X sky130_fd_sc_hd__mux2_1
X_19913_ _20194_/B _18651_/Y _19911_/X _19912_/Y vssd1 vssd1 vccd1 vccd1 _19913_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_174_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19844_ _22485_/A _19721_/X _19838_/X _19843_/X _19758_/X vssd1 vssd1 vccd1 vccd1
+ _25667_/D sky130_fd_sc_hd__o221a_1
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19775_ _19805_/A _19805_/B vssd1 vssd1 vccd1 vccd1 _19853_/B sky130_fd_sc_hd__xnor2_1
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16987_ _16987_/A vssd1 vssd1 vccd1 vccd1 _16987_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18726_ _18726_/A _18726_/B vssd1 vssd1 vccd1 vccd1 _18787_/B sky130_fd_sc_hd__xor2_4
XTAP_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15938_ _26501_/Q _26373_/Q _15938_/S vssd1 vssd1 vccd1 vccd1 _15939_/B sky130_fd_sc_hd__mux2_1
XFILLER_36_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18657_ _19930_/A _19261_/B vssd1 vssd1 vccd1 vccd1 _18657_/X sky130_fd_sc_hd__or2_1
X_15869_ _17809_/A _20034_/A _15868_/Y vssd1 vssd1 vccd1 vccd1 _16040_/B sky130_fd_sc_hd__a21oi_4
XFILLER_252_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17608_ _17608_/A vssd1 vssd1 vccd1 vccd1 _17608_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18588_ _25733_/Q _25732_/Q _18588_/C vssd1 vssd1 vccd1 vccd1 _18650_/B sky130_fd_sc_hd__and3_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17539_ _17548_/A _17539_/B vssd1 vssd1 vccd1 vccd1 _25568_/D sky130_fd_sc_hd__nor2_1
XFILLER_269_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20550_ _23731_/A vssd1 vssd1 vccd1 vccd1 _20550_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_220_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19209_ _18554_/X _19207_/X _19208_/Y vssd1 vssd1 vccd1 vccd1 _19209_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20481_ _19748_/X _20480_/Y _19755_/X vssd1 vssd1 vccd1 vccd1 _20481_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_158_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22220_ _26188_/Q _22201_/X _22206_/X _22219_/X _22203_/X vssd1 vssd1 vccd1 vccd1
+ _22220_/X sky130_fd_sc_hd__a221o_1
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22151_ _26169_/Q _22136_/X _22150_/X _22148_/X vssd1 vssd1 vccd1 vccd1 _26169_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_161_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput420 _25955_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[19] sky130_fd_sc_hd__buf_2
XFILLER_279_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput431 _25965_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[29] sky130_fd_sc_hd__buf_2
X_21102_ _21138_/A vssd1 vssd1 vccd1 vccd1 _21118_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput442 _25994_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_stall_o sky130_fd_sc_hd__buf_2
Xoutput453 _25736_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[12] sky130_fd_sc_hd__buf_2
X_22082_ _26149_/Q _20939_/X _22088_/S vssd1 vssd1 vccd1 vccd1 _22083_/A sky130_fd_sc_hd__mux2_1
Xoutput464 _25746_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[22] sky130_fd_sc_hd__buf_2
Xoutput475 _25727_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[3] sky130_fd_sc_hd__buf_2
X_21033_ _25886_/Q _20926_/X _21037_/S vssd1 vssd1 vccd1 vccd1 _21034_/A sky130_fd_sc_hd__mux2_1
Xoutput486 _17057_/X vssd1 vssd1 vccd1 vccd1 wmask0[2] sky130_fd_sc_hd__buf_2
X_25910_ _27122_/CLK _25910_/D vssd1 vssd1 vccd1 vccd1 _25910_/Q sky130_fd_sc_hd__dfxtp_4
X_26890_ _27278_/CLK _26890_/D vssd1 vssd1 vccd1 vccd1 _26890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25841_ _27307_/CLK _25841_/D vssd1 vssd1 vccd1 vccd1 _25841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22984_ _26465_/Q _22672_/X _22984_/S vssd1 vssd1 vccd1 vccd1 _22985_/A sky130_fd_sc_hd__mux2_1
X_25772_ _27277_/CLK _25772_/D vssd1 vssd1 vccd1 vccd1 _25772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24723_ _24723_/A vssd1 vssd1 vccd1 vccd1 _24742_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_271_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21935_ _21946_/A vssd1 vssd1 vccd1 vccd1 _21944_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_55_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21866_ _17482_/A _21866_/B _21866_/C vssd1 vssd1 vccd1 vccd1 _21885_/B sky130_fd_sc_hd__and3b_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24654_ _24654_/A _24654_/B vssd1 vssd1 vccd1 vccd1 _24654_/Y sky130_fd_sc_hd__nand2_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20817_ _20817_/A vssd1 vssd1 vccd1 vccd1 _25804_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23605_ _23605_/A vssd1 vssd1 vccd1 vccd1 _26713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21797_ _26029_/Q _20866_/X _21805_/S vssd1 vssd1 vccd1 vccd1 _21798_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24585_ _24585_/A _24595_/B vssd1 vssd1 vccd1 vccd1 _24585_/Y sky130_fd_sc_hd__nand2_1
XFILLER_196_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26324_ _26326_/CLK _26324_/D vssd1 vssd1 vccd1 vccd1 _26324_/Q sky130_fd_sc_hd__dfxtp_2
X_20748_ _20546_/X _25771_/Q _20750_/S vssd1 vssd1 vccd1 vccd1 _20749_/A sky130_fd_sc_hd__mux2_1
X_23536_ _23536_/A vssd1 vssd1 vccd1 vccd1 _23536_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_195_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26255_ _26257_/CLK _26255_/D vssd1 vssd1 vccd1 vccd1 _26255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23467_ _26665_/Q _23079_/X _23469_/S vssd1 vssd1 vccd1 vccd1 _23468_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20679_ _20679_/A _20683_/B vssd1 vssd1 vccd1 vccd1 _20679_/X sky130_fd_sc_hd__or2_1
XFILLER_149_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13220_ _13284_/A vssd1 vssd1 vccd1 vccd1 _13221_/A sky130_fd_sc_hd__clkbuf_2
X_22418_ _22459_/A vssd1 vssd1 vccd1 vccd1 _22418_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25206_ _25218_/A _25206_/B _25206_/C _25206_/D vssd1 vssd1 vccd1 vccd1 _25228_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_195_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26186_ _26186_/CLK _26186_/D vssd1 vssd1 vccd1 vccd1 _26186_/Q sky130_fd_sc_hd__dfxtp_1
X_23398_ _23398_/A vssd1 vssd1 vccd1 vccd1 _26634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13151_ _26339_/Q _26599_/Q _15555_/S vssd1 vssd1 vccd1 vccd1 _13151_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22349_ _22335_/Y _22346_/X _22347_/X _22348_/X vssd1 vssd1 vccd1 vccd1 _26228_/D
+ sky130_fd_sc_hd__o211a_1
X_25137_ _25137_/A vssd1 vssd1 vccd1 vccd1 _25137_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13082_ _13082_/A vssd1 vssd1 vccd1 vccd1 _13083_/A sky130_fd_sc_hd__clkbuf_2
X_25068_ _24690_/Y _25043_/X _25067_/Y _25055_/X vssd1 vssd1 vccd1 vccd1 _25068_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_112_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24019_ _24019_/A vssd1 vssd1 vccd1 vccd1 _26881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16910_ _16910_/A vssd1 vssd1 vccd1 vccd1 _16910_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17890_ _14567_/A _17851_/B _17990_/A vssd1 vssd1 vccd1 vccd1 _17890_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16841_ _16910_/A _16841_/B vssd1 vssd1 vccd1 vccd1 _16940_/A sky130_fd_sc_hd__or2_1
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19560_ _19551_/X _19340_/X _19559_/X _19555_/X vssd1 vssd1 vccd1 vccd1 _25657_/D
+ sky130_fd_sc_hd__o211a_1
X_16772_ _25684_/Q vssd1 vssd1 vccd1 vccd1 _22522_/A sky130_fd_sc_hd__buf_2
XFILLER_219_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13984_ _25698_/Q _15820_/B _15716_/S vssd1 vssd1 vccd1 vccd1 _13984_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18511_ _19896_/B _18508_/X _18509_/X _27174_/Q _18510_/X vssd1 vssd1 vccd1 vccd1
+ _18511_/X sky130_fd_sc_hd__a221o_1
XFILLER_246_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15723_ _12769_/A _26891_/Q _26763_/Q _15807_/S vssd1 vssd1 vccd1 vccd1 _15723_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19491_ _25631_/Q _19497_/B vssd1 vssd1 vccd1 vccd1 _19491_/X sky130_fd_sc_hd__or2_1
X_12935_ _14031_/A vssd1 vssd1 vccd1 vccd1 _17592_/B sky130_fd_sc_hd__clkbuf_4
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18442_ _25507_/Q _18439_/X _18441_/X _25539_/Q vssd1 vssd1 vccd1 vccd1 _18442_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _15652_/X _15653_/X _16079_/S vssd1 vssd1 vccd1 vccd1 _15654_/X sky130_fd_sc_hd__mux2_1
XFILLER_234_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12866_ _12866_/A _12866_/B vssd1 vssd1 vccd1 vccd1 _12866_/X sky130_fd_sc_hd__and2_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _16292_/B vssd1 vssd1 vccd1 vccd1 _16409_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18373_ _18366_/X _18372_/X _14128_/B vssd1 vssd1 vccd1 vccd1 _18373_/X sky130_fd_sc_hd__a21o_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _26505_/Q _26377_/Q _15596_/S vssd1 vssd1 vccd1 vccd1 _15586_/B sky130_fd_sc_hd__mux2_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _12992_/A vssd1 vssd1 vccd1 vccd1 _13309_/A sky130_fd_sc_hd__buf_4
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _25528_/Q _17324_/B vssd1 vssd1 vccd1 vccd1 _17331_/C sky130_fd_sc_hd__and2_1
X_14536_ _26652_/Q _25692_/Q _14536_/S vssd1 vssd1 vccd1 vccd1 _14536_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17255_ _25506_/Q _17252_/A _17254_/Y vssd1 vssd1 vccd1 vccd1 _25506_/D sky130_fd_sc_hd__o21a_1
XFILLER_105_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14467_ _26621_/Q _26717_/Q _14474_/S vssd1 vssd1 vccd1 vccd1 _14468_/B sky130_fd_sc_hd__mux2_1
XFILLER_175_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16206_ _17791_/A _16206_/B vssd1 vssd1 vccd1 vccd1 _16206_/Y sky130_fd_sc_hd__nand2_1
X_13418_ _25807_/Q _15555_/S _13402_/A _13417_/X vssd1 vssd1 vccd1 vccd1 _13418_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17186_ _20978_/A vssd1 vssd1 vccd1 vccd1 _20657_/A sky130_fd_sc_hd__buf_4
XFILLER_155_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14398_ _25726_/Q _14560_/S vssd1 vssd1 vccd1 vccd1 _14398_/X sky130_fd_sc_hd__or2_2
XFILLER_143_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16137_ _16241_/S _16134_/X _16136_/X _15020_/A vssd1 vssd1 vccd1 vccd1 _16137_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_128_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13349_ _13835_/A vssd1 vssd1 vccd1 vccd1 _13488_/A sky130_fd_sc_hd__buf_2
XFILLER_142_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16068_ _16066_/X _16067_/X _16079_/S vssd1 vssd1 vccd1 vccd1 _16068_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15019_ _15019_/A vssd1 vssd1 vccd1 vccd1 _15020_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_130_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19827_ _19661_/X _19825_/X _19771_/X _20641_/A vssd1 vssd1 vccd1 vccd1 _19829_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19758_ _22480_/B vssd1 vssd1 vccd1 vccd1 _19758_/X sky130_fd_sc_hd__buf_4
XFILLER_272_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18709_ _19946_/A _18843_/D vssd1 vssd1 vccd1 vccd1 _18710_/B sky130_fd_sc_hd__or2_1
XFILLER_204_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19689_ _20000_/A vssd1 vssd1 vccd1 vccd1 _19820_/S sky130_fd_sc_hd__buf_2
XFILLER_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21720_ _22817_/C _22817_/A _25478_/Q vssd1 vssd1 vccd1 vccd1 _23139_/A sky130_fd_sc_hd__or3b_4
XFILLER_262_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21651_ _25968_/Q vssd1 vssd1 vccd1 vccd1 _21651_/Y sky130_fd_sc_hd__inv_2
XFILLER_224_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20602_ _20601_/X _25718_/Q _20614_/S vssd1 vssd1 vccd1 vccd1 _20603_/A sky130_fd_sc_hd__mux2_1
X_24370_ _25600_/Q _21872_/X _24370_/S vssd1 vssd1 vccd1 vccd1 _24649_/B sky130_fd_sc_hd__mux2_4
XFILLER_33_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21582_ _21552_/X _21566_/X _21580_/Y _21581_/X vssd1 vssd1 vccd1 vccd1 _21582_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_149_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23321_ _23321_/A vssd1 vssd1 vccd1 vccd1 _26600_/D sky130_fd_sc_hd__clkbuf_1
X_20533_ _23718_/A vssd1 vssd1 vccd1 vccd1 _20533_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_166_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26040_ _26599_/CLK _26040_/D vssd1 vssd1 vccd1 vccd1 _26040_/Q sky130_fd_sc_hd__dfxtp_4
X_23252_ _23252_/A vssd1 vssd1 vccd1 vccd1 _26569_/D sky130_fd_sc_hd__clkbuf_1
X_20464_ _25691_/Q vssd1 vssd1 vccd1 vccd1 _22535_/A sky130_fd_sc_hd__inv_2
XFILLER_118_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22203_ _22203_/A vssd1 vssd1 vccd1 vccd1 _22203_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23183_ _26539_/Q _23098_/X _23183_/S vssd1 vssd1 vccd1 vccd1 _23184_/A sky130_fd_sc_hd__mux2_1
X_20395_ _25688_/Q vssd1 vssd1 vccd1 vccd1 _20420_/B sky130_fd_sc_hd__buf_2
XFILLER_133_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22134_ _26163_/Q _22122_/X _22124_/X input257/X _22118_/X vssd1 vssd1 vccd1 vccd1
+ _22134_/X sky130_fd_sc_hd__a221o_1
XFILLER_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26942_ _26980_/CLK _26942_/D vssd1 vssd1 vccd1 vccd1 _26942_/Q sky130_fd_sc_hd__dfxtp_1
X_22065_ _22065_/A vssd1 vssd1 vccd1 vccd1 _26141_/D sky130_fd_sc_hd__clkbuf_1
Xoutput294 _16991_/X vssd1 vssd1 vccd1 vccd1 addr1[0] sky130_fd_sc_hd__buf_2
XINSDIODE2_1 _18613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21016_ _21016_/A vssd1 vssd1 vccd1 vccd1 _25878_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26873_ _27324_/CLK _26873_/D vssd1 vssd1 vccd1 vccd1 _26873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25824_ _25824_/CLK _25824_/D vssd1 vssd1 vccd1 vccd1 _25824_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_74_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25755_ _26292_/CLK _25755_/D vssd1 vssd1 vccd1 vccd1 _25755_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22967_ _26457_/Q _22647_/X _22973_/S vssd1 vssd1 vccd1 vccd1 _22968_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ _18076_/A vssd1 vssd1 vccd1 vccd1 _17995_/A sky130_fd_sc_hd__buf_4
X_24706_ _24706_/A vssd1 vssd1 vccd1 vccd1 _24725_/A sky130_fd_sc_hd__buf_2
X_21918_ _20542_/X _26076_/Q _21922_/S vssd1 vssd1 vccd1 vccd1 _21919_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25686_ _26286_/CLK _25686_/D vssd1 vssd1 vccd1 vccd1 _25686_/Q sky130_fd_sc_hd__dfxtp_1
X_22898_ _22898_/A vssd1 vssd1 vccd1 vccd1 _26426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24637_ _25119_/A vssd1 vssd1 vccd1 vccd1 _25065_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_230_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21849_ _26053_/Q _20948_/X _21849_/S vssd1 vssd1 vccd1 vccd1 _21850_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15370_ _14622_/A _15353_/X _15360_/X _15369_/X _14682_/A vssd1 vssd1 vccd1 vccd1
+ _15370_/X sky130_fd_sc_hd__a311o_1
X_24568_ _27043_/Q _24562_/X _24565_/Y _24567_/X vssd1 vssd1 vccd1 vccd1 _27043_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26307_ _26307_/CLK _26307_/D vssd1 vssd1 vccd1 vccd1 _26307_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_184_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14321_ _14403_/A _14321_/B vssd1 vssd1 vccd1 vccd1 _14321_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23519_ _23519_/A vssd1 vssd1 vccd1 vccd1 _26686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27287_ _27287_/CLK _27287_/D vssd1 vssd1 vccd1 vccd1 _27287_/Q sky130_fd_sc_hd__dfxtp_1
X_24499_ _24551_/A vssd1 vssd1 vccd1 vccd1 _24499_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_278_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17040_ _17035_/X _16935_/B _17039_/X input230/X vssd1 vssd1 vccd1 vccd1 _17040_/X
+ sky130_fd_sc_hd__a22o_4
X_26238_ _26238_/CLK _26238_/D vssd1 vssd1 vccd1 vccd1 _26238_/Q sky130_fd_sc_hd__dfxtp_1
X_14252_ _26331_/Q _26591_/Q _14252_/S vssd1 vssd1 vccd1 vccd1 _14252_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13203_ _20868_/B _13244_/A _13277_/A _22817_/C _13202_/X vssd1 vssd1 vccd1 vccd1
+ _13204_/C sky130_fd_sc_hd__a221oi_2
XFILLER_137_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26169_ _27264_/CLK _26169_/D vssd1 vssd1 vccd1 vccd1 _26169_/Q sky130_fd_sc_hd__dfxtp_1
X_14183_ _14440_/S _14171_/X _14175_/X _14355_/A _14182_/X vssd1 vssd1 vccd1 vccd1
+ _14183_/X sky130_fd_sc_hd__a311o_1
XFILLER_87_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_13134_ _13134_/A vssd1 vssd1 vccd1 vccd1 _13135_/A sky130_fd_sc_hd__clkbuf_4
X_18991_ _27054_/Q _18747_/X _18988_/X _18990_/X _18761_/X vssd1 vssd1 vccd1 vccd1
+ _18991_/X sky130_fd_sc_hd__o221a_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13065_ _13065_/A vssd1 vssd1 vccd1 vccd1 _15460_/S sky130_fd_sc_hd__buf_2
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17942_ _18202_/A vssd1 vssd1 vccd1 vccd1 _18210_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_215_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17873_ _17869_/X _17870_/X _18070_/S vssd1 vssd1 vccd1 vccd1 _17873_/X sky130_fd_sc_hd__mux2_2
X_19612_ _27062_/Q _19616_/B _19612_/C vssd1 vssd1 vccd1 vccd1 _19614_/C sky130_fd_sc_hd__and3_1
X_16824_ _16828_/A _16824_/B _16868_/B vssd1 vssd1 vccd1 vccd1 _16825_/A sky130_fd_sc_hd__and3_4
XFILLER_254_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19543_ _25651_/Q _19549_/B vssd1 vssd1 vccd1 vccd1 _19543_/X sky130_fd_sc_hd__or2_1
XFILLER_235_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16755_ _25678_/Q vssd1 vssd1 vccd1 vccd1 _22509_/A sky130_fd_sc_hd__buf_2
Xclkbuf_4_0_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_253_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13967_ _26070_/Q _25875_/Q _16005_/S vssd1 vssd1 vccd1 vccd1 _13967_/X sky130_fd_sc_hd__mux2_1
XFILLER_207_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15706_ _15706_/A _15706_/B _15706_/C vssd1 vssd1 vccd1 vccd1 _15706_/X sky130_fd_sc_hd__or3_1
XFILLER_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12918_ _14133_/A vssd1 vssd1 vccd1 vccd1 _17623_/B sky130_fd_sc_hd__clkbuf_2
X_19474_ _18912_/A _19472_/Y _18998_/X vssd1 vssd1 vccd1 vccd1 _19474_/X sky130_fd_sc_hd__o21a_1
X_16686_ _21190_/A vssd1 vssd1 vccd1 vccd1 _16769_/A sky130_fd_sc_hd__clkbuf_2
X_13898_ _13896_/X _13897_/X _14246_/S vssd1 vssd1 vccd1 vccd1 _13898_/X sky130_fd_sc_hd__mux2_1
XFILLER_234_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18425_ _19046_/B _19572_/B _18424_/X _18359_/X vssd1 vssd1 vccd1 vccd1 _18425_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_206_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15637_ _14870_/A _15634_/X _15636_/X _14659_/A vssd1 vssd1 vccd1 vccd1 _15637_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12849_ _25909_/Q _12899_/A _12846_/X _12891_/A _12869_/A vssd1 vssd1 vccd1 vccd1
+ _12849_/X sky130_fd_sc_hd__o221a_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18356_ _18356_/A vssd1 vssd1 vccd1 vccd1 _19289_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15568_ _15562_/X _15564_/X _15567_/X _16072_/S _12702_/A vssd1 vssd1 vccd1 vccd1
+ _15568_/X sky130_fd_sc_hd__o221a_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17307_ _25522_/Q _17305_/B _17306_/Y vssd1 vssd1 vccd1 vccd1 _25522_/D sky130_fd_sc_hd__o21a_1
X_14519_ _13083_/A _26876_/Q _26748_/Q _14332_/S vssd1 vssd1 vccd1 vccd1 _14519_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18287_ _25728_/Q _18287_/B vssd1 vssd1 vccd1 vccd1 _18288_/B sky130_fd_sc_hd__nor2_1
X_15499_ _15317_/A _15496_/X _15498_/X _15312_/A vssd1 vssd1 vccd1 vccd1 _15499_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_266_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17238_ _25176_/A vssd1 vssd1 vccd1 vccd1 _25109_/A sky130_fd_sc_hd__buf_6
XFILLER_174_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17169_ _21429_/A _17159_/X _17168_/Y _17134_/X vssd1 vssd1 vccd1 vccd1 _25482_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20180_ _27152_/Q _27086_/Q vssd1 vssd1 vccd1 vccd1 _20180_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23870_ _23870_/A vssd1 vssd1 vccd1 vccd1 _26815_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22821_ _26392_/Q _22640_/X _22829_/S vssd1 vssd1 vccd1 vccd1 _22822_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25540_ _25545_/CLK _25540_/D vssd1 vssd1 vccd1 vccd1 _25540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22752_ _26362_/Q _22650_/X _22756_/S vssd1 vssd1 vccd1 vccd1 _22753_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21703_ _25990_/Q _17456_/A _21707_/S vssd1 vssd1 vccd1 vccd1 _21704_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22683_ _26340_/Q _22682_/X _22689_/S vssd1 vssd1 vccd1 vccd1 _22684_/A sky130_fd_sc_hd__mux2_1
X_25471_ _25590_/CLK _25471_/D vssd1 vssd1 vccd1 vccd1 _25471_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_212_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27210_ _27228_/CLK _27210_/D vssd1 vssd1 vccd1 vccd1 _27210_/Q sky130_fd_sc_hd__dfxtp_1
X_24422_ _26303_/Q _24382_/X _24383_/X input216/X _24384_/X vssd1 vssd1 vccd1 vccd1
+ _24422_/X sky130_fd_sc_hd__a221o_1
X_21634_ _21276_/A _21633_/X _21603_/X vssd1 vssd1 vccd1 vccd1 _21634_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_100_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_139_wb_clk_i _25501_/CLK vssd1 vssd1 vccd1 vccd1 _25867_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_166_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27141_ _27164_/CLK _27141_/D vssd1 vssd1 vccd1 vccd1 _27141_/Q sky130_fd_sc_hd__dfxtp_1
X_21565_ _21544_/X _21564_/X _21537_/X vssd1 vssd1 vccd1 vccd1 _21565_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_178_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24353_ _24457_/A _25491_/Q _17703_/X _24989_/A _24352_/X vssd1 vssd1 vccd1 vccd1
+ _24633_/C sky130_fd_sc_hd__a2111o_1
XFILLER_60_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23304_ _23361_/S vssd1 vssd1 vccd1 vccd1 _23313_/S sky130_fd_sc_hd__clkbuf_4
X_20516_ _23530_/A vssd1 vssd1 vccd1 vccd1 _23706_/A sky130_fd_sc_hd__clkbuf_4
X_24284_ _26985_/Q _26984_/Q _24284_/C vssd1 vssd1 vccd1 vccd1 _24286_/B sky130_fd_sc_hd__and3_1
XFILLER_154_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27072_ _27176_/CLK _27072_/D vssd1 vssd1 vccd1 vccd1 _27072_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_219_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21496_ _21430_/X _19072_/X _21431_/X _25816_/Q _21483_/X vssd1 vssd1 vccd1 vccd1
+ _21496_/X sky130_fd_sc_hd__a221o_1
XFILLER_5_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23235_ _23281_/S vssd1 vssd1 vccd1 vccd1 _23244_/S sky130_fd_sc_hd__buf_6
X_26023_ _26483_/CLK _26023_/D vssd1 vssd1 vccd1 vccd1 _26023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20447_ _20448_/A _20448_/B vssd1 vssd1 vccd1 vccd1 _20471_/A sky130_fd_sc_hd__nand2_1
XFILLER_107_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23166_ _26531_/Q _23073_/X _23172_/S vssd1 vssd1 vccd1 vccd1 _23167_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20378_ _20694_/A _19698_/X _20377_/X _20357_/A vssd1 vssd1 vccd1 vccd1 _20379_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_133_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22117_ _22203_/A vssd1 vssd1 vccd1 vccd1 _22155_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_268_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23097_ _23097_/A vssd1 vssd1 vccd1 vccd1 _26506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_279_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22048_ _22048_/A vssd1 vssd1 vccd1 vccd1 _26133_/D sky130_fd_sc_hd__clkbuf_1
X_26925_ _26925_/CLK _26925_/D vssd1 vssd1 vccd1 vccd1 _26925_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26856_ _26856_/CLK _26856_/D vssd1 vssd1 vccd1 vccd1 _26856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14870_ _14870_/A vssd1 vssd1 vccd1 vccd1 _16320_/S sky130_fd_sc_hd__clkbuf_4
XTAP_5789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13821_ _13821_/A _13821_/B vssd1 vssd1 vccd1 vccd1 _13821_/X sky130_fd_sc_hd__or2_1
X_25807_ _26913_/CLK _25807_/D vssd1 vssd1 vccd1 vccd1 _25807_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_47_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26787_ _27238_/CLK _26787_/D vssd1 vssd1 vccd1 vccd1 _26787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23999_ _23999_/A vssd1 vssd1 vccd1 vccd1 _26873_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_251_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16540_ _16538_/X _16539_/X _16540_/S vssd1 vssd1 vccd1 vccd1 _16540_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_108 _21628_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13752_ _16639_/A _13750_/X _13751_/X vssd1 vssd1 vccd1 vccd1 _23536_/A sky130_fd_sc_hd__a21o_4
X_25738_ _26282_/CLK _25738_/D vssd1 vssd1 vccd1 vccd1 _25738_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_119 _23032_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_6_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_204_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12703_ _12703_/A vssd1 vssd1 vccd1 vccd1 _12704_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16471_ _12777_/A _26907_/Q _26779_/Q _16490_/B _16484_/A vssd1 vssd1 vccd1 vccd1
+ _16471_/X sky130_fd_sc_hd__a221o_1
XFILLER_245_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13683_ _13683_/A vssd1 vssd1 vccd1 vccd1 _13683_/X sky130_fd_sc_hd__clkbuf_2
X_25669_ _25670_/CLK _25669_/D vssd1 vssd1 vccd1 vccd1 _25669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18210_ _18208_/X _18209_/X _18210_/S vssd1 vssd1 vccd1 vccd1 _18210_/X sky130_fd_sc_hd__mux2_1
X_15422_ _27315_/Q _26572_/Q _15422_/S vssd1 vssd1 vccd1 vccd1 _15422_/X sky130_fd_sc_hd__mux2_1
XPHY_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19190_ _19189_/Y _16606_/Y _19453_/S vssd1 vssd1 vccd1 vccd1 _19190_/X sky130_fd_sc_hd__mux2_1
XPHY_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18141_ _19196_/A _18136_/Y _18140_/X _18035_/A _19076_/A vssd1 vssd1 vccd1 vccd1
+ _18141_/X sky130_fd_sc_hd__o32a_2
X_15353_ _16401_/S _15350_/X _15352_/X _15019_/A vssd1 vssd1 vccd1 vccd1 _15353_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14304_ _13521_/A _25761_/Q _14365_/S _26847_/Q _14390_/S vssd1 vssd1 vccd1 vccd1
+ _14304_/X sky130_fd_sc_hd__o221a_1
XFILLER_200_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18072_ _18068_/X _18071_/X _18318_/S vssd1 vssd1 vccd1 vccd1 _18073_/B sky130_fd_sc_hd__mux2_1
XFILLER_184_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15284_ _15165_/X _15282_/X _15283_/X vssd1 vssd1 vccd1 vccd1 _15285_/B sky130_fd_sc_hd__o21ai_1
XFILLER_184_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17023_ _17021_/X _16864_/B _17017_/X input217/X vssd1 vssd1 vccd1 vccd1 _17023_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14235_ _17966_/A _14570_/B vssd1 vssd1 vccd1 vccd1 _18324_/B sky130_fd_sc_hd__nor2_2
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14166_ _13614_/A _14161_/X _14165_/Y _15885_/A vssd1 vssd1 vccd1 vccd1 _14166_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13117_ _27306_/Q _26563_/Q _15540_/S vssd1 vssd1 vccd1 vccd1 _13117_/X sky130_fd_sc_hd__mux2_1
X_14097_ _13890_/A _26689_/Q _26817_/Q _15714_/A _13048_/A vssd1 vssd1 vccd1 vccd1
+ _14097_/X sky130_fd_sc_hd__a221o_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18974_ _19252_/A vssd1 vssd1 vccd1 vccd1 _19448_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_258_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13048_ _13048_/A vssd1 vssd1 vccd1 vccd1 _13049_/A sky130_fd_sc_hd__clkbuf_4
X_17925_ _18063_/S vssd1 vssd1 vccd1 vccd1 _18042_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_140_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17856_ _17856_/A _19585_/S vssd1 vssd1 vccd1 vccd1 _17856_/X sky130_fd_sc_hd__or2b_1
XFILLER_39_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16807_ _16812_/A vssd1 vssd1 vccd1 vccd1 _16810_/A sky130_fd_sc_hd__buf_2
XFILLER_281_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17787_ _17787_/A _17787_/B vssd1 vssd1 vccd1 vccd1 _17787_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14999_ _14890_/A _25786_/Q _14905_/S _26872_/Q _14917_/X vssd1 vssd1 vccd1 vccd1
+ _14999_/X sky130_fd_sc_hd__o221a_1
XFILLER_281_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19526_ _19552_/A vssd1 vssd1 vccd1 vccd1 _19536_/B sky130_fd_sc_hd__clkbuf_1
X_16738_ _22494_/A _16726_/X _16727_/X _18678_/A vssd1 vssd1 vccd1 vccd1 _16738_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_241_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19457_ _16550_/A _17997_/A _19455_/X vssd1 vssd1 vccd1 vccd1 _19457_/X sky130_fd_sc_hd__a21o_1
X_16669_ _16669_/A _16669_/B vssd1 vssd1 vccd1 vccd1 _21198_/A sky130_fd_sc_hd__nand2_4
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18408_ _19256_/A _18357_/A _18376_/X _18407_/X vssd1 vssd1 vccd1 vccd1 _18408_/X
+ sky130_fd_sc_hd__a211o_1
X_19388_ _19388_/A _19423_/B vssd1 vssd1 vccd1 vccd1 _19388_/X sky130_fd_sc_hd__or2_1
XFILLER_188_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18339_ _18339_/A vssd1 vssd1 vccd1 vccd1 _18340_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_187_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21350_ _21350_/A vssd1 vssd1 vccd1 vccd1 _21350_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20301_ _20301_/A _20302_/A vssd1 vssd1 vccd1 vccd1 _20301_/Y sky130_fd_sc_hd__nor2_1
X_21281_ _21559_/B vssd1 vssd1 vccd1 vccd1 _21332_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23020_ _26481_/Q _22723_/X _23028_/S vssd1 vssd1 vccd1 vccd1 _23021_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20232_ _20305_/A _20260_/B _20300_/B vssd1 vssd1 vccd1 vccd1 _20232_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_150_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20163_ _22509_/A _20078_/X _20155_/X _20162_/X _20076_/X vssd1 vssd1 vccd1 vccd1
+ _25678_/D sky130_fd_sc_hd__o221a_1
XFILLER_249_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24971_ _27157_/Q _24953_/X _24969_/Y _24970_/X vssd1 vssd1 vccd1 vccd1 _27157_/D
+ sky130_fd_sc_hd__o211a_1
X_20094_ _25740_/Q _20355_/A _20093_/X _20119_/B vssd1 vssd1 vccd1 vccd1 _20095_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_58_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26710_ _27322_/CLK _26710_/D vssd1 vssd1 vccd1 vccd1 _26710_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23922_ _23773_/X _26839_/Q _23926_/S vssd1 vssd1 vccd1 vccd1 _23923_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26641_ _27316_/CLK _26641_/D vssd1 vssd1 vccd1 vccd1 _26641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23853_ _23853_/A vssd1 vssd1 vccd1 vccd1 _26808_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22804_ _22804_/A vssd1 vssd1 vccd1 vccd1 _26385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26572_ _27315_/CLK _26572_/D vssd1 vssd1 vccd1 vccd1 _26572_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20996_ _25869_/Q _20866_/X _21004_/S vssd1 vssd1 vccd1 vccd1 _20997_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23784_ _23784_/A vssd1 vssd1 vccd1 vccd1 _26778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_260_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25523_ _25985_/CLK _25523_/D vssd1 vssd1 vccd1 vccd1 _25523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22735_ _22735_/A vssd1 vssd1 vccd1 vccd1 _26356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25454_ _25454_/A vssd1 vssd1 vccd1 vccd1 _27321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22666_ _23709_/A vssd1 vssd1 vccd1 vccd1 _22666_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24405_ _26300_/Q _21881_/X _21883_/X input244/X _24404_/X vssd1 vssd1 vccd1 vccd1
+ _24405_/X sky130_fd_sc_hd__a221o_1
XFILLER_185_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21617_ _21354_/A _21566_/X _21616_/Y _21581_/X vssd1 vssd1 vccd1 vccd1 _21617_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_200_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25385_ _27291_/Q _23776_/A _25387_/S vssd1 vssd1 vccd1 vccd1 _25386_/A sky130_fd_sc_hd__mux2_1
X_22597_ _26314_/Q _22604_/B vssd1 vssd1 vccd1 vccd1 _22597_/Y sky130_fd_sc_hd__nand2_1
X_27124_ _27130_/CLK _27124_/D vssd1 vssd1 vccd1 vccd1 _27124_/Q sky130_fd_sc_hd__dfxtp_4
X_24336_ _27003_/Q _24334_/B _24335_/Y vssd1 vssd1 vccd1 vccd1 _27003_/D sky130_fd_sc_hd__o21a_1
XFILLER_127_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21548_ _21509_/X _19207_/X _21510_/X _25820_/Q _21547_/X vssd1 vssd1 vccd1 vccd1
+ _21548_/X sky130_fd_sc_hd__a221o_1
XFILLER_217_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27055_ _27062_/CLK _27055_/D vssd1 vssd1 vccd1 vccd1 _27055_/Q sky130_fd_sc_hd__dfxtp_2
X_24267_ _24285_/A _24267_/B _24268_/B vssd1 vssd1 vccd1 vccd1 _26979_/D sky130_fd_sc_hd__nor3_1
X_21479_ _25953_/Q _21443_/X _21478_/Y _21467_/X vssd1 vssd1 vccd1 vccd1 _25953_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_4_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26006_ _27307_/CLK _26006_/D vssd1 vssd1 vccd1 vccd1 _26006_/Q sky130_fd_sc_hd__dfxtp_2
X_14020_ _13636_/B _16830_/B _14019_/X _15948_/B vssd1 vssd1 vccd1 vccd1 _17798_/A
+ sky130_fd_sc_hd__o211a_1
X_23218_ _26554_/Q _23044_/X _23222_/S vssd1 vssd1 vccd1 vccd1 _23219_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24198_ _24216_/A _24203_/C vssd1 vssd1 vccd1 vccd1 _24198_/Y sky130_fd_sc_hd__nor2_1
XFILLER_150_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23149_ _23149_/A vssd1 vssd1 vccd1 vccd1 _26523_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27304_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_268_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15971_ _27275_/Q _26468_/Q _15971_/S vssd1 vssd1 vccd1 vccd1 _15971_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17710_ _18116_/A _17735_/A _17735_/B vssd1 vssd1 vccd1 vccd1 _17711_/C sky130_fd_sc_hd__nor3_1
XTAP_5553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26908_ _26908_/CLK _26908_/D vssd1 vssd1 vccd1 vccd1 _26908_/Q sky130_fd_sc_hd__dfxtp_2
X_14922_ _27292_/Q _26485_/Q _14996_/S vssd1 vssd1 vccd1 vccd1 _14922_/X sky130_fd_sc_hd__mux2_1
XTAP_5564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18690_ _19196_/A vssd1 vssd1 vccd1 vccd1 _19482_/B sky130_fd_sc_hd__buf_2
XTAP_5575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17641_ _17650_/A _17641_/B vssd1 vssd1 vccd1 vccd1 _25592_/D sky130_fd_sc_hd__nor2_1
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26839_ _26932_/CLK _26839_/D vssd1 vssd1 vccd1 vccd1 _26839_/Q sky130_fd_sc_hd__dfxtp_1
X_14853_ _16384_/S vssd1 vssd1 vccd1 vccd1 _14876_/S sky130_fd_sc_hd__clkbuf_2
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _13802_/X _13558_/A _13578_/X _25605_/Q _13803_/X vssd1 vssd1 vccd1 vccd1
+ _23533_/A sky130_fd_sc_hd__a221o_4
XFILLER_17_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17572_ _19636_/A vssd1 vssd1 vccd1 vccd1 _17572_/X sky130_fd_sc_hd__clkbuf_1
X_14784_ _16513_/A _26126_/Q _26027_/Q _14767_/S _14773_/A vssd1 vssd1 vccd1 vccd1
+ _14784_/X sky130_fd_sc_hd__a221o_1
XFILLER_251_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19311_ _18947_/A _19309_/Y _18998_/A vssd1 vssd1 vccd1 vccd1 _19311_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16523_ _26127_/Q _26028_/Q _16523_/S vssd1 vssd1 vccd1 vccd1 _16523_/X sky130_fd_sc_hd__mux2_1
XFILLER_232_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13735_ _13704_/X _13717_/X _13734_/X vssd1 vssd1 vccd1 vccd1 _13735_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19242_ _18602_/X _18495_/B _18497_/X _18597_/X _19241_/X vssd1 vssd1 vccd1 vccd1
+ _19242_/X sky130_fd_sc_hd__o221a_1
XFILLER_149_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16454_ _19322_/A _16454_/B vssd1 vssd1 vccd1 vccd1 _17846_/D sky130_fd_sc_hd__nor2_1
X_13666_ _15588_/A _25838_/Q _26038_/Q _15915_/S _13644_/X vssd1 vssd1 vccd1 vccd1
+ _13666_/X sky130_fd_sc_hd__a221o_1
X_15405_ _15318_/X _15400_/X _15404_/X _15313_/X vssd1 vssd1 vccd1 vccd1 _15405_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19173_ _20252_/A _19442_/B vssd1 vssd1 vccd1 vccd1 _19173_/Y sky130_fd_sc_hd__nor2_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ _26515_/Q _26387_/Q _16385_/S vssd1 vssd1 vccd1 vccd1 _16385_/X sky130_fd_sc_hd__mux2_1
X_13597_ _26917_/Q _26401_/Q _15971_/S vssd1 vssd1 vccd1 vccd1 _13597_/X sky130_fd_sc_hd__mux2_1
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18124_ _18458_/A vssd1 vssd1 vccd1 vccd1 _18568_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15336_ _14807_/A _15319_/X _15325_/X _15335_/X _14786_/A vssd1 vssd1 vccd1 vccd1
+ _15336_/X sky130_fd_sc_hd__a311o_1
XFILLER_185_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18055_ _18598_/S vssd1 vssd1 vccd1 vccd1 _18684_/S sky130_fd_sc_hd__clkbuf_2
X_15267_ _26086_/Q _16134_/S _15265_/X _15266_/X vssd1 vssd1 vccd1 vccd1 _15267_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17006_ _17016_/A vssd1 vssd1 vccd1 vccd1 _17006_/X sky130_fd_sc_hd__clkbuf_2
X_14218_ _13937_/X _25762_/Q _15759_/S _26848_/Q _14309_/S vssd1 vssd1 vccd1 vccd1
+ _14218_/X sky130_fd_sc_hd__o221a_1
XFILLER_126_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15198_ _16259_/S vssd1 vssd1 vccd1 vccd1 _16255_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_113_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14149_ _26100_/Q _26001_/Q _14265_/S vssd1 vssd1 vccd1 vccd1 _14149_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_258_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18957_ _17287_/X _18559_/A _18954_/X _18956_/X _18574_/A vssd1 vssd1 vccd1 vccd1
+ _18957_/X sky130_fd_sc_hd__o221a_1
XFILLER_98_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17908_ _17906_/X _17907_/X _18070_/S vssd1 vssd1 vccd1 vccd1 _17908_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18888_ _19455_/C _18720_/X _18886_/Y _18887_/Y _18788_/X vssd1 vssd1 vccd1 vccd1
+ _18888_/X sky130_fd_sc_hd__a221o_4
XFILLER_39_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17839_ _18978_/A _17837_/X _17838_/X vssd1 vssd1 vccd1 vccd1 _17839_/X sky130_fd_sc_hd__o21a_1
XFILLER_187_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20850_ _25821_/Q vssd1 vssd1 vccd1 vccd1 _20851_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_282_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19509_ _19499_/X _18576_/X _19508_/X _19502_/X vssd1 vssd1 vccd1 vccd1 _25638_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_212_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20781_ _20609_/X _25786_/Q _20783_/S vssd1 vssd1 vccd1 vccd1 _20782_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_450 _17054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_461 _18969_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_472 _22533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22520_ _22520_/A _22524_/B vssd1 vssd1 vccd1 vccd1 _22521_/A sky130_fd_sc_hd__and2_1
XFILLER_195_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_483 _19728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_494 _16681_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22451_ _26204_/Q _22446_/X _22450_/X _22442_/X vssd1 vssd1 vccd1 vccd1 _26252_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21402_ _25480_/Q _21416_/B vssd1 vssd1 vccd1 vccd1 _21402_/X sky130_fd_sc_hd__or2_1
X_22382_ _22390_/A vssd1 vssd1 vccd1 vccd1 _22405_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25170_ _27198_/Q _25137_/X _25169_/X vssd1 vssd1 vccd1 vccd1 _27198_/D sky130_fd_sc_hd__o21ba_1
XFILLER_157_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21333_ _21284_/X _18524_/X _21286_/X _25804_/Q _21322_/X vssd1 vssd1 vccd1 vccd1
+ _21333_/X sky130_fd_sc_hd__a221o_1
X_24121_ _24121_/A vssd1 vssd1 vccd1 vccd1 _26927_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21264_ _21264_/A vssd1 vssd1 vccd1 vccd1 _21873_/A sky130_fd_sc_hd__buf_2
X_24052_ _24052_/A vssd1 vssd1 vccd1 vccd1 _26896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23003_ _23003_/A vssd1 vssd1 vccd1 vccd1 _26473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20215_ _27153_/Q _27087_/Q vssd1 vssd1 vccd1 vccd1 _20218_/B sky130_fd_sc_hd__nor2_1
XFILLER_278_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21195_ _21195_/A _21195_/B _21195_/C vssd1 vssd1 vccd1 vccd1 _21195_/Y sky130_fd_sc_hd__nor3_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20146_ _20118_/B _20126_/A _20145_/X vssd1 vssd1 vccd1 vccd1 _20148_/B sky130_fd_sc_hd__a21oi_1
XFILLER_265_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24954_ _24954_/A vssd1 vssd1 vccd1 vccd1 _24972_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_20077_ _22502_/A _19876_/X _20068_/X _20075_/X _20076_/X vssd1 vssd1 vccd1 vccd1
+ _25675_/D sky130_fd_sc_hd__o221a_1
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23905_ _23905_/A vssd1 vssd1 vccd1 vccd1 _26831_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24885_ _20694_/A _19963_/X _25151_/A _24779_/A vssd1 vssd1 vccd1 vccd1 _24885_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_261_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26624_ _26880_/CLK _26624_/D vssd1 vssd1 vccd1 vccd1 _26624_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23836_ _23836_/A vssd1 vssd1 vccd1 vccd1 _26800_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_154_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27087_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26555_ _27298_/CLK _26555_/D vssd1 vssd1 vccd1 vccd1 _26555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_260_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23767_ _23767_/A vssd1 vssd1 vccd1 vccd1 _23780_/S sky130_fd_sc_hd__buf_6
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20979_ _20986_/C vssd1 vssd1 vccd1 vccd1 _25867_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_214_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13520_ _13520_/A vssd1 vssd1 vccd1 vccd1 _13521_/A sky130_fd_sc_hd__clkbuf_2
X_25506_ _27014_/CLK _25506_/D vssd1 vssd1 vccd1 vccd1 _25506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22718_ _26351_/Q _22717_/X _22721_/S vssd1 vssd1 vccd1 vccd1 _22719_/A sky130_fd_sc_hd__mux2_1
X_26486_ _27326_/CLK _26486_/D vssd1 vssd1 vccd1 vccd1 _26486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23698_ _23698_/A vssd1 vssd1 vccd1 vccd1 _26751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13451_ _13711_/A _13451_/B vssd1 vssd1 vccd1 vccd1 _13451_/Y sky130_fd_sc_hd__nand2_1
X_25437_ _23747_/X _27314_/Q _25437_/S vssd1 vssd1 vccd1 vccd1 _25438_/A sky130_fd_sc_hd__mux2_1
X_22649_ _22649_/A vssd1 vssd1 vccd1 vccd1 _26329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16170_ _16170_/A _16921_/A vssd1 vssd1 vccd1 vccd1 _16170_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13382_ _17824_/A _13380_/Y _13381_/Y vssd1 vssd1 vccd1 vccd1 _17817_/D sky130_fd_sc_hd__a21o_1
X_25368_ _27283_/Q _23750_/A _25376_/S vssd1 vssd1 vccd1 vccd1 _25369_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15121_ _26678_/Q _25718_/Q _15121_/S vssd1 vssd1 vccd1 vccd1 _15121_/X sky130_fd_sc_hd__mux2_1
X_27107_ _27110_/CLK _27107_/D vssd1 vssd1 vccd1 vccd1 _27107_/Q sky130_fd_sc_hd__dfxtp_2
X_24319_ _24327_/A _24319_/B _24320_/B vssd1 vssd1 vccd1 vccd1 _26997_/D sky130_fd_sc_hd__nor3_1
XFILLER_182_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25299_ _25299_/A vssd1 vssd1 vccd1 vccd1 _27252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27038_ _27044_/CLK _27038_/D vssd1 vssd1 vccd1 vccd1 _27038_/Q sky130_fd_sc_hd__dfxtp_1
X_15052_ _15351_/B vssd1 vssd1 vccd1 vccd1 _16380_/B sky130_fd_sc_hd__buf_6
XFILLER_182_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14003_ _13135_/A _14000_/X _14002_/X _13857_/X vssd1 vssd1 vccd1 vccd1 _14003_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_141_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19860_ _19860_/A _19860_/B vssd1 vssd1 vccd1 vccd1 _19860_/X sky130_fd_sc_hd__or2_1
X_18811_ _18811_/A vssd1 vssd1 vccd1 vccd1 _18811_/X sky130_fd_sc_hd__clkbuf_2
X_19791_ _19683_/X _19789_/Y _19790_/X _19651_/X vssd1 vssd1 vccd1 vccd1 _19791_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_284_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18742_ _18806_/A vssd1 vssd1 vccd1 vccd1 _18742_/X sky130_fd_sc_hd__clkbuf_2
X_15954_ _15954_/A _15954_/B _15954_/C vssd1 vssd1 vccd1 vccd1 _15954_/X sky130_fd_sc_hd__or3_1
XTAP_5350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput150 dout1[49] vssd1 vssd1 vccd1 vccd1 input150/X sky130_fd_sc_hd__clkbuf_2
XTAP_5361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_283_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput161 dout1[59] vssd1 vssd1 vccd1 vccd1 input161/X sky130_fd_sc_hd__clkbuf_2
XTAP_5372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput172 irq[10] vssd1 vssd1 vccd1 vccd1 _19613_/C sky130_fd_sc_hd__buf_4
X_14905_ _26681_/Q _25721_/Q _14905_/S vssd1 vssd1 vccd1 vccd1 _14905_/X sky130_fd_sc_hd__mux2_1
XTAP_5394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18673_ _18673_/A vssd1 vssd1 vccd1 vccd1 _25608_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15885_ _15885_/A _15885_/B _15885_/C vssd1 vssd1 vccd1 vccd1 _15885_/X sky130_fd_sc_hd__or3_1
Xinput183 irq[6] vssd1 vssd1 vccd1 vccd1 input183/X sky130_fd_sc_hd__clkbuf_8
XFILLER_36_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput194 localMemory_wb_adr_i[13] vssd1 vssd1 vccd1 vccd1 input194/X sky130_fd_sc_hd__clkbuf_1
XFILLER_236_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14836_ _25659_/Q _24351_/B _14613_/X vssd1 vssd1 vccd1 vccd1 _14836_/X sky130_fd_sc_hd__a21o_1
X_17624_ _25925_/Q _17544_/X _17623_/X vssd1 vssd1 vccd1 vccd1 _17624_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_251_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _17653_/A vssd1 vssd1 vccd1 vccd1 _17592_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14767_ _26650_/Q _26746_/Q _14767_/S vssd1 vssd1 vccd1 vccd1 _14767_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16506_ _16488_/X _16505_/X _14593_/X vssd1 vssd1 vccd1 vccd1 _16506_/X sky130_fd_sc_hd__a21o_1
X_13718_ _27271_/Q _26464_/Q _16067_/S vssd1 vssd1 vccd1 vccd1 _13718_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17486_ _17486_/A vssd1 vssd1 vccd1 vccd1 _21208_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14698_ _25859_/Q _26059_/Q _14699_/S vssd1 vssd1 vccd1 vccd1 _14698_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19225_ _27029_/Q _18514_/A _19224_/X _18455_/A vssd1 vssd1 vccd1 vccd1 _19225_/X
+ sky130_fd_sc_hd__a22o_1
X_16437_ _15321_/X _25856_/Q _26056_/Q _15209_/S _15210_/X vssd1 vssd1 vccd1 vccd1
+ _16437_/X sky130_fd_sc_hd__a221o_1
XFILLER_258_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13649_ _12738_/D _26597_/Q _15931_/S _26337_/Q _14223_/S vssd1 vssd1 vccd1 vccd1
+ _13649_/X sky130_fd_sc_hd__o221a_1
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19156_ _19156_/A _19156_/B vssd1 vssd1 vccd1 vccd1 _19183_/B sky130_fd_sc_hd__xnor2_4
X_16368_ _20690_/A _19268_/A _16368_/S vssd1 vssd1 vccd1 vccd1 _17783_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18107_ _18391_/A vssd1 vssd1 vccd1 vccd1 _19058_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15319_ _15313_/X _15314_/X _15316_/X _15318_/X vssd1 vssd1 vccd1 vccd1 _15319_/X
+ sky130_fd_sc_hd__a211o_1
X_19087_ _19087_/A vssd1 vssd1 vccd1 vccd1 _19087_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16299_ _15065_/X _26417_/Q _16324_/S _16298_/X vssd1 vssd1 vccd1 vccd1 _16299_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18038_ _18184_/B _19290_/A vssd1 vssd1 vccd1 vccd1 _18038_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20000_ _20000_/A vssd1 vssd1 vccd1 vccd1 _20219_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_114_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19989_ _27113_/Q _19877_/X _19967_/X _19988_/Y vssd1 vssd1 vccd1 vccd1 _19989_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21951_ _20605_/X _26091_/Q _21955_/S vssd1 vssd1 vccd1 vccd1 _21952_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20902_ _20902_/A vssd1 vssd1 vccd1 vccd1 _25838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_255_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24670_ _24678_/A _24670_/B vssd1 vssd1 vccd1 vccd1 _27075_/D sky130_fd_sc_hd__nor2_1
X_21882_ _24456_/A vssd1 vssd1 vccd1 vccd1 _24474_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_254_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23621_ _26719_/Q _23520_/X _23623_/S vssd1 vssd1 vccd1 vccd1 _23622_/A sky130_fd_sc_hd__mux2_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20833_ _20833_/A vssd1 vssd1 vccd1 vccd1 _25812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26340_ _26468_/CLK _26340_/D vssd1 vssd1 vccd1 vccd1 _26340_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_196_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23552_ _23552_/A vssd1 vssd1 vccd1 vccd1 _23552_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20764_ _20575_/X _25778_/Q _20772_/S vssd1 vssd1 vccd1 vccd1 _20765_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_280 _25810_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_291 _25821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22503_ _22503_/A vssd1 vssd1 vccd1 vccd1 _26276_/D sky130_fd_sc_hd__clkbuf_1
X_26271_ _26271_/CLK _26271_/D vssd1 vssd1 vccd1 vccd1 _26271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20695_ _26288_/Q _20686_/X _20694_/X _20684_/X vssd1 vssd1 vccd1 vccd1 _25751_/D
+ sky130_fd_sc_hd__o211a_1
X_23483_ _26672_/Q _23101_/X _23491_/S vssd1 vssd1 vccd1 vccd1 _23484_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_13_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_13_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_167_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25222_ _27218_/Q _25217_/X _25220_/X _25221_/X vssd1 vssd1 vccd1 vccd1 _27218_/D
+ sky130_fd_sc_hd__o211a_1
X_22434_ _26246_/Q _22444_/B vssd1 vssd1 vccd1 vccd1 _22434_/X sky130_fd_sc_hd__or2_1
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25153_ _20420_/B _24639_/A _25139_/X _16575_/A _12781_/X vssd1 vssd1 vccd1 vccd1
+ _25153_/X sky130_fd_sc_hd__a221o_1
X_22365_ _22368_/A _22365_/B vssd1 vssd1 vccd1 vccd1 _22366_/A sky130_fd_sc_hd__and2_1
X_24104_ _24104_/A vssd1 vssd1 vccd1 vccd1 _26919_/D sky130_fd_sc_hd__clkbuf_1
X_21316_ input98/X input73/X _21327_/S vssd1 vssd1 vccd1 vccd1 _21316_/X sky130_fd_sc_hd__mux2_8
X_22296_ _26211_/Q _22284_/X _22295_/X _22288_/X vssd1 vssd1 vccd1 vccd1 _26211_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25084_ _27181_/Q _25058_/X _25083_/X vssd1 vssd1 vccd1 vccd1 _27181_/D sky130_fd_sc_hd__o21ba_1
XFILLER_2_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24035_ _26889_/Q _23552_/X _24037_/S vssd1 vssd1 vccd1 vccd1 _24036_/A sky130_fd_sc_hd__mux2_1
X_21247_ _21247_/A vssd1 vssd1 vccd1 vccd1 _21507_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21178_ _25930_/Q _21166_/X _21167_/X input30/X vssd1 vssd1 vccd1 vccd1 _21179_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_132_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20129_ _19763_/X _20113_/X _20128_/Y _20067_/A vssd1 vssd1 vccd1 vccd1 _20129_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_89_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25986_ _25992_/CLK _25986_/D vssd1 vssd1 vccd1 vccd1 _25986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _14610_/A vssd1 vssd1 vccd1 vccd1 _12951_/X sky130_fd_sc_hd__clkbuf_2
X_24937_ _19957_/A _24930_/X _24936_/Y _24921_/X vssd1 vssd1 vccd1 vccd1 _27144_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15670_ _15670_/A vssd1 vssd1 vccd1 vccd1 _15672_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _25474_/Q _25472_/Q _12822_/A vssd1 vssd1 vccd1 vccd1 _12947_/B sky130_fd_sc_hd__o21ba_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24868_ _24866_/Y _24867_/X _24854_/X vssd1 vssd1 vccd1 vccd1 _27123_/D sky130_fd_sc_hd__a21oi_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14621_/A vssd1 vssd1 vccd1 vccd1 _14622_/A sky130_fd_sc_hd__buf_2
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26607_ _26796_/CLK _26607_/D vssd1 vssd1 vccd1 vccd1 _26607_/Q sky130_fd_sc_hd__dfxtp_1
X_23819_ _23728_/X _26793_/Q _23821_/S vssd1 vssd1 vccd1 vccd1 _23820_/A sky130_fd_sc_hd__mux2_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24799_ _20635_/A _24789_/X _24659_/Y _24791_/X vssd1 vssd1 vccd1 vccd1 _24799_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _17336_/X _17341_/C _25533_/Q vssd1 vssd1 vccd1 vccd1 _17342_/B sky130_fd_sc_hd__a21oi_1
XFILLER_199_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14550_/X _14551_/X _14552_/S vssd1 vssd1 vccd1 vccd1 _14552_/X sky130_fd_sc_hd__mux2_1
X_26538_ _26823_/CLK _26538_/D vssd1 vssd1 vccd1 vccd1 _26538_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13503_ _26530_/Q _26138_/Q _13792_/S vssd1 vssd1 vccd1 vccd1 _13503_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _17268_/X _17273_/C _17270_/Y vssd1 vssd1 vccd1 vccd1 _25511_/D sky130_fd_sc_hd__o21a_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26469_ _26601_/CLK _26469_/D vssd1 vssd1 vccd1 vccd1 _26469_/Q sky130_fd_sc_hd__dfxtp_2
X_14483_ _15948_/B _18059_/B _14563_/A vssd1 vssd1 vccd1 vccd1 _16586_/B sky130_fd_sc_hd__a21o_2
XFILLER_202_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19010_ _16624_/B _18978_/B _17838_/X vssd1 vssd1 vccd1 vccd1 _19011_/B sky130_fd_sc_hd__a21bo_1
XFILLER_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16222_ _26803_/Q _26447_/Q _16223_/S vssd1 vssd1 vccd1 vccd1 _16222_/X sky130_fd_sc_hd__mux2_1
X_13434_ _15473_/S _13430_/X _13432_/X _13433_/X vssd1 vssd1 vccd1 vccd1 _13434_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_201_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16153_ _15044_/A _16151_/X _16152_/X vssd1 vssd1 vccd1 vccd1 _16153_/X sky130_fd_sc_hd__o21a_1
X_13365_ _13365_/A vssd1 vssd1 vccd1 vccd1 _13366_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_166_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_wb_clk_i clkbuf_4_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27310_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_182_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15104_ _15841_/S vssd1 vssd1 vccd1 vccd1 _16182_/S sky130_fd_sc_hd__buf_2
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16084_ _16170_/A _16908_/A vssd1 vssd1 vccd1 vccd1 _16084_/Y sky130_fd_sc_hd__nor2_4
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13296_ _13951_/S vssd1 vssd1 vccd1 vccd1 _15768_/S sky130_fd_sc_hd__clkbuf_4
X_19912_ _19912_/A _20227_/B vssd1 vssd1 vccd1 vccd1 _19912_/Y sky130_fd_sc_hd__nor2_1
X_15035_ _15276_/S vssd1 vssd1 vccd1 vccd1 _16225_/S sky130_fd_sc_hd__buf_4
XFILLER_142_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19843_ _19748_/X _19842_/X _19755_/X vssd1 vssd1 vccd1 vccd1 _19843_/X sky130_fd_sc_hd__a21o_1
XFILLER_268_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19774_ _19774_/A _19774_/B vssd1 vssd1 vccd1 vccd1 _19805_/B sky130_fd_sc_hd__and2_1
XFILLER_209_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16986_ _16986_/A _16986_/B vssd1 vssd1 vccd1 vccd1 _16987_/A sky130_fd_sc_hd__and2_1
XFILLER_256_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18725_ _18726_/A _18725_/B vssd1 vssd1 vccd1 vccd1 _19579_/A sky130_fd_sc_hd__xnor2_1
XTAP_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15937_ _26077_/Q _25882_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15937_/X sky130_fd_sc_hd__mux2_1
XTAP_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18656_ _27143_/Q vssd1 vssd1 vccd1 vccd1 _19930_/A sky130_fd_sc_hd__clkbuf_4
X_15868_ _25738_/Q _15868_/B vssd1 vssd1 vccd1 vccd1 _15868_/Y sky130_fd_sc_hd__nor2_1
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17607_ _17615_/A _17607_/B vssd1 vssd1 vccd1 vccd1 _25583_/D sky130_fd_sc_hd__nor2_1
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14819_ _14804_/X _14812_/X _14815_/X _14818_/X vssd1 vssd1 vccd1 vccd1 _14819_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_252_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15799_ _15473_/S _15796_/X _15798_/X _13433_/X vssd1 vssd1 vccd1 vccd1 _15799_/X
+ sky130_fd_sc_hd__a211o_1
X_18587_ _18587_/A vssd1 vssd1 vccd1 vccd1 _25606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_280_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17538_ _25568_/Q _17529_/X _17516_/X _17537_/Y vssd1 vssd1 vccd1 vccd1 _17539_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_189_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17469_ _26251_/Q _17453_/A _17459_/A _25979_/Q vssd1 vssd1 vccd1 vccd1 _17706_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_20_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19208_ _20280_/A _19472_/B vssd1 vssd1 vccd1 vccd1 _19208_/Y sky130_fd_sc_hd__nor2_1
X_20480_ _27164_/Q _20480_/B vssd1 vssd1 vccd1 vccd1 _20480_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_177_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19139_ _18555_/X _19129_/X _19138_/X vssd1 vssd1 vccd1 vccd1 _19139_/X sky130_fd_sc_hd__a21o_4
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22150_ _26168_/Q _22113_/X _22140_/X input262/X _22137_/X vssd1 vssd1 vccd1 vccd1
+ _22150_/X sky130_fd_sc_hd__a221o_1
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput410 _25936_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[0] sky130_fd_sc_hd__buf_2
Xoutput421 _25937_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[1] sky130_fd_sc_hd__buf_2
XFILLER_161_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21101_ _21101_/A vssd1 vssd1 vccd1 vccd1 _25908_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput432 _25938_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[2] sky130_fd_sc_hd__buf_2
XFILLER_218_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput443 _12781_/X vssd1 vssd1 vccd1 vccd1 probe_env[0] sky130_fd_sc_hd__buf_2
X_22081_ _22081_/A vssd1 vssd1 vccd1 vccd1 _26148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput454 _25737_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[13] sky130_fd_sc_hd__buf_2
Xoutput465 _25747_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[23] sky130_fd_sc_hd__buf_2
XFILLER_259_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21032_ _21032_/A vssd1 vssd1 vccd1 vccd1 _25885_/D sky130_fd_sc_hd__clkbuf_1
Xoutput476 _25728_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[4] sky130_fd_sc_hd__buf_2
Xoutput487 _17059_/X vssd1 vssd1 vccd1 vccd1 wmask0[3] sky130_fd_sc_hd__buf_2
XFILLER_114_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25840_ _26467_/CLK _25840_/D vssd1 vssd1 vccd1 vccd1 _25840_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_41_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25771_ _27307_/CLK _25771_/D vssd1 vssd1 vccd1 vccd1 _25771_/Q sky130_fd_sc_hd__dfxtp_4
X_22983_ _22983_/A vssd1 vssd1 vccd1 vccd1 _26464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24722_ _24722_/A _24722_/B vssd1 vssd1 vccd1 vccd1 _27087_/D sky130_fd_sc_hd__nor2_1
XFILLER_228_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21934_ _21934_/A vssd1 vssd1 vccd1 vccd1 _26083_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24653_ _17444_/C _12778_/B _19640_/A _24635_/A _24771_/A vssd1 vssd1 vccd1 vccd1
+ _24654_/B sky130_fd_sc_hd__o311a_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21865_ _21865_/A vssd1 vssd1 vccd1 vccd1 _26060_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_256_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23604_ _26713_/Q _23603_/X _23604_/S vssd1 vssd1 vccd1 vccd1 _23605_/A sky130_fd_sc_hd__mux2_1
X_20816_ _25804_/Q vssd1 vssd1 vccd1 vccd1 _20817_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_169_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24584_ _24610_/A vssd1 vssd1 vccd1 vccd1 _24595_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21796_ _21864_/S vssd1 vssd1 vccd1 vccd1 _21805_/S sky130_fd_sc_hd__buf_2
XFILLER_24_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26323_ _26327_/CLK _26323_/D vssd1 vssd1 vccd1 vccd1 _26323_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_195_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23535_ _23535_/A vssd1 vssd1 vccd1 vccd1 _26691_/D sky130_fd_sc_hd__clkbuf_1
X_20747_ _20747_/A vssd1 vssd1 vccd1 vccd1 _25770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26254_ _26257_/CLK _26254_/D vssd1 vssd1 vccd1 vccd1 _26254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23466_ _23466_/A vssd1 vssd1 vccd1 vccd1 _26664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20678_ _26281_/Q _20673_/X _20677_/X _20671_/X vssd1 vssd1 vccd1 vccd1 _25744_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25205_ _24707_/B _25198_/X _25204_/X _27214_/Q _25199_/X vssd1 vssd1 vccd1 vccd1
+ _27214_/D sky130_fd_sc_hd__o221a_1
X_22417_ _22638_/A _26219_/Q _22554_/A _22419_/D vssd1 vssd1 vccd1 vccd1 _22459_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26185_ _26186_/CLK _26185_/D vssd1 vssd1 vccd1 vccd1 _26185_/Q sky130_fd_sc_hd__dfxtp_1
X_23397_ _26634_/Q _23082_/X _23397_/S vssd1 vssd1 vccd1 vccd1 _23398_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13150_ _15796_/S vssd1 vssd1 vccd1 vccd1 _15555_/S sky130_fd_sc_hd__buf_4
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25136_ _27191_/Q _25112_/X _25135_/X vssd1 vssd1 vccd1 vccd1 _27191_/D sky130_fd_sc_hd__o21ba_1
X_22348_ _22428_/A vssd1 vssd1 vccd1 vccd1 _22348_/X sky130_fd_sc_hd__buf_2
XFILLER_3_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13081_ _15559_/S vssd1 vssd1 vccd1 vccd1 _15645_/S sky130_fd_sc_hd__buf_2
XFILLER_151_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25067_ _20652_/A _25059_/X _25066_/X vssd1 vssd1 vccd1 vccd1 _25067_/Y sky130_fd_sc_hd__o21ai_1
X_22279_ _22310_/A vssd1 vssd1 vccd1 vccd1 _22279_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24018_ _26881_/Q _23526_/X _24026_/S vssd1 vssd1 vccd1 vccd1 _24019_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ _16840_/A vssd1 vssd1 vccd1 vccd1 _16840_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16771_ _22520_/A _16769_/X _16770_/X _16606_/Y vssd1 vssd1 vccd1 vccd1 _16771_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_120_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13983_ _26658_/Q _15797_/B vssd1 vssd1 vccd1 vccd1 _13983_/X sky130_fd_sc_hd__or2_1
X_25969_ _27156_/CLK _25969_/D vssd1 vssd1 vccd1 vccd1 _25969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15722_ _26667_/Q _15800_/S _15721_/X _13050_/A vssd1 vssd1 vccd1 vccd1 _15722_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18510_ _18510_/A vssd1 vssd1 vccd1 vccd1 _18510_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_207_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12934_ _12934_/A vssd1 vssd1 vccd1 vccd1 _14031_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ _19484_/X _17764_/X _19487_/X _19489_/X vssd1 vssd1 vccd1 vccd1 _25630_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_207_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18441_ _18441_/A vssd1 vssd1 vccd1 vccd1 _18441_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15653_ _26112_/Q _26013_/Q _15653_/S vssd1 vssd1 vccd1 vccd1 _15653_/X sky130_fd_sc_hd__mux2_1
X_12865_ _12862_/A _15706_/A _15708_/A _12942_/A _12866_/B vssd1 vssd1 vccd1 vccd1
+ _12865_/X sky130_fd_sc_hd__o221a_1
XFILLER_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14604_ _14604_/A _14604_/B vssd1 vssd1 vccd1 vccd1 _16292_/B sky130_fd_sc_hd__or2_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _18368_/X _18371_/X _18372_/S vssd1 vssd1 vccd1 vccd1 _18372_/X sky130_fd_sc_hd__mux2_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _15843_/A vssd1 vssd1 vccd1 vccd1 _15670_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _25597_/Q vssd1 vssd1 vccd1 vccd1 _12992_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _17332_/A _17323_/B _17324_/B vssd1 vssd1 vccd1 vccd1 _25527_/D sky130_fd_sc_hd__nor3_1
XFILLER_199_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _14535_/A _14535_/B _14535_/C vssd1 vssd1 vccd1 vccd1 _14535_/X sky130_fd_sc_hd__or3_1
XFILLER_186_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17254_ _17285_/A _17256_/B vssd1 vssd1 vccd1 vccd1 _17254_/Y sky130_fd_sc_hd__nor2_1
X_14466_ _13344_/A _14464_/X _14465_/X _13939_/A vssd1 vssd1 vccd1 vccd1 _14466_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16205_ _17791_/A _16206_/B vssd1 vssd1 vccd1 vccd1 _16207_/A sky130_fd_sc_hd__nor2_2
X_13417_ _27241_/Q _15468_/B vssd1 vssd1 vccd1 vccd1 _13417_/X sky130_fd_sc_hd__or2_1
XFILLER_139_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17185_ _25489_/Q _17185_/B vssd1 vssd1 vccd1 vccd1 _17185_/X sky130_fd_sc_hd__or2_1
XFILLER_128_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14397_ _13465_/A _23517_/A _14396_/X _13683_/A vssd1 vssd1 vccd1 vccd1 _19665_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_155_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16136_ _15167_/X _26413_/Q _15142_/A _16135_/X vssd1 vssd1 vccd1 vccd1 _16136_/X
+ sky130_fd_sc_hd__o211a_1
X_13348_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13835_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_255_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16067_ _25848_/Q _26048_/Q _16067_/S vssd1 vssd1 vccd1 vccd1 _16067_/X sky130_fd_sc_hd__mux2_1
X_13279_ _15859_/A vssd1 vssd1 vccd1 vccd1 _15576_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_142_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15018_ _12775_/A _26418_/Q _15060_/S _15017_/X vssd1 vssd1 vccd1 vccd1 _15018_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19826_ _25731_/Q vssd1 vssd1 vccd1 vccd1 _20641_/A sky130_fd_sc_hd__buf_8
XFILLER_68_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19757_ _22515_/A vssd1 vssd1 vccd1 vccd1 _22480_/B sky130_fd_sc_hd__clkbuf_2
X_16969_ _16868_/X _16954_/X _16956_/X _16867_/X _16968_/X vssd1 vssd1 vccd1 vccd1
+ _16970_/C sky130_fd_sc_hd__a221o_1
XFILLER_244_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18708_ _19946_/A _18843_/D vssd1 vssd1 vccd1 vccd1 _18781_/B sky130_fd_sc_hd__nand2_2
X_19688_ _27134_/Q _25173_/A _27133_/Q vssd1 vssd1 vccd1 vccd1 _20000_/A sky130_fd_sc_hd__or3b_4
XFILLER_253_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18639_ _18684_/S _18199_/X _17966_/A vssd1 vssd1 vccd1 vccd1 _18639_/X sky130_fd_sc_hd__a21o_1
XFILLER_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21650_ _25967_/Q _21273_/A _21649_/Y _17283_/A vssd1 vssd1 vccd1 vccd1 _25967_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_80_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20601_ _23770_/A vssd1 vssd1 vccd1 vccd1 _20601_/X sky130_fd_sc_hd__clkbuf_2
X_21581_ _21581_/A vssd1 vssd1 vccd1 vccd1 _21581_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23320_ _20542_/X _26600_/Q _23324_/S vssd1 vssd1 vccd1 vccd1 _23321_/A sky130_fd_sc_hd__mux2_1
X_20532_ _23542_/A vssd1 vssd1 vccd1 vccd1 _23718_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_193_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23251_ _26569_/Q _23092_/X _23255_/S vssd1 vssd1 vccd1 vccd1 _23252_/A sky130_fd_sc_hd__mux2_1
X_20463_ _22533_/A _20003_/X _20454_/X _20462_/X _20346_/X vssd1 vssd1 vccd1 vccd1
+ _25690_/D sky130_fd_sc_hd__o221a_1
XFILLER_192_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22202_ input2/X input268/X _22207_/S vssd1 vssd1 vccd1 vccd1 _22202_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23182_ _23182_/A vssd1 vssd1 vccd1 vccd1 _26538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20394_ _22528_/A _20003_/X _20386_/X _20393_/X _20346_/X vssd1 vssd1 vccd1 vccd1
+ _25687_/D sky130_fd_sc_hd__o221a_1
XFILLER_106_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22133_ _26163_/Q _22110_/X _22129_/X _22132_/X vssd1 vssd1 vccd1 vccd1 _26163_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_161_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26941_ _26974_/CLK _26941_/D vssd1 vssd1 vccd1 vccd1 _26941_/Q sky130_fd_sc_hd__dfxtp_1
X_22064_ _26141_/Q _20913_/X _22066_/S vssd1 vssd1 vccd1 vccd1 _22065_/A sky130_fd_sc_hd__mux2_1
Xoutput295 _16992_/X vssd1 vssd1 vccd1 vccd1 addr1[1] sky130_fd_sc_hd__buf_2
XFILLER_275_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_2 _19896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21015_ _25878_/Q _20900_/X _21015_/S vssd1 vssd1 vccd1 vccd1 _21016_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26872_ _27259_/CLK _26872_/D vssd1 vssd1 vccd1 vccd1 _26872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25823_ _26744_/CLK _25823_/D vssd1 vssd1 vccd1 vccd1 _25823_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25754_ _26292_/CLK _25754_/D vssd1 vssd1 vccd1 vccd1 _25754_/Q sky130_fd_sc_hd__dfxtp_4
X_22966_ _22966_/A vssd1 vssd1 vccd1 vccd1 _26456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24705_ _24722_/A _24705_/B vssd1 vssd1 vccd1 vccd1 _27083_/D sky130_fd_sc_hd__nor2_1
X_21917_ _21917_/A vssd1 vssd1 vccd1 vccd1 _26075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25685_ _25690_/CLK _25685_/D vssd1 vssd1 vccd1 vccd1 _25685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22897_ _26426_/Q _22650_/X _22901_/S vssd1 vssd1 vccd1 vccd1 _22898_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24636_ _24636_/A vssd1 vssd1 vccd1 vccd1 _24636_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_169_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21848_ _21848_/A vssd1 vssd1 vccd1 vccd1 _26052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24567_ _24619_/A vssd1 vssd1 vccd1 vccd1 _24567_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21779_ _20596_/X _26022_/Q _21787_/S vssd1 vssd1 vccd1 vccd1 _21780_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26306_ _26307_/CLK _26306_/D vssd1 vssd1 vccd1 vccd1 _26306_/Q sky130_fd_sc_hd__dfxtp_2
X_14320_ input129/X input134/X _14320_/S vssd1 vssd1 vccd1 vccd1 _14321_/B sky130_fd_sc_hd__mux2_8
XFILLER_157_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23518_ _26686_/Q _23517_/X _23524_/S vssd1 vssd1 vccd1 vccd1 _23519_/A sky130_fd_sc_hd__mux2_1
X_27286_ _27287_/CLK _27286_/D vssd1 vssd1 vccd1 vccd1 _27286_/Q sky130_fd_sc_hd__dfxtp_1
X_24498_ _24518_/A _24611_/A vssd1 vssd1 vccd1 vccd1 _24498_/Y sky130_fd_sc_hd__nand2_1
X_26237_ _26238_/CLK _26237_/D vssd1 vssd1 vccd1 vccd1 _26237_/Q sky130_fd_sc_hd__dfxtp_1
X_14251_ _13863_/X _14246_/X _14250_/X _13112_/A vssd1 vssd1 vccd1 vccd1 _14251_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23449_ _23506_/S vssd1 vssd1 vccd1 vccd1 _23458_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_172_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13202_ _23363_/B _13365_/A _13336_/A _21793_/A _13201_/X vssd1 vssd1 vccd1 vccd1
+ _13202_/X sky130_fd_sc_hd__a221o_1
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26168_ _27264_/CLK _26168_/D vssd1 vssd1 vccd1 vccd1 _26168_/Q sky130_fd_sc_hd__dfxtp_1
X_14182_ _13141_/A _14178_/X _14181_/X _14522_/S vssd1 vssd1 vccd1 vccd1 _14182_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13133_ _14330_/A vssd1 vssd1 vccd1 vccd1 _13134_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_174_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25119_ _25119_/A vssd1 vssd1 vccd1 vccd1 _25119_/X sky130_fd_sc_hd__clkbuf_2
X_26099_ _26592_/CLK _26099_/D vssd1 vssd1 vccd1 vccd1 _26099_/Q sky130_fd_sc_hd__dfxtp_1
X_18990_ _27022_/Q _18756_/X _18989_/X _18759_/X vssd1 vssd1 vccd1 vccd1 _18990_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _14246_/S vssd1 vssd1 vccd1 vccd1 _13065_/A sky130_fd_sc_hd__buf_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _17941_/A vssd1 vssd1 vccd1 vccd1 _18202_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_78_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17872_ _18058_/S vssd1 vssd1 vccd1 vccd1 _18070_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_238_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19611_ _27065_/Q _19616_/B _19611_/C vssd1 vssd1 vccd1 vccd1 _19614_/B sky130_fd_sc_hd__and3_1
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16823_ _16838_/A _16823_/B vssd1 vssd1 vccd1 vccd1 _16868_/B sky130_fd_sc_hd__nor2_4
XFILLER_226_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19542_ _19538_/X _19099_/X _19540_/X _19541_/X vssd1 vssd1 vccd1 vccd1 _25650_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13966_ _13966_/A vssd1 vssd1 vccd1 vccd1 _15516_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_207_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16754_ _22507_/A _16742_/X _16743_/X _16637_/C vssd1 vssd1 vccd1 vccd1 _16754_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15705_ _12912_/A _15704_/Y _12929_/A vssd1 vssd1 vccd1 vccd1 _15705_/X sky130_fd_sc_hd__a21o_1
X_12917_ _13389_/A vssd1 vssd1 vccd1 vccd1 _14133_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16685_ _22530_/A _16685_/B vssd1 vssd1 vccd1 vccd1 _21190_/A sky130_fd_sc_hd__nor2_4
X_19473_ _17673_/X _19471_/X _19472_/Y vssd1 vssd1 vccd1 vccd1 _19473_/Y sky130_fd_sc_hd__a21oi_1
X_13897_ _26103_/Q _26004_/Q _14245_/S vssd1 vssd1 vccd1 vccd1 _13897_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18424_ _18424_/A _19289_/B vssd1 vssd1 vccd1 vccd1 _18424_/X sky130_fd_sc_hd__or2_1
X_12848_ _12872_/A _14131_/A vssd1 vssd1 vccd1 vccd1 _12869_/A sky130_fd_sc_hd__nor2_1
X_15636_ _26080_/Q _15623_/B _15546_/S _15635_/X vssd1 vssd1 vccd1 vccd1 _15636_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15567_ _15565_/X _15566_/X _15567_/S vssd1 vssd1 vccd1 vccd1 _15567_/X sky130_fd_sc_hd__mux2_1
X_18355_ _16717_/A _18328_/A _17802_/A _18354_/Y vssd1 vssd1 vccd1 vccd1 _19572_/A
+ sky130_fd_sc_hd__a211oi_2
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _25113_/A vssd1 vssd1 vccd1 vccd1 _25106_/A sky130_fd_sc_hd__inv_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17306_ _17334_/A _17312_/C vssd1 vssd1 vccd1 vccd1 _17306_/Y sky130_fd_sc_hd__nor2_1
X_14518_ _26620_/Q _26716_/Q _14518_/S vssd1 vssd1 vccd1 vccd1 _14518_/X sky130_fd_sc_hd__mux2_1
X_15498_ _15509_/A _15498_/B vssd1 vssd1 vccd1 vccd1 _15498_/X sky130_fd_sc_hd__or2_1
XFILLER_30_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18286_ _25728_/Q _18287_/B vssd1 vssd1 vccd1 vccd1 _18432_/C sky130_fd_sc_hd__and2_1
XFILLER_266_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14449_ _25870_/Q _14449_/B vssd1 vssd1 vccd1 vccd1 _14449_/X sky130_fd_sc_hd__or2_1
X_17237_ _17242_/A _17242_/B _17236_/Y vssd1 vssd1 vccd1 vccd1 _25502_/D sky130_fd_sc_hd__o21a_1
XFILLER_134_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17168_ _19392_/A _17195_/B vssd1 vssd1 vccd1 vccd1 _17168_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16119_ _16093_/Y _16101_/Y _16118_/Y _13314_/X _13466_/X vssd1 vssd1 vccd1 vccd1
+ _16119_/Y sky130_fd_sc_hd__o221ai_4
X_17099_ _22340_/S _26229_/Q _17078_/X _17098_/X vssd1 vssd1 vccd1 vccd1 _17099_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_171_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_257_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19809_ _19809_/A _19830_/B vssd1 vssd1 vccd1 vccd1 _19809_/Y sky130_fd_sc_hd__nand2_1
XFILLER_229_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22820_ _22888_/S vssd1 vssd1 vccd1 vccd1 _22829_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_226_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22751_ _22751_/A vssd1 vssd1 vccd1 vccd1 _26361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21702_ _21702_/A vssd1 vssd1 vccd1 vccd1 _25989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25470_ _25598_/CLK _25470_/D vssd1 vssd1 vccd1 vccd1 _25470_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_53_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22682_ _23725_/A vssd1 vssd1 vccd1 vccd1 _22682_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_212_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24421_ _24506_/A vssd1 vssd1 vccd1 vccd1 _24421_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21633_ _25754_/Q _21278_/A _21563_/A _21632_/X vssd1 vssd1 vccd1 vccd1 _21633_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_240_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27140_ _27166_/CLK _27140_/D vssd1 vssd1 vccd1 vccd1 _27140_/Q sky130_fd_sc_hd__dfxtp_1
X_24352_ _17483_/Y _17684_/B _24351_/Y _24340_/S vssd1 vssd1 vccd1 vccd1 _24352_/X
+ sky130_fd_sc_hd__o22a_1
X_21564_ _19246_/A _21545_/X _21561_/X _21563_/X vssd1 vssd1 vccd1 vccd1 _21564_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23303_ _23303_/A vssd1 vssd1 vccd1 vccd1 _26592_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20515_ _20515_/A vssd1 vssd1 vccd1 vccd1 _25697_/D sky130_fd_sc_hd__clkbuf_1
X_27071_ _27203_/CLK _27071_/D vssd1 vssd1 vccd1 vccd1 _27071_/Q sky130_fd_sc_hd__dfxtp_1
X_24283_ _26984_/Q _24284_/C _26985_/Q vssd1 vssd1 vccd1 vccd1 _24285_/B sky130_fd_sc_hd__a21oi_1
XFILLER_197_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21495_ _25487_/Q _21495_/B vssd1 vssd1 vccd1 vccd1 _21495_/X sky130_fd_sc_hd__or2_1
XFILLER_181_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26022_ _27259_/CLK _26022_/D vssd1 vssd1 vccd1 vccd1 _26022_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_179_wb_clk_i clkbuf_4_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26715_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23234_ _23234_/A vssd1 vssd1 vccd1 vccd1 _26561_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20446_ _25754_/Q _20355_/X _20445_/Y _20357_/X vssd1 vssd1 vccd1 vccd1 _20448_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_109_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_108_wb_clk_i clkbuf_4_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26257_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_134_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_279_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23165_ _23165_/A vssd1 vssd1 vccd1 vccd1 _26530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20377_ _19341_/A _18019_/X _19348_/X _20376_/Y vssd1 vssd1 vccd1 vccd1 _20377_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22116_ _22121_/A _22239_/B vssd1 vssd1 vccd1 vccd1 _22203_/A sky130_fd_sc_hd__or2_1
XFILLER_133_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23096_ _26506_/Q _23095_/X _23099_/S vssd1 vssd1 vccd1 vccd1 _23097_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22047_ _26133_/Q _20887_/X _22055_/S vssd1 vssd1 vccd1 vccd1 _22048_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26924_ _27311_/CLK _26924_/D vssd1 vssd1 vccd1 vccd1 _26924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26855_ _27306_/CLK _26855_/D vssd1 vssd1 vccd1 vccd1 _26855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_275_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13820_ _26627_/Q _26723_/Q _13951_/S vssd1 vssd1 vccd1 vccd1 _13821_/B sky130_fd_sc_hd__mux2_1
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25806_ _27295_/CLK _25806_/D vssd1 vssd1 vccd1 vccd1 _25806_/Q sky130_fd_sc_hd__dfxtp_4
X_26786_ _27238_/CLK _26786_/D vssd1 vssd1 vccd1 vccd1 _26786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23998_ _26873_/Q _23603_/X _23998_/S vssd1 vssd1 vccd1 vccd1 _23999_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13751_ _25638_/Q _16130_/B _13578_/X _25606_/Q vssd1 vssd1 vccd1 vccd1 _13751_/X
+ sky130_fd_sc_hd__a22o_1
X_25737_ _25737_/CLK _25737_/D vssd1 vssd1 vccd1 vccd1 _25737_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_109 _21878_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22949_ _22949_/A vssd1 vssd1 vccd1 vccd1 _26449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12702_ _12702_/A vssd1 vssd1 vccd1 vccd1 _12703_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_216_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16470_ _16498_/S vssd1 vssd1 vccd1 vccd1 _16490_/B sky130_fd_sc_hd__clkbuf_2
X_13682_ _14820_/A _13662_/X _13671_/X _13681_/X _14722_/A vssd1 vssd1 vccd1 vccd1
+ _13682_/X sky130_fd_sc_hd__a221o_4
X_25668_ _25670_/CLK _25668_/D vssd1 vssd1 vccd1 vccd1 _25668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15421_ _15227_/S _15419_/X _15420_/X _16185_/A vssd1 vssd1 vccd1 vccd1 _15421_/X
+ sky130_fd_sc_hd__a31o_1
XPHY_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24619_ _24619_/A vssd1 vssd1 vccd1 vccd1 _24619_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25599_ _25599_/CLK _25599_/D vssd1 vssd1 vccd1 vccd1 _25599_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15352_ _15167_/X _26412_/Q _15142_/A _15351_/X vssd1 vssd1 vccd1 vccd1 _15352_/X
+ sky130_fd_sc_hd__o211a_1
X_18140_ _18910_/A _18135_/X _18705_/A vssd1 vssd1 vccd1 vccd1 _18140_/X sky130_fd_sc_hd__o21ba_1
XFILLER_157_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14303_ _25800_/Q _27234_/Q _14310_/S vssd1 vssd1 vccd1 vccd1 _14303_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18071_ _18069_/X _18070_/X _18071_/S vssd1 vssd1 vccd1 vccd1 _18071_/X sky130_fd_sc_hd__mux2_1
X_27269_ _27269_/CLK _27269_/D vssd1 vssd1 vccd1 vccd1 _27269_/Q sky130_fd_sc_hd__dfxtp_1
X_15283_ _15065_/A _26706_/Q _26834_/Q _16134_/S _15169_/X vssd1 vssd1 vccd1 vccd1
+ _15283_/X sky130_fd_sc_hd__a221o_1
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17022_ _17021_/X _16857_/B _17017_/X input216/X vssd1 vssd1 vccd1 vccd1 _17022_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_8_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14234_ _17800_/C vssd1 vssd1 vccd1 vccd1 _14570_/B sky130_fd_sc_hd__buf_2
XFILLER_138_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14165_ _14165_/A _14165_/B vssd1 vssd1 vccd1 vccd1 _14165_/Y sky130_fd_sc_hd__nand2_1
XFILLER_259_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13116_ _15566_/S vssd1 vssd1 vccd1 vccd1 _15540_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_98_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14096_ _26625_/Q _26721_/Q _14265_/S vssd1 vssd1 vccd1 vccd1 _14096_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18973_ _18973_/A vssd1 vssd1 vccd1 vccd1 _18973_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13047_ _13610_/A vssd1 vssd1 vccd1 vccd1 _13048_/A sky130_fd_sc_hd__buf_2
X_17924_ _14567_/A _17851_/B _17949_/S vssd1 vssd1 vccd1 vccd1 _17924_/X sky130_fd_sc_hd__mux2_1
XFILLER_252_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17855_ _19452_/A _19452_/B _17857_/A vssd1 vssd1 vccd1 vccd1 _19585_/S sky130_fd_sc_hd__a21oi_1
XFILLER_78_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16806_ _16887_/A vssd1 vssd1 vccd1 vccd1 _16812_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17786_ _17786_/A vssd1 vssd1 vccd1 vccd1 _17787_/B sky130_fd_sc_hd__inv_2
XFILLER_282_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14998_ _25825_/Q _27259_/Q _15005_/S vssd1 vssd1 vccd1 vccd1 _14998_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19525_ _19551_/A vssd1 vssd1 vccd1 vccd1 _19525_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16737_ _25671_/Q vssd1 vssd1 vccd1 vccd1 _22494_/A sky130_fd_sc_hd__buf_2
X_13949_ _13252_/A _26882_/Q _26754_/Q _15938_/S _13943_/X vssd1 vssd1 vccd1 vccd1
+ _13949_/X sky130_fd_sc_hd__a221o_1
XFILLER_35_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_281_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19456_ _16550_/A _19455_/X _17927_/Y vssd1 vssd1 vccd1 vccd1 _19456_/X sky130_fd_sc_hd__a21o_1
XFILLER_222_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16668_ _20977_/A _16668_/B vssd1 vssd1 vccd1 vccd1 _16669_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_250_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18407_ _18891_/A _19768_/A _19768_/B _18406_/X _18005_/A vssd1 vssd1 vccd1 vccd1
+ _18407_/X sky130_fd_sc_hd__a311o_1
XFILLER_222_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15619_ _25646_/Q _16130_/B vssd1 vssd1 vccd1 vccd1 _15619_/X sky130_fd_sc_hd__and2_1
XFILLER_22_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19387_ _25626_/Q _18719_/A _19386_/X _19352_/X vssd1 vssd1 vccd1 vccd1 _25626_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_250_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16599_ _16603_/B vssd1 vssd1 vccd1 vccd1 _19639_/B sky130_fd_sc_hd__buf_2
XFILLER_194_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18338_ _18338_/A vssd1 vssd1 vccd1 vccd1 _18630_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_6_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27253_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_147_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18269_ _18269_/A _18269_/B vssd1 vssd1 vccd1 vccd1 _18269_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20300_ _20300_/A _20300_/B _20300_/C _20300_/D vssd1 vssd1 vccd1 vccd1 _20302_/A
+ sky130_fd_sc_hd__or4_1
X_21280_ _21507_/A vssd1 vssd1 vccd1 vccd1 _21559_/B sky130_fd_sc_hd__clkbuf_2
X_20231_ _20305_/A _20260_/B _20300_/B vssd1 vssd1 vccd1 vccd1 _20231_/X sky130_fd_sc_hd__or3_1
XFILLER_190_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20162_ _19894_/X _20161_/X _19902_/X vssd1 vssd1 vccd1 vccd1 _20162_/X sky130_fd_sc_hd__a21o_1
XFILLER_277_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24970_ _25221_/A vssd1 vssd1 vccd1 vccd1 _24970_/X sky130_fd_sc_hd__clkbuf_2
X_20093_ _20376_/A _18965_/X _18019_/X _15698_/Y vssd1 vssd1 vccd1 vccd1 _20093_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_58_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23921_ _23921_/A vssd1 vssd1 vccd1 vccd1 _26838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_273_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_257_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26640_ _27315_/CLK _26640_/D vssd1 vssd1 vccd1 vccd1 _26640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23852_ _23776_/X _26808_/Q _23854_/S vssd1 vssd1 vccd1 vccd1 _23853_/A sky130_fd_sc_hd__mux2_1
XFILLER_273_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22803_ _26385_/Q _22723_/X _22811_/S vssd1 vssd1 vccd1 vccd1 _22804_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26571_ _26799_/CLK _26571_/D vssd1 vssd1 vccd1 vccd1 _26571_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23783_ _23782_/X _26778_/Q _23786_/S vssd1 vssd1 vccd1 vccd1 _23784_/A sky130_fd_sc_hd__mux2_1
XFILLER_272_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20995_ _21063_/S vssd1 vssd1 vccd1 vccd1 _21004_/S sky130_fd_sc_hd__buf_2
XFILLER_260_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25522_ _27022_/CLK _25522_/D vssd1 vssd1 vccd1 vccd1 _25522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22734_ _26356_/Q _22733_/X _22737_/S vssd1 vssd1 vccd1 vccd1 _22735_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25453_ _23770_/X _27321_/Q _25459_/S vssd1 vssd1 vccd1 vccd1 _25454_/A sky130_fd_sc_hd__mux2_1
X_22665_ _22665_/A vssd1 vssd1 vccd1 vccd1 _26334_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24404_ _24501_/A vssd1 vssd1 vccd1 vccd1 _24404_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_231_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21616_ _21616_/A vssd1 vssd1 vccd1 vccd1 _21616_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25384_ _25384_/A vssd1 vssd1 vccd1 vccd1 _27290_/D sky130_fd_sc_hd__clkbuf_1
X_22596_ _22593_/X _22595_/Y _22587_/X vssd1 vssd1 vccd1 vccd1 _26313_/D sky130_fd_sc_hd__a21oi_1
X_27123_ _27130_/CLK _27123_/D vssd1 vssd1 vccd1 vccd1 _27123_/Q sky130_fd_sc_hd__dfxtp_4
X_24335_ _24335_/A _24335_/B vssd1 vssd1 vccd1 vccd1 _24335_/Y sky130_fd_sc_hd__nor2_1
XFILLER_166_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21547_ _21547_/A vssd1 vssd1 vccd1 vccd1 _21547_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27054_ _27062_/CLK _27054_/D vssd1 vssd1 vccd1 vccd1 _27054_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_193_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24266_ _26979_/Q _26978_/Q _24266_/C vssd1 vssd1 vccd1 vccd1 _24268_/B sky130_fd_sc_hd__and3_1
XFILLER_153_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21478_ _21474_/Y _21477_/X _21425_/X vssd1 vssd1 vccd1 vccd1 _21478_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_5_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26005_ _27276_/CLK _26005_/D vssd1 vssd1 vccd1 vccd1 _26005_/Q sky130_fd_sc_hd__dfxtp_4
X_23217_ _23217_/A vssd1 vssd1 vccd1 vccd1 _26553_/D sky130_fd_sc_hd__clkbuf_1
X_20429_ _20467_/C _20421_/Y _19941_/X _20428_/X vssd1 vssd1 vccd1 vccd1 _20429_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24197_ _26956_/Q _26955_/Q _24197_/C vssd1 vssd1 vccd1 vccd1 _24203_/C sky130_fd_sc_hd__and3_1
XFILLER_181_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23148_ _26523_/Q _23047_/X _23150_/S vssd1 vssd1 vccd1 vccd1 _23149_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15970_ _15968_/X _15969_/X _15970_/S vssd1 vssd1 vccd1 vccd1 _15970_/X sky130_fd_sc_hd__mux2_1
X_23079_ _23552_/A vssd1 vssd1 vccd1 vccd1 _23079_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14921_ _26093_/Q _25898_/Q _15003_/S vssd1 vssd1 vccd1 vccd1 _14921_/X sky130_fd_sc_hd__mux2_1
X_26907_ _26939_/CLK _26907_/D vssd1 vssd1 vccd1 vccd1 _26907_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_76_wb_clk_i clkbuf_4_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _26909_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_249_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _17444_/A _17635_/X _17604_/X _17639_/Y vssd1 vssd1 vccd1 vccd1 _17641_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_5598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26838_ _27322_/CLK _26838_/D vssd1 vssd1 vccd1 vccd1 _26838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14852_ _14693_/S _14849_/X _14851_/X _14662_/A vssd1 vssd1 vccd1 vccd1 _14852_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_75_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13803_ _25637_/Q _13803_/B vssd1 vssd1 vccd1 vccd1 _13803_/X sky130_fd_sc_hd__and2_1
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14783_ _26550_/Q _26158_/Q _16510_/A vssd1 vssd1 vccd1 vccd1 _14783_/X sky130_fd_sc_hd__mux2_1
X_17571_ _17575_/A _17571_/B vssd1 vssd1 vccd1 vccd1 _25574_/D sky130_fd_sc_hd__nor2_1
XFILLER_44_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26769_ _27316_/CLK _26769_/D vssd1 vssd1 vccd1 vccd1 _26769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19310_ _18741_/X _19308_/X _19309_/Y vssd1 vssd1 vccd1 vccd1 _19310_/Y sky130_fd_sc_hd__a21oi_1
X_13734_ _14677_/A _13722_/X _13726_/X _14681_/A _13733_/X vssd1 vssd1 vccd1 vccd1
+ _13734_/X sky130_fd_sc_hd__a311o_2
X_16522_ _26551_/Q _26159_/Q _16523_/S vssd1 vssd1 vccd1 vccd1 _16522_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19241_ _17782_/A _17781_/A _18733_/X _19240_/X vssd1 vssd1 vccd1 vccd1 _19241_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13665_ _14221_/S vssd1 vssd1 vccd1 vccd1 _15915_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16453_ _16453_/A _17780_/B vssd1 vssd1 vccd1 vccd1 _16454_/B sky130_fd_sc_hd__nor2_1
XFILLER_220_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _15417_/A _15404_/B vssd1 vssd1 vccd1 vccd1 _15404_/X sky130_fd_sc_hd__or2_1
X_19172_ _18806_/X _19162_/X _19171_/X vssd1 vssd1 vccd1 vccd1 _19172_/X sky130_fd_sc_hd__a21o_4
X_16384_ _26355_/Q _26615_/Q _16384_/S vssd1 vssd1 vccd1 vccd1 _16384_/X sky130_fd_sc_hd__mux2_1
X_13596_ _27304_/Q _26561_/Q _15816_/S vssd1 vssd1 vccd1 vccd1 _13596_/X sky130_fd_sc_hd__mux2_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18123_ _27038_/Q _19055_/A _18115_/X _19066_/A vssd1 vssd1 vccd1 vccd1 _18123_/X
+ sky130_fd_sc_hd__o211a_1
X_15335_ _15318_/X _15329_/X _15334_/X _14817_/A vssd1 vssd1 vccd1 vccd1 _15335_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_200_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18054_ _18050_/X _18053_/X _18318_/S vssd1 vssd1 vccd1 vccd1 _18054_/X sky130_fd_sc_hd__mux2_1
X_15266_ _25891_/Q _16154_/B vssd1 vssd1 vccd1 vccd1 _15266_/X sky130_fd_sc_hd__or2_1
XFILLER_117_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14217_ _25801_/Q _27235_/Q _15775_/S vssd1 vssd1 vccd1 vccd1 _14217_/X sky130_fd_sc_hd__mux2_1
X_17005_ _16784_/X _17001_/X _16848_/B _17003_/X input226/X vssd1 vssd1 vccd1 vccd1
+ _17005_/X sky130_fd_sc_hd__a32o_4
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15197_ _15197_/A vssd1 vssd1 vccd1 vccd1 _16259_/S sky130_fd_sc_hd__buf_6
XFILLER_126_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14148_ _26524_/Q _26132_/Q _14265_/S vssd1 vssd1 vccd1 vccd1 _14148_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18956_ _25549_/Q _18568_/A _18955_/X _19069_/A _18572_/A vssd1 vssd1 vccd1 vccd1
+ _18956_/X sky130_fd_sc_hd__a221o_1
X_14079_ _13465_/A _23526_/A _14078_/X _13683_/A vssd1 vssd1 vccd1 vccd1 _19769_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_67_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17907_ _17818_/B _16287_/B _17954_/S vssd1 vssd1 vccd1 vccd1 _17907_/X sky130_fd_sc_hd__mux2_1
XFILLER_273_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18887_ _19042_/A _18887_/B vssd1 vssd1 vccd1 vccd1 _18887_/Y sky130_fd_sc_hd__nand2_1
X_17838_ _17838_/A _16043_/B vssd1 vssd1 vccd1 vccd1 _17838_/X sky130_fd_sc_hd__or2b_1
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17769_ _17769_/A _18076_/B vssd1 vssd1 vccd1 vccd1 _18945_/A sky130_fd_sc_hd__nand2_1
XFILLER_270_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19508_ _25638_/Q _19510_/B vssd1 vssd1 vccd1 vccd1 _19508_/X sky130_fd_sc_hd__or2_1
XFILLER_207_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20780_ _20780_/A vssd1 vssd1 vccd1 vccd1 _25785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_440 _25730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_451 _17057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19439_ _25563_/Q _18763_/X _19438_/X _18767_/X _18768_/X vssd1 vssd1 vccd1 vccd1
+ _19439_/X sky130_fd_sc_hd__a221o_1
XFILLER_179_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_462 _19000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_473 _17712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_484 _21195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_495 _16681_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22450_ _26252_/Q _22457_/B vssd1 vssd1 vccd1 vccd1 _22450_/X sky130_fd_sc_hd__or2_1
XFILLER_195_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21401_ _25947_/Q _21378_/X _21398_/Y _21400_/X vssd1 vssd1 vccd1 vccd1 _25947_/D
+ sky130_fd_sc_hd__a211o_1
X_22381_ _22381_/A vssd1 vssd1 vccd1 vccd1 _22381_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24120_ _26927_/Q _23571_/X _24120_/S vssd1 vssd1 vccd1 vccd1 _24121_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21332_ _25475_/Q _21332_/B vssd1 vssd1 vccd1 vccd1 _21332_/X sky130_fd_sc_hd__or2_1
XFILLER_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24051_ _26896_/Q _23574_/X _24059_/S vssd1 vssd1 vccd1 vccd1 _24052_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21263_ _25937_/Q _21202_/X _21261_/Y _21262_/X vssd1 vssd1 vccd1 vccd1 _25937_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_150_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23002_ _26473_/Q _22698_/X _23006_/S vssd1 vssd1 vccd1 vccd1 _23003_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20214_ _27153_/Q _27087_/Q vssd1 vssd1 vccd1 vccd1 _20218_/A sky130_fd_sc_hd__and2_1
XFILLER_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21194_ _21197_/A _21194_/B vssd1 vssd1 vccd1 vccd1 _25934_/D sky130_fd_sc_hd__nor2_1
XFILLER_278_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_249_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20145_ _20118_/A _20126_/A _20126_/B vssd1 vssd1 vccd1 vccd1 _20145_/X sky130_fd_sc_hd__a21bo_1
XFILLER_89_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24953_ _24957_/A vssd1 vssd1 vccd1 vccd1 _24953_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ _21718_/A vssd1 vssd1 vccd1 vccd1 _20076_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23904_ _23747_/X _26831_/Q _23904_/S vssd1 vssd1 vccd1 vccd1 _23905_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24884_ _27128_/Q _24890_/B vssd1 vssd1 vccd1 vccd1 _24884_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26623_ _27299_/CLK _26623_/D vssd1 vssd1 vccd1 vccd1 _26623_/Q sky130_fd_sc_hd__dfxtp_1
X_23835_ _23750_/X _26800_/Q _23843_/S vssd1 vssd1 vccd1 vccd1 _23836_/A sky130_fd_sc_hd__mux2_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26554_ _27297_/CLK _26554_/D vssd1 vssd1 vccd1 vccd1 _26554_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23766_ _23766_/A vssd1 vssd1 vccd1 vccd1 _23766_/X sky130_fd_sc_hd__buf_2
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20978_ _20978_/A _20978_/B _21870_/A vssd1 vssd1 vccd1 vccd1 _20986_/C sky130_fd_sc_hd__and3_1
XFILLER_213_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25505_ _27014_/CLK _25505_/D vssd1 vssd1 vccd1 vccd1 _25505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22717_ _23760_/A vssd1 vssd1 vccd1 vccd1 _22717_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26485_ _27292_/CLK _26485_/D vssd1 vssd1 vccd1 vccd1 _26485_/Q sky130_fd_sc_hd__dfxtp_1
X_23697_ _23696_/X _26751_/Q _23700_/S vssd1 vssd1 vccd1 vccd1 _23698_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_194_wb_clk_i clkbuf_4_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27319_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13450_ _12745_/A _13448_/X _13449_/X vssd1 vssd1 vccd1 vccd1 _13451_/B sky130_fd_sc_hd__o21ai_1
XFILLER_213_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25436_ _25436_/A vssd1 vssd1 vccd1 vccd1 _27313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22648_ _26329_/Q _22647_/X _22657_/S vssd1 vssd1 vccd1 vccd1 _22649_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_123_wb_clk_i clkbuf_4_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27014_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13381_ _19947_/A _17824_/A vssd1 vssd1 vccd1 vccd1 _13381_/Y sky130_fd_sc_hd__nor2_1
X_25367_ _25378_/A vssd1 vssd1 vccd1 vccd1 _25376_/S sky130_fd_sc_hd__clkbuf_4
X_22579_ _22567_/X _22578_/Y _22574_/X vssd1 vssd1 vccd1 vccd1 _26307_/D sky130_fd_sc_hd__a21oi_1
XFILLER_210_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15120_ _15118_/X _15119_/X _15120_/S vssd1 vssd1 vccd1 vccd1 _15120_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24318_ _26997_/Q _26996_/Q _24318_/C vssd1 vssd1 vccd1 vccd1 _24320_/B sky130_fd_sc_hd__and3_1
X_27106_ _27110_/CLK _27106_/D vssd1 vssd1 vccd1 vccd1 _27106_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_181_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25298_ _23754_/X _27252_/Q _25304_/S vssd1 vssd1 vccd1 vccd1 _25299_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27037_ _27137_/CLK _27037_/D vssd1 vssd1 vccd1 vccd1 _27037_/Q sky130_fd_sc_hd__dfxtp_1
X_15051_ _15540_/S vssd1 vssd1 vccd1 vccd1 _15351_/B sky130_fd_sc_hd__clkbuf_4
X_24249_ _26972_/Q _24250_/C _26973_/Q vssd1 vssd1 vccd1 vccd1 _24251_/B sky130_fd_sc_hd__a21oi_1
XFILLER_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14002_ _13085_/A _26398_/Q _14246_/S _14001_/X vssd1 vssd1 vccd1 vccd1 _14002_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18810_ _18810_/A vssd1 vssd1 vccd1 vccd1 _18810_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19790_ _19790_/A _19870_/B vssd1 vssd1 vccd1 vccd1 _19790_/X sky130_fd_sc_hd__or2_1
XFILLER_110_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18741_ _18741_/A vssd1 vssd1 vccd1 vccd1 _18741_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15953_ _12912_/A _15345_/X _12929_/A vssd1 vssd1 vccd1 vccd1 _15953_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput140 dout1[3] vssd1 vssd1 vccd1 vccd1 input140/X sky130_fd_sc_hd__clkbuf_1
XTAP_5362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput151 dout1[4] vssd1 vssd1 vccd1 vccd1 input151/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput162 dout1[5] vssd1 vssd1 vccd1 vccd1 input162/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14904_ _16439_/A _14904_/B _14904_/C vssd1 vssd1 vccd1 vccd1 _14904_/Y sky130_fd_sc_hd__nor3_1
XTAP_5384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput173 irq[11] vssd1 vssd1 vccd1 vccd1 _19620_/C sky130_fd_sc_hd__buf_4
X_18672_ _22368_/A _18672_/B vssd1 vssd1 vccd1 vccd1 _18673_/A sky130_fd_sc_hd__and2_1
XTAP_5395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ _15982_/S _15882_/X _15883_/X _14165_/A vssd1 vssd1 vccd1 vccd1 _15885_/C
+ sky130_fd_sc_hd__o211a_1
Xinput184 irq[7] vssd1 vssd1 vccd1 vccd1 _19623_/C sky130_fd_sc_hd__buf_4
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput195 localMemory_wb_adr_i[14] vssd1 vssd1 vccd1 vccd1 input195/X sky130_fd_sc_hd__clkbuf_1
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17623_ _17653_/A _17623_/B _17623_/C vssd1 vssd1 vccd1 vccd1 _17623_/X sky130_fd_sc_hd__or3_1
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ _16409_/B _15873_/C vssd1 vssd1 vccd1 vccd1 _14835_/Y sky130_fd_sc_hd__nor2_1
XFILLER_236_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _17554_/A vssd1 vssd1 vccd1 vccd1 _17554_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14766_ _14766_/A vssd1 vssd1 vccd1 vccd1 _16517_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16505_ _17197_/A _16492_/X _16496_/X _16504_/X _14683_/X vssd1 vssd1 vccd1 vccd1
+ _16505_/X sky130_fd_sc_hd__a311o_1
X_13717_ _13717_/A _13717_/B _13717_/C vssd1 vssd1 vccd1 vccd1 _13717_/X sky130_fd_sc_hd__or3_1
XFILLER_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17485_ _26245_/Q _17455_/A _21206_/A _25973_/Q vssd1 vssd1 vccd1 vccd1 _17486_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14697_ _14690_/X _14693_/X _16476_/S vssd1 vssd1 vccd1 vccd1 _14697_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19224_ _27157_/Q _19367_/B vssd1 vssd1 vccd1 vccd1 _19224_/X sky130_fd_sc_hd__or2_1
X_16436_ _26807_/Q _26451_/Q _16436_/S vssd1 vssd1 vccd1 vccd1 _16436_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13648_ _13951_/S vssd1 vssd1 vccd1 vccd1 _15931_/S sky130_fd_sc_hd__buf_2
XFILLER_32_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _19155_/A _19155_/B vssd1 vssd1 vccd1 vccd1 _19579_/D sky130_fd_sc_hd__xnor2_2
X_13579_ _25639_/Q _15532_/B _13578_/X _25607_/Q vssd1 vssd1 vccd1 vccd1 _13579_/X
+ sky130_fd_sc_hd__a22o_1
X_16367_ _14724_/A _16296_/Y _16366_/Y _14827_/X vssd1 vssd1 vccd1 vccd1 _19268_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_185_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18106_ _18949_/B vssd1 vssd1 vccd1 vccd1 _19331_/B sky130_fd_sc_hd__clkbuf_2
X_15318_ _15318_/A vssd1 vssd1 vccd1 vccd1 _15318_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16298_ _26933_/Q _16400_/S vssd1 vssd1 vccd1 vccd1 _16298_/X sky130_fd_sc_hd__or2_1
X_19086_ _25617_/Q _18971_/X _19085_/X _19007_/X vssd1 vssd1 vccd1 vccd1 _25617_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_274_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18037_ _18358_/A vssd1 vssd1 vccd1 vccd1 _18037_/X sky130_fd_sc_hd__clkbuf_2
X_15249_ _25620_/Q _14596_/A _15248_/X _14617_/A vssd1 vssd1 vccd1 vccd1 _23581_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_173_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19988_ _19763_/X _19983_/X _20007_/B _19987_/X vssd1 vssd1 vccd1 vccd1 _19988_/Y
+ sky130_fd_sc_hd__o31ai_2
XFILLER_114_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18939_ _18861_/X _18938_/X _15702_/A vssd1 vssd1 vccd1 vccd1 _18940_/B sky130_fd_sc_hd__a21oi_2
XFILLER_268_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_267_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21950_ _21950_/A vssd1 vssd1 vccd1 vccd1 _26090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_255_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20901_ _25838_/Q _20900_/X _20901_/S vssd1 vssd1 vccd1 vccd1 _20902_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_254_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21881_ _24473_/A vssd1 vssd1 vccd1 vccd1 _21881_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23620_ _23620_/A vssd1 vssd1 vccd1 vccd1 _26718_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20832_ _25812_/Q vssd1 vssd1 vccd1 vccd1 _20833_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23551_ _23551_/A vssd1 vssd1 vccd1 vccd1 _26696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20763_ _20774_/A vssd1 vssd1 vccd1 vccd1 _20772_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_196_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_270 _18058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_281 _25812_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22502_ _22502_/A _22502_/B vssd1 vssd1 vccd1 vccd1 _22503_/A sky130_fd_sc_hd__and2_1
XFILLER_35_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_292 _25822_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26270_ _26271_/CLK _26270_/D vssd1 vssd1 vccd1 vccd1 _26270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23482_ _23493_/A vssd1 vssd1 vccd1 vccd1 _23491_/S sky130_fd_sc_hd__buf_4
XFILLER_161_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20694_ _20694_/A _20707_/C vssd1 vssd1 vccd1 vccd1 _20694_/X sky130_fd_sc_hd__or2_1
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25221_ _25221_/A vssd1 vssd1 vccd1 vccd1 _25221_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22433_ _22460_/A vssd1 vssd1 vccd1 vccd1 _22444_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25152_ _27194_/Q _25137_/X _25150_/X _25151_/Y _22380_/X vssd1 vssd1 vccd1 vccd1
+ _27194_/D sky130_fd_sc_hd__o221a_1
X_22364_ _17085_/C _26225_/Q _22376_/S vssd1 vssd1 vccd1 vccd1 _22365_/B sky130_fd_sc_hd__mux2_1
XFILLER_248_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24103_ _26919_/Q _23546_/X _24109_/S vssd1 vssd1 vccd1 vccd1 _24104_/A sky130_fd_sc_hd__mux2_1
X_21315_ _21276_/X _21314_/X _21227_/X vssd1 vssd1 vccd1 vccd1 _21315_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_164_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25083_ _24703_/Y _25070_/X _25081_/Y _25082_/X vssd1 vssd1 vccd1 vccd1 _25083_/X
+ sky130_fd_sc_hd__a31o_1
X_22295_ _26210_/Q _22294_/X _22285_/X _26311_/Q _22286_/X vssd1 vssd1 vccd1 vccd1
+ _22295_/X sky130_fd_sc_hd__a221o_1
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24034_ _24034_/A vssd1 vssd1 vccd1 vccd1 _26888_/D sky130_fd_sc_hd__clkbuf_1
X_21246_ _21277_/A vssd1 vssd1 vccd1 vccd1 _21545_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21177_ _21177_/A vssd1 vssd1 vccd1 vccd1 _25929_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_277_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20128_ _19879_/X _20127_/X _19890_/X vssd1 vssd1 vccd1 vccd1 _20128_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_104_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_265_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25985_ _25985_/CLK _25985_/D vssd1 vssd1 vccd1 vccd1 _25985_/Q sky130_fd_sc_hd__dfxtp_2
X_12950_ _14486_/B vssd1 vssd1 vccd1 vccd1 _14610_/A sky130_fd_sc_hd__buf_2
XFILLER_58_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24936_ _24936_/A _24951_/B vssd1 vssd1 vccd1 vccd1 _24936_/Y sky130_fd_sc_hd__nand2_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20059_ _13641_/B _19914_/X _19774_/B _20089_/A vssd1 vssd1 vccd1 vccd1 _20084_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_261_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12881_ _12822_/A _25473_/Q vssd1 vssd1 vccd1 vccd1 _12962_/C sky130_fd_sc_hd__and2b_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24867_ _20681_/A _19963_/X _24736_/Y _24779_/A vssd1 vssd1 vccd1 vccd1 _24867_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26606_ _27313_/CLK _26606_/D vssd1 vssd1 vccd1 vccd1 _26606_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _23606_/A vssd1 vssd1 vccd1 vccd1 _14620_/Y sky130_fd_sc_hd__inv_2
X_23818_ _23818_/A vssd1 vssd1 vccd1 vccd1 _26792_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24798_ _27105_/Q _24798_/B vssd1 vssd1 vccd1 vccd1 _24798_/Y sky130_fd_sc_hd__nand2_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14551_ _27263_/Q _26456_/Q _14551_/S vssd1 vssd1 vccd1 vccd1 _14551_/X sky130_fd_sc_hd__mux2_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26537_ _27280_/CLK _26537_/D vssd1 vssd1 vccd1 vccd1 _26537_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23749_ _23749_/A vssd1 vssd1 vccd1 vccd1 _26767_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _13485_/X _13500_/X _13501_/X _12755_/A vssd1 vssd1 vccd1 vccd1 _13506_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_198_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _17268_/X _17273_/C _17269_/X vssd1 vssd1 vccd1 vccd1 _17270_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _13179_/A _14480_/X _14481_/X vssd1 vssd1 vccd1 vccd1 _14563_/A sky130_fd_sc_hd__o21a_1
X_26468_ _26468_/CLK _26468_/D vssd1 vssd1 vccd1 vccd1 _26468_/Q sky130_fd_sc_hd__dfxtp_2
X_13433_ _13857_/A vssd1 vssd1 vccd1 vccd1 _13433_/X sky130_fd_sc_hd__clkbuf_2
X_16221_ _16217_/X _16220_/X _16221_/S vssd1 vssd1 vccd1 vccd1 _16221_/X sky130_fd_sc_hd__mux2_1
X_25419_ _25419_/A vssd1 vssd1 vccd1 vccd1 _27305_/D sky130_fd_sc_hd__clkbuf_1
X_26399_ _26433_/CLK _26399_/D vssd1 vssd1 vccd1 vccd1 _26399_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_195_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16152_ _12773_/A _26705_/Q _26833_/Q _16319_/S _15048_/A vssd1 vssd1 vccd1 vccd1
+ _16152_/X sky130_fd_sc_hd__a221o_1
X_13364_ _14741_/A _26855_/Q _25769_/Q _15299_/S _15317_/A vssd1 vssd1 vccd1 vccd1
+ _13364_/X sky130_fd_sc_hd__a221o_1
XFILLER_139_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15103_ _14818_/X _15087_/X _15090_/X _15102_/X vssd1 vssd1 vccd1 vccd1 _15103_/X
+ sky130_fd_sc_hd__a31o_1
X_16083_ _15073_/A _23571_/A _16082_/X _15388_/A vssd1 vssd1 vccd1 vccd1 _16908_/A
+ sky130_fd_sc_hd__o211ai_4
X_13295_ _14452_/S vssd1 vssd1 vccd1 vccd1 _13951_/S sky130_fd_sc_hd__buf_2
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19911_ _19911_/A vssd1 vssd1 vccd1 vccd1 _19911_/X sky130_fd_sc_hd__clkbuf_2
X_15034_ _16305_/A vssd1 vssd1 vccd1 vccd1 _15276_/S sky130_fd_sc_hd__buf_2
XFILLER_107_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_91_wb_clk_i _25501_/CLK vssd1 vssd1 vccd1 vccd1 _25660_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19842_ _19839_/A _19841_/Y _19870_/B vssd1 vssd1 vccd1 vccd1 _19842_/X sky130_fd_sc_hd__mux2_4
XFILLER_3_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_wb_clk_i clkbuf_4_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27252_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19773_ _19881_/A _19770_/X _19771_/X _20637_/A vssd1 vssd1 vccd1 vccd1 _19805_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16985_ _16939_/A _16982_/X _16984_/X vssd1 vssd1 vccd1 vccd1 _16986_/B sky130_fd_sc_hd__o21a_2
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18724_ _18724_/A _18724_/B vssd1 vssd1 vccd1 vccd1 _18725_/B sky130_fd_sc_hd__nor2_1
XFILLER_110_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15936_ _15606_/X _15934_/X _15935_/X _13545_/A vssd1 vssd1 vccd1 vccd1 _15936_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_260_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_280_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18655_ _27111_/Q _18504_/X _18653_/X _18654_/X vssd1 vssd1 vccd1 vccd1 _18655_/X
+ sky130_fd_sc_hd__o22a_2
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15867_ _13207_/A _23555_/A _15866_/Y vssd1 vssd1 vccd1 vccd1 _20034_/A sky130_fd_sc_hd__o21ai_4
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17606_ _15441_/X _17584_/X _17604_/X _17605_/X vssd1 vssd1 vccd1 vccd1 _17607_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14818_ _14818_/A vssd1 vssd1 vccd1 vccd1 _14818_/X sky130_fd_sc_hd__buf_4
XFILLER_280_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18586_ _18630_/A _18586_/B vssd1 vssd1 vccd1 vccd1 _18587_/A sky130_fd_sc_hd__and2_1
X_15798_ _12770_/A _26406_/Q _13431_/X _15797_/X vssd1 vssd1 vccd1 vccd1 _15798_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_212_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17537_ _17534_/X _17556_/B _14240_/X _17536_/X _25905_/Q vssd1 vssd1 vccd1 vccd1
+ _17537_/Y sky130_fd_sc_hd__o32ai_4
X_14749_ _14991_/S vssd1 vssd1 vccd1 vccd1 _14813_/S sky130_fd_sc_hd__buf_2
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17468_ _26249_/Q _17455_/A _17461_/A _25977_/Q vssd1 vssd1 vccd1 vccd1 _17470_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_177_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19207_ _18555_/X _19197_/X _19206_/X vssd1 vssd1 vccd1 vccd1 _19207_/X sky130_fd_sc_hd__a21o_4
XFILLER_34_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16419_ _25896_/Q _16419_/B vssd1 vssd1 vccd1 vccd1 _16419_/X sky130_fd_sc_hd__or2_1
X_17399_ _25550_/Q _25551_/Q _17399_/C vssd1 vssd1 vccd1 vccd1 _17401_/B sky130_fd_sc_hd__and3_1
XFILLER_192_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19138_ _25522_/Q _18559_/X _19135_/X _19137_/X _18574_/X vssd1 vssd1 vccd1 vccd1
+ _19138_/X sky130_fd_sc_hd__o221a_1
XFILLER_157_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19069_ _19069_/A vssd1 vssd1 vccd1 vccd1 _19069_/X sky130_fd_sc_hd__clkbuf_2
Xoutput400 _17049_/X vssd1 vssd1 vccd1 vccd1 din0[31] sky130_fd_sc_hd__buf_2
Xoutput411 _25946_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[10] sky130_fd_sc_hd__buf_2
XFILLER_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21100_ _21100_/A _21100_/B vssd1 vssd1 vccd1 vccd1 _21101_/A sky130_fd_sc_hd__or2_1
Xoutput422 _25956_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[20] sky130_fd_sc_hd__buf_2
XFILLER_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput433 _25966_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[30] sky130_fd_sc_hd__buf_2
X_22080_ _26148_/Q _20935_/X _22088_/S vssd1 vssd1 vccd1 vccd1 _22081_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput444 _12763_/Y vssd1 vssd1 vccd1 vccd1 probe_env[1] sky130_fd_sc_hd__buf_2
Xoutput455 _25738_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[14] sky130_fd_sc_hd__buf_2
XFILLER_160_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput466 _25748_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[24] sky130_fd_sc_hd__buf_2
XFILLER_160_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21031_ _25885_/Q _20923_/X _21037_/S vssd1 vssd1 vccd1 vccd1 _21032_/A sky130_fd_sc_hd__mux2_1
Xoutput477 _25729_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[5] sky130_fd_sc_hd__buf_2
XFILLER_248_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22982_ _26464_/Q _22669_/X _22984_/S vssd1 vssd1 vccd1 vccd1 _22983_/A sky130_fd_sc_hd__mux2_1
X_25770_ _27307_/CLK _25770_/D vssd1 vssd1 vccd1 vccd1 _25770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24721_ _27087_/Q _24701_/X _24719_/Y _24720_/X vssd1 vssd1 vccd1 vccd1 _24722_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_21933_ _20571_/X _26083_/Q _21933_/S vssd1 vssd1 vccd1 vccd1 _21934_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24652_ _24777_/A _24915_/A vssd1 vssd1 vccd1 vccd1 _24654_/A sky130_fd_sc_hd__or2_4
XFILLER_242_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21864_ _26060_/Q _20970_/X _21864_/S vssd1 vssd1 vccd1 vccd1 _21865_/A sky130_fd_sc_hd__mux2_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23603_ _23603_/A vssd1 vssd1 vccd1 vccd1 _23603_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_270_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20815_ _20815_/A vssd1 vssd1 vccd1 vccd1 _25803_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24583_ _27049_/Q _24576_/X _24582_/Y _24580_/X vssd1 vssd1 vccd1 vccd1 _27049_/D
+ sky130_fd_sc_hd__o211a_1
X_21795_ _21851_/A vssd1 vssd1 vccd1 vccd1 _21864_/S sky130_fd_sc_hd__buf_8
XFILLER_249_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_26322_ _26322_/CLK _26322_/D vssd1 vssd1 vccd1 vccd1 _26322_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_223_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23534_ _26691_/Q _23533_/X _23540_/S vssd1 vssd1 vccd1 vccd1 _23535_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20746_ _20542_/X _25770_/Q _20750_/S vssd1 vssd1 vccd1 vccd1 _20747_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26253_ _26257_/CLK _26253_/D vssd1 vssd1 vccd1 vccd1 _26253_/Q sky130_fd_sc_hd__dfxtp_1
X_23465_ _26664_/Q _23076_/X _23469_/S vssd1 vssd1 vccd1 vccd1 _23466_/A sky130_fd_sc_hd__mux2_1
X_20677_ _20677_/A _20683_/B vssd1 vssd1 vccd1 vccd1 _20677_/X sky130_fd_sc_hd__or2_1
XFILLER_183_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25204_ _25225_/A vssd1 vssd1 vccd1 vccd1 _25204_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22416_ _26230_/Q _22416_/B _22416_/C vssd1 vssd1 vccd1 vccd1 _22419_/D sky130_fd_sc_hd__nand3_2
XFILLER_155_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26184_ _26319_/CLK _26184_/D vssd1 vssd1 vccd1 vccd1 _26184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23396_ _23396_/A vssd1 vssd1 vccd1 vccd1 _26633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25135_ _24746_/Y _25124_/X _25134_/Y _17339_/A vssd1 vssd1 vccd1 vccd1 _25135_/X
+ sky130_fd_sc_hd__a31o_1
X_22347_ _22379_/A _17078_/X _26228_/Q vssd1 vssd1 vccd1 vccd1 _22347_/X sky130_fd_sc_hd__a21o_1
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13080_ _26663_/Q _15255_/A _13079_/X _15168_/A vssd1 vssd1 vccd1 vccd1 _13080_/X
+ sky130_fd_sc_hd__o211a_1
X_25066_ _22494_/A _25065_/X _25060_/X _18678_/A _25052_/X vssd1 vssd1 vccd1 vccd1
+ _25066_/X sky130_fd_sc_hd__a221o_1
X_22278_ _26205_/Q _22269_/X _22277_/X _22273_/X vssd1 vssd1 vccd1 vccd1 _26205_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24017_ _24074_/S vssd1 vssd1 vccd1 vccd1 _24026_/S sky130_fd_sc_hd__clkbuf_4
X_21229_ _25867_/Q vssd1 vssd1 vccd1 vccd1 _21552_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_278_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16770_ _16770_/A vssd1 vssd1 vccd1 vccd1 _16770_/X sky130_fd_sc_hd__clkbuf_2
X_13982_ _13085_/A _26882_/Q _26754_/Q _13043_/A vssd1 vssd1 vccd1 vccd1 _13982_/X
+ sky130_fd_sc_hd__a22o_1
X_25968_ _27227_/CLK _25968_/D vssd1 vssd1 vccd1 vccd1 _25968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_265_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15721_ _25707_/Q _15984_/B vssd1 vssd1 vccd1 vccd1 _15721_/X sky130_fd_sc_hd__or2_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12933_ _14131_/A _12933_/B vssd1 vssd1 vccd1 vccd1 _13559_/B sky130_fd_sc_hd__nor2_1
X_24919_ _27137_/Q _24902_/X _24918_/Y vssd1 vssd1 vccd1 vccd1 _27137_/D sky130_fd_sc_hd__o21a_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25899_ _27293_/CLK _25899_/D vssd1 vssd1 vccd1 vccd1 _25899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18440_ _18440_/A vssd1 vssd1 vccd1 vccd1 _18441_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _26536_/Q _26144_/Q _15653_/S vssd1 vssd1 vccd1 vccd1 _15652_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12864_ _25599_/Q _25598_/Q vssd1 vssd1 vccd1 vccd1 _12942_/A sky130_fd_sc_hd__or2_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14603_ _14603_/A vssd1 vssd1 vccd1 vccd1 _14604_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18371_ _18371_/A vssd1 vssd1 vccd1 vccd1 _18371_/X sky130_fd_sc_hd__buf_4
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _26081_/Q _25886_/Q _16176_/S vssd1 vssd1 vccd1 vccd1 _15583_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _12808_/A _25569_/Q vssd1 vssd1 vccd1 vccd1 _17129_/A sky130_fd_sc_hd__nand2_1
XFILLER_215_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _25526_/Q _25527_/Q _17322_/C vssd1 vssd1 vccd1 vccd1 _17324_/B sky130_fd_sc_hd__and3_1
XFILLER_18_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14534_ _13941_/A _14532_/X _14533_/X _13945_/A vssd1 vssd1 vccd1 vccd1 _14535_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17253_ _25505_/Q _25506_/Q _17253_/C vssd1 vssd1 vccd1 vccd1 _17256_/B sky130_fd_sc_hd__and3_1
X_14465_ _13937_/A _25830_/Q _26030_/Q _16021_/S _13336_/A vssd1 vssd1 vccd1 vccd1
+ _14465_/X sky130_fd_sc_hd__a221o_1
XFILLER_186_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16204_ _25745_/Q _20227_/A _16204_/S vssd1 vssd1 vccd1 vccd1 _16206_/B sky130_fd_sc_hd__mux2_2
X_13416_ _26854_/Q _25768_/Q _13719_/A vssd1 vssd1 vccd1 vccd1 _13416_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14396_ _13545_/A _14379_/X _14395_/X vssd1 vssd1 vccd1 vccd1 _14396_/X sky130_fd_sc_hd__a21o_1
X_17184_ _16493_/S _17170_/X _17183_/X _17175_/X vssd1 vssd1 vccd1 vccd1 _25488_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13347_ _13347_/A vssd1 vssd1 vccd1 vccd1 _15308_/S sky130_fd_sc_hd__clkbuf_8
X_16135_ _26929_/Q _16135_/B vssd1 vssd1 vccd1 vccd1 _16135_/X sky130_fd_sc_hd__or2_1
XFILLER_6_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13278_ _13278_/A vssd1 vssd1 vccd1 vccd1 _15859_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16066_ _26799_/Q _26443_/Q _16069_/S vssd1 vssd1 vccd1 vccd1 _16066_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15017_ _26934_/Q _16385_/S vssd1 vssd1 vccd1 vccd1 _15017_/X sky130_fd_sc_hd__or2_1
XFILLER_284_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19825_ _19882_/B _18531_/X _19671_/A _19824_/Y vssd1 vssd1 vccd1 vccd1 _19825_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_97_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_271_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19756_ _19748_/X _19754_/X _19755_/X vssd1 vssd1 vccd1 vccd1 _19756_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16968_ _16983_/A _16973_/B _16968_/C vssd1 vssd1 vccd1 vccd1 _16968_/X sky130_fd_sc_hd__and3_1
XFILLER_272_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18707_ _25735_/Q vssd1 vssd1 vccd1 vccd1 _19946_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_225_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15919_ _13254_/A _26109_/Q _26010_/Q _16113_/A _15769_/A vssd1 vssd1 vccd1 vccd1
+ _15919_/X sky130_fd_sc_hd__a221o_1
XFILLER_209_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19687_ _19687_/A _19687_/B vssd1 vssd1 vccd1 vccd1 _19687_/Y sky130_fd_sc_hd__nor2_1
X_16899_ _16924_/A _16899_/B vssd1 vssd1 vccd1 vccd1 _16900_/A sky130_fd_sc_hd__and2_1
XFILLER_253_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18638_ _16735_/X _19354_/B _18637_/X vssd1 vssd1 vccd1 vccd1 _18638_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_252_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18569_ _18569_/A vssd1 vssd1 vccd1 vccd1 _18569_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_206_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20600_ _23594_/A vssd1 vssd1 vccd1 vccd1 _23770_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_21580_ _21580_/A vssd1 vssd1 vccd1 vccd1 _21580_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20531_ _20531_/A vssd1 vssd1 vccd1 vccd1 _25701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23250_ _23250_/A vssd1 vssd1 vccd1 vccd1 _26568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20462_ _19683_/X _20461_/X _19718_/X vssd1 vssd1 vccd1 vccd1 _20462_/X sky130_fd_sc_hd__a21o_1
XFILLER_146_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22201_ _22249_/A vssd1 vssd1 vccd1 vccd1 _22201_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_180_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23181_ _26538_/Q _23095_/X _23183_/S vssd1 vssd1 vccd1 vccd1 _23182_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20393_ _19683_/X _20392_/X _19718_/X vssd1 vssd1 vccd1 vccd1 _20393_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22132_ _22195_/A vssd1 vssd1 vccd1 vccd1 _22132_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22063_ _22063_/A vssd1 vssd1 vccd1 vccd1 _26140_/D sky130_fd_sc_hd__clkbuf_1
X_26940_ _26940_/CLK _26940_/D vssd1 vssd1 vccd1 vccd1 _26940_/Q sky130_fd_sc_hd__dfxtp_4
Xoutput285 _17062_/X vssd1 vssd1 vccd1 vccd1 addr0[0] sky130_fd_sc_hd__buf_2
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21014_ _21014_/A vssd1 vssd1 vccd1 vccd1 _25877_/D sky130_fd_sc_hd__clkbuf_1
Xoutput296 _16993_/X vssd1 vssd1 vccd1 vccd1 addr1[2] sky130_fd_sc_hd__buf_2
XINSDIODE2_3 _22368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26871_ _27319_/CLK _26871_/D vssd1 vssd1 vccd1 vccd1 _26871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_275_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25822_ _26715_/CLK _25822_/D vssd1 vssd1 vccd1 vccd1 _25822_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_114_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_263_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22965_ _26456_/Q _22640_/X _22973_/S vssd1 vssd1 vccd1 vccd1 _22966_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25753_ _26292_/CLK _25753_/D vssd1 vssd1 vccd1 vccd1 _25753_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24704_ _27083_/Q _24701_/X _24703_/Y _24697_/X vssd1 vssd1 vccd1 vccd1 _24705_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_271_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21916_ _20538_/X _26075_/Q _21922_/S vssd1 vssd1 vccd1 vccd1 _21917_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22896_ _22896_/A vssd1 vssd1 vccd1 vccd1 _26425_/D sky130_fd_sc_hd__clkbuf_1
X_25684_ _26286_/CLK _25684_/D vssd1 vssd1 vccd1 vccd1 _25684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_270_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21847_ _26052_/Q _20945_/X _21849_/S vssd1 vssd1 vccd1 vccd1 _21848_/A sky130_fd_sc_hd__mux2_1
X_24635_ _24635_/A vssd1 vssd1 vccd1 vccd1 _24636_/A sky130_fd_sc_hd__buf_2
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24566_ _24630_/A vssd1 vssd1 vccd1 vccd1 _24619_/A sky130_fd_sc_hd__buf_2
X_21778_ _21778_/A vssd1 vssd1 vccd1 vccd1 _21787_/S sky130_fd_sc_hd__buf_6
X_26305_ _26307_/CLK _26305_/D vssd1 vssd1 vccd1 vccd1 _26305_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_11_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20729_ _20729_/A vssd1 vssd1 vccd1 vccd1 _25762_/D sky130_fd_sc_hd__clkbuf_1
X_23517_ _23517_/A vssd1 vssd1 vccd1 vccd1 _23517_/X sky130_fd_sc_hd__buf_2
X_24497_ _24739_/B vssd1 vssd1 vccd1 vccd1 _24611_/A sky130_fd_sc_hd__inv_2
X_27285_ _27285_/CLK _27285_/D vssd1 vssd1 vccd1 vccd1 _27285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_278_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14250_ _13134_/A _14247_/X _14249_/X _13857_/A vssd1 vssd1 vccd1 vccd1 _14250_/X
+ sky130_fd_sc_hd__a211o_1
X_26236_ _26520_/CLK _26236_/D vssd1 vssd1 vccd1 vccd1 _26236_/Q sky130_fd_sc_hd__dfxtp_4
X_23448_ _23448_/A vssd1 vssd1 vccd1 vccd1 _26656_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13201_ _13773_/A _22817_/C _20485_/A _13209_/A vssd1 vssd1 vccd1 vccd1 _13201_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14181_ _14330_/A _14179_/X _14180_/X _14111_/A vssd1 vssd1 vccd1 vccd1 _14181_/X
+ sky130_fd_sc_hd__a211o_1
X_26167_ _27264_/CLK _26167_/D vssd1 vssd1 vccd1 vccd1 _26167_/Q sky130_fd_sc_hd__dfxtp_1
X_23379_ _23379_/A vssd1 vssd1 vccd1 vccd1 _26625_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13132_ _14515_/S vssd1 vssd1 vccd1 vccd1 _14330_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_25118_ _27187_/Q _25112_/X _25117_/X vssd1 vssd1 vccd1 vccd1 _27187_/D sky130_fd_sc_hd__o21ba_1
X_26098_ _26240_/CLK _26098_/D vssd1 vssd1 vccd1 vccd1 _26098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13063_ _14264_/S vssd1 vssd1 vccd1 vccd1 _14246_/S sky130_fd_sc_hd__buf_2
X_17940_ _17935_/X _17939_/X _18071_/S vssd1 vssd1 vccd1 vccd1 _17940_/X sky130_fd_sc_hd__mux2_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25049_ _20643_/A _25031_/X _25048_/X vssd1 vssd1 vccd1 vccd1 _25049_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17871_ _17871_/A vssd1 vssd1 vccd1 vccd1 _18058_/S sky130_fd_sc_hd__buf_2
XFILLER_120_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19610_ _26061_/Q vssd1 vssd1 vccd1 vccd1 _19616_/B sky130_fd_sc_hd__clkbuf_1
X_16822_ _16822_/A vssd1 vssd1 vccd1 vccd1 _16822_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19541_ _19541_/A vssd1 vssd1 vccd1 vccd1 _19541_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16753_ _25677_/Q vssd1 vssd1 vccd1 vccd1 _22507_/A sky130_fd_sc_hd__buf_2
X_13965_ _15760_/A _13961_/X _13964_/X _13529_/A vssd1 vssd1 vccd1 vccd1 _13965_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_219_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15704_ _15704_/A _15871_/A vssd1 vssd1 vccd1 vccd1 _15704_/Y sky130_fd_sc_hd__nand2_1
X_12916_ _13922_/B vssd1 vssd1 vccd1 vccd1 _12916_/X sky130_fd_sc_hd__clkbuf_2
X_19472_ _19472_/A _19472_/B vssd1 vssd1 vccd1 vccd1 _19472_/Y sky130_fd_sc_hd__nor2_1
XFILLER_250_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16684_ _25688_/Q vssd1 vssd1 vccd1 vccd1 _22530_/A sky130_fd_sc_hd__inv_2
XFILLER_94_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13896_ _26527_/Q _26135_/Q _14253_/S vssd1 vssd1 vccd1 vccd1 _13896_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18423_ _18423_/A _18423_/B vssd1 vssd1 vccd1 vccd1 _19572_/B sky130_fd_sc_hd__xnor2_2
X_15635_ _25885_/Q _15635_/B vssd1 vssd1 vccd1 vccd1 _15635_/X sky130_fd_sc_hd__or2_1
XFILLER_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _25599_/Q vssd1 vssd1 vccd1 vccd1 _12872_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _17986_/A _14570_/B _18328_/A _16717_/A vssd1 vssd1 vccd1 vccd1 _18354_/Y
+ sky130_fd_sc_hd__a211oi_1
X_15566_ _26113_/Q _26014_/Q _15566_/S vssd1 vssd1 vccd1 vccd1 _15566_/X sky130_fd_sc_hd__mux2_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _17712_/B _12778_/B vssd1 vssd1 vccd1 vccd1 _25113_/A sky130_fd_sc_hd__or2_4
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _25522_/Q _17305_/B vssd1 vssd1 vccd1 vccd1 _17312_/C sky130_fd_sc_hd__and2_1
XFILLER_175_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14517_ _13083_/A _26684_/Q _26812_/Q _14332_/S vssd1 vssd1 vccd1 vccd1 _14517_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18285_ _18285_/A vssd1 vssd1 vccd1 vccd1 _18285_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15497_ _26506_/Q _26378_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15498_/B sky130_fd_sc_hd__mux2_1
XFILLER_175_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17236_ _17242_/A _17242_/B _17235_/X vssd1 vssd1 vccd1 vccd1 _17236_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14448_ _27264_/Q _26457_/Q _14452_/S vssd1 vssd1 vccd1 vccd1 _14448_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17167_ _18077_/A vssd1 vssd1 vccd1 vccd1 _19392_/A sky130_fd_sc_hd__buf_4
X_14379_ _13543_/A _14368_/X _14371_/X _14378_/X vssd1 vssd1 vccd1 vccd1 _14379_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_116_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16118_ _16105_/X _16108_/X _16117_/Y vssd1 vssd1 vccd1 vccd1 _16118_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17098_ _26224_/Q _22239_/A _17088_/X _17094_/X _22230_/C vssd1 vssd1 vccd1 vccd1
+ _17098_/X sky130_fd_sc_hd__o221a_1
XFILLER_143_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16049_ _27314_/Q _26571_/Q _16053_/S vssd1 vssd1 vccd1 vccd1 _16049_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19808_ _19808_/A _19808_/B vssd1 vssd1 vccd1 vccd1 _19830_/B sky130_fd_sc_hd__nand2_1
XFILLER_257_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19739_ _19725_/X _19737_/X _19738_/X vssd1 vssd1 vccd1 vccd1 _19745_/A sky130_fd_sc_hd__a21o_1
X_22750_ _26361_/Q _22647_/X _22756_/S vssd1 vssd1 vccd1 vccd1 _22751_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21701_ _25989_/Q _17456_/B _21707_/S vssd1 vssd1 vccd1 vccd1 _21702_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22681_ _22681_/A vssd1 vssd1 vccd1 vccd1 _26339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24420_ _27014_/Q _24391_/X _24419_/Y _24415_/X vssd1 vssd1 vccd1 vccd1 _27014_/D
+ sky130_fd_sc_hd__o211a_1
X_21632_ _21630_/Y _21631_/X _21589_/X vssd1 vssd1 vccd1 vccd1 _21632_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24351_ _26940_/Q _24351_/B vssd1 vssd1 vccd1 vccd1 _24351_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21563_ _21563_/A vssd1 vssd1 vccd1 vccd1 _21563_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23302_ _20508_/X _26592_/Q _23302_/S vssd1 vssd1 vccd1 vccd1 _23303_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20514_ _20512_/X _25697_/Q _20530_/S vssd1 vssd1 vccd1 vccd1 _20515_/A sky130_fd_sc_hd__mux2_1
X_27070_ _27203_/CLK _27070_/D vssd1 vssd1 vccd1 vccd1 _27070_/Q sky130_fd_sc_hd__dfxtp_1
X_24282_ _26984_/Q _24284_/C _24281_/Y vssd1 vssd1 vccd1 vccd1 _26984_/D sky130_fd_sc_hd__o21a_1
X_21494_ _25954_/Q _21443_/X _21493_/Y _21467_/X vssd1 vssd1 vccd1 vccd1 _25954_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_154_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23233_ _26561_/Q _23066_/X _23233_/S vssd1 vssd1 vccd1 vccd1 _23234_/A sky130_fd_sc_hd__mux2_1
X_26021_ _27329_/A _26021_/D vssd1 vssd1 vccd1 vccd1 _26021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20445_ _19442_/A _18092_/A _19422_/X _20328_/X vssd1 vssd1 vccd1 vccd1 _20445_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_180_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23164_ _26530_/Q _23069_/X _23172_/S vssd1 vssd1 vccd1 vccd1 _23165_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20376_ _20376_/A vssd1 vssd1 vccd1 vccd1 _20376_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22115_ _22206_/A vssd1 vssd1 vccd1 vccd1 _22115_/X sky130_fd_sc_hd__buf_2
XFILLER_192_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23095_ _23568_/A vssd1 vssd1 vccd1 vccd1 _23095_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_148_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27203_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22046_ _22103_/S vssd1 vssd1 vccd1 vccd1 _22055_/S sky130_fd_sc_hd__clkbuf_4
X_26923_ _27311_/CLK _26923_/D vssd1 vssd1 vccd1 vccd1 _26923_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26854_ _27278_/CLK _26854_/D vssd1 vssd1 vccd1 vccd1 _26854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_13_0_wb_clk_i _25501_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_13_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25805_ _26917_/CLK _25805_/D vssd1 vssd1 vccd1 vccd1 _25805_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_217_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26785_ _27301_/CLK _26785_/D vssd1 vssd1 vccd1 vccd1 _26785_/Q sky130_fd_sc_hd__dfxtp_1
X_23997_ _23997_/A vssd1 vssd1 vccd1 vccd1 _26872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_263_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_284_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13750_ _12871_/A _13740_/Y _13745_/Y _14486_/C _13575_/X vssd1 vssd1 vccd1 vccd1
+ _13750_/X sky130_fd_sc_hd__o32a_1
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25736_ _25737_/CLK _25736_/D vssd1 vssd1 vccd1 vccd1 _25736_/Q sky130_fd_sc_hd__dfxtp_4
X_22948_ _26449_/Q _22723_/X _22956_/S vssd1 vssd1 vccd1 vccd1 _22949_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12701_ _14362_/A vssd1 vssd1 vccd1 vccd1 _12702_/A sky130_fd_sc_hd__buf_4
XFILLER_188_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13681_ _14777_/A _13674_/X _13680_/X _13367_/A vssd1 vssd1 vccd1 vccd1 _13681_/X
+ sky130_fd_sc_hd__o31a_1
X_25667_ _25670_/CLK _25667_/D vssd1 vssd1 vccd1 vccd1 _25667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22879_ _22879_/A vssd1 vssd1 vccd1 vccd1 _26418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15420_ _15406_/X _26116_/Q _26017_/Q _16440_/S _15417_/A vssd1 vssd1 vccd1 vccd1
+ _15420_/X sky130_fd_sc_hd__a221o_1
XPHY_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24618_ _24974_/A _24621_/B vssd1 vssd1 vccd1 vccd1 _24618_/Y sky130_fd_sc_hd__nand2_1
XPHY_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25598_ _25598_/CLK _25598_/D vssd1 vssd1 vccd1 vccd1 _25598_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15351_ _26928_/Q _15351_/B vssd1 vssd1 vccd1 vccd1 _15351_/X sky130_fd_sc_hd__or2_1
XFILLER_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24549_ _27037_/Q _24546_/X _24548_/Y _24523_/X vssd1 vssd1 vccd1 vccd1 _27037_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14302_ _14300_/X _14301_/X _14309_/S vssd1 vssd1 vccd1 vccd1 _14302_/X sky130_fd_sc_hd__mux2_1
X_18070_ _17937_/X _17933_/X _18070_/S vssd1 vssd1 vccd1 vccd1 _18070_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27268_ _27269_/CLK _27268_/D vssd1 vssd1 vccd1 vccd1 _27268_/Q sky130_fd_sc_hd__dfxtp_1
X_15282_ _26642_/Q _26738_/Q _16325_/S vssd1 vssd1 vccd1 vccd1 _15282_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17021_ _17063_/A vssd1 vssd1 vccd1 vccd1 _17021_/X sky130_fd_sc_hd__clkbuf_2
X_26219_ _26222_/CLK _26219_/D vssd1 vssd1 vccd1 vccd1 _26219_/Q sky130_fd_sc_hd__dfxtp_2
X_14233_ _14566_/A _19728_/A _14232_/X vssd1 vssd1 vccd1 vccd1 _17800_/C sky130_fd_sc_hd__o21a_1
XFILLER_137_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27199_ _27203_/CLK _27199_/D vssd1 vssd1 vccd1 vccd1 _27199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14164_ _13884_/S _14162_/X _14163_/X vssd1 vssd1 vccd1 vccd1 _14165_/B sky130_fd_sc_hd__o21ai_1
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13115_ _15546_/S vssd1 vssd1 vccd1 vccd1 _15031_/A sky130_fd_sc_hd__buf_4
XFILLER_113_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14095_ _14095_/A vssd1 vssd1 vccd1 vccd1 _14265_/S sky130_fd_sc_hd__clkbuf_4
X_18972_ _19218_/A vssd1 vssd1 vccd1 vccd1 _18972_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13046_ _25586_/Q vssd1 vssd1 vccd1 vccd1 _13610_/A sky130_fd_sc_hd__inv_2
X_17923_ _17950_/S vssd1 vssd1 vccd1 vccd1 _17949_/S sky130_fd_sc_hd__buf_2
XFILLER_279_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_285_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17854_ _14831_/A _17779_/Y _17853_/X vssd1 vssd1 vccd1 vccd1 _19452_/B sky130_fd_sc_hd__a21bo_2
XFILLER_227_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16805_ _16785_/Y _16804_/Y _16693_/X vssd1 vssd1 vccd1 vccd1 _16805_/X sky130_fd_sc_hd__a21o_1
XFILLER_226_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17785_ _17846_/C _19276_/A _17784_/Y vssd1 vssd1 vccd1 vccd1 _17785_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14997_ _14995_/X _14996_/X _15004_/S vssd1 vssd1 vccd1 vccd1 _14997_/X sky130_fd_sc_hd__mux2_1
XFILLER_219_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19524_ _19512_/X _18876_/X _19523_/X _19515_/X vssd1 vssd1 vccd1 vccd1 _25644_/D
+ sky130_fd_sc_hd__o211a_1
X_16736_ _22491_/A _16726_/X _16727_/X _16735_/X vssd1 vssd1 vccd1 vccd1 _16736_/X
+ sky130_fd_sc_hd__a22o_1
X_13948_ _26658_/Q _25698_/Q _14221_/S vssd1 vssd1 vccd1 vccd1 _13948_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19455_ _17995_/B _19455_/B _19455_/C vssd1 vssd1 vccd1 vccd1 _19455_/X sky130_fd_sc_hd__and3b_1
X_16667_ _25995_/Q vssd1 vssd1 vccd1 vccd1 _16668_/B sky130_fd_sc_hd__buf_2
XFILLER_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13879_ _26787_/Q _26431_/Q _14008_/S vssd1 vssd1 vccd1 vccd1 _13879_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18406_ _18382_/X _18386_/Y _18405_/X _17671_/X vssd1 vssd1 vccd1 vccd1 _18406_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_201_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15618_ _15245_/X _13744_/X _14604_/A vssd1 vssd1 vccd1 vccd1 _15618_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_179_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19386_ _17443_/B _19218_/X _19384_/Y _19385_/Y _19253_/X vssd1 vssd1 vccd1 vccd1
+ _19386_/X sky130_fd_sc_hd__a221o_2
X_16598_ _16932_/B _16782_/A _16957_/A _17971_/D _16597_/X vssd1 vssd1 vccd1 vccd1
+ _16603_/B sky130_fd_sc_hd__o221a_1
XFILLER_194_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18337_ _18337_/A vssd1 vssd1 vccd1 vccd1 _25602_/D sky130_fd_sc_hd__clkbuf_1
X_15549_ _25886_/Q _16061_/B vssd1 vssd1 vccd1 vccd1 _15549_/X sky130_fd_sc_hd__or2_1
XFILLER_188_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18268_ _18260_/X _18267_/X _18685_/S vssd1 vssd1 vccd1 vccd1 _18269_/B sky130_fd_sc_hd__mux2_2
XFILLER_163_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17219_ _17219_/A _17224_/B vssd1 vssd1 vccd1 vccd1 _17219_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18199_ _18196_/X _18197_/X _18348_/S vssd1 vssd1 vccd1 vccd1 _18199_/X sky130_fd_sc_hd__mux2_1
X_20230_ _20299_/A _20259_/B vssd1 vssd1 vccd1 vccd1 _20300_/B sky130_fd_sc_hd__xnor2_1
XFILLER_116_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20161_ _27151_/Q _20160_/X _20371_/S vssd1 vssd1 vccd1 vccd1 _20161_/X sky130_fd_sc_hd__mux2_2
XFILLER_226_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20092_ _20092_/A _20092_/B vssd1 vssd1 vccd1 vccd1 _20376_/A sky130_fd_sc_hd__nor2_2
XFILLER_276_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23920_ _23770_/X _26838_/Q _23926_/S vssd1 vssd1 vccd1 vccd1 _23921_/A sky130_fd_sc_hd__mux2_1
XFILLER_257_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23851_ _23851_/A vssd1 vssd1 vccd1 vccd1 _26807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_22802_ _22802_/A vssd1 vssd1 vccd1 vccd1 _22811_/S sky130_fd_sc_hd__buf_4
X_26570_ _27313_/CLK _26570_/D vssd1 vssd1 vccd1 vccd1 _26570_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23782_ _23782_/A vssd1 vssd1 vccd1 vccd1 _23782_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20994_ _21050_/A vssd1 vssd1 vccd1 vccd1 _21063_/S sky130_fd_sc_hd__buf_6
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25521_ _27022_/CLK _25521_/D vssd1 vssd1 vccd1 vccd1 _25521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22733_ _23776_/A vssd1 vssd1 vccd1 vccd1 _22733_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22664_ _26334_/Q _22663_/X _22673_/S vssd1 vssd1 vccd1 vccd1 _22665_/A sky130_fd_sc_hd__mux2_1
X_25452_ _25452_/A vssd1 vssd1 vccd1 vccd1 _27320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24403_ _27011_/Q _24391_/X _24402_/Y _24379_/X vssd1 vssd1 vccd1 vccd1 _27011_/D
+ sky130_fd_sc_hd__o211a_1
X_21615_ input63/X input99/X _21615_/S vssd1 vssd1 vccd1 vccd1 _21616_/A sky130_fd_sc_hd__mux2_8
XFILLER_197_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22595_ _26313_/Q _22604_/B vssd1 vssd1 vccd1 vccd1 _22595_/Y sky130_fd_sc_hd__nand2_1
X_25383_ _27290_/Q _23773_/A _25387_/S vssd1 vssd1 vccd1 vccd1 _25384_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_27122_ _27122_/CLK _27122_/D vssd1 vssd1 vccd1 vccd1 _27122_/Q sky130_fd_sc_hd__dfxtp_4
X_24334_ _27003_/Q _24334_/B vssd1 vssd1 vccd1 vccd1 _24335_/B sky130_fd_sc_hd__and2_1
X_21546_ _25491_/Q _21574_/B vssd1 vssd1 vccd1 vccd1 _21546_/X sky130_fd_sc_hd__or2_1
XFILLER_194_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24265_ _26978_/Q _24266_/C _26979_/Q vssd1 vssd1 vccd1 vccd1 _24267_/B sky130_fd_sc_hd__a21oi_1
X_27053_ _27062_/CLK _27053_/D vssd1 vssd1 vccd1 vccd1 _27053_/Q sky130_fd_sc_hd__dfxtp_2
X_21477_ _21421_/X _21462_/X _21476_/Y _21451_/X vssd1 vssd1 vccd1 vccd1 _21477_/X
+ sky130_fd_sc_hd__a31o_1
X_26004_ _26595_/CLK _26004_/D vssd1 vssd1 vccd1 vccd1 _26004_/Q sky130_fd_sc_hd__dfxtp_1
X_23216_ _26553_/Q _23041_/X _23222_/S vssd1 vssd1 vccd1 vccd1 _23217_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20428_ _19796_/X _20427_/X _19890_/X vssd1 vssd1 vccd1 vccd1 _20428_/X sky130_fd_sc_hd__a21o_1
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24196_ _26955_/Q _24197_/C _24195_/Y vssd1 vssd1 vccd1 vccd1 _26955_/D sky130_fd_sc_hd__o21a_1
XFILLER_107_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23147_ _23147_/A vssd1 vssd1 vccd1 vccd1 _26522_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20359_ _20359_/A _20399_/A vssd1 vssd1 vccd1 vccd1 _20398_/A sky130_fd_sc_hd__xnor2_1
XFILLER_106_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23078_ _23078_/A vssd1 vssd1 vccd1 vccd1 _26500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14920_ _14794_/A _14915_/X _14919_/X _17181_/A vssd1 vssd1 vccd1 vccd1 _14920_/X
+ sky130_fd_sc_hd__o211a_1
X_26906_ _27259_/CLK _26906_/D vssd1 vssd1 vccd1 vccd1 _26906_/Q sky130_fd_sc_hd__dfxtp_1
X_22029_ _26126_/Q _20967_/X _22031_/S vssd1 vssd1 vccd1 vccd1 _22030_/A sky130_fd_sc_hd__mux2_1
XTAP_5544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26837_ _27253_/CLK _26837_/D vssd1 vssd1 vccd1 vccd1 _26837_/Q sky130_fd_sc_hd__dfxtp_1
X_14851_ _25826_/Q _14963_/S _14969_/S _14850_/X vssd1 vssd1 vccd1 vccd1 _14851_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13802_ _12835_/Y _15704_/A _12849_/X _12857_/X vssd1 vssd1 vccd1 vccd1 _13802_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_21_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17570_ _25574_/Q _17564_/X _17540_/X _17569_/X vssd1 vssd1 vccd1 vccd1 _17571_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26768_ _27253_/CLK _26768_/D vssd1 vssd1 vccd1 vccd1 _26768_/Q sky130_fd_sc_hd__dfxtp_1
X_14782_ _16517_/A _14780_/X _14781_/X _12758_/A vssd1 vssd1 vccd1 vccd1 _14782_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_189_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16521_ _16521_/A _16521_/B _16521_/C vssd1 vssd1 vccd1 vccd1 _16521_/X sky130_fd_sc_hd__or3_1
XFILLER_232_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13733_ _14647_/A _13729_/X _13732_/X _13114_/A vssd1 vssd1 vccd1 vccd1 _13733_/X
+ sky130_fd_sc_hd__o211a_1
X_25719_ _27322_/CLK _25719_/D vssd1 vssd1 vccd1 vccd1 _25719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26699_ _27311_/CLK _26699_/D vssd1 vssd1 vccd1 vccd1 _26699_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _27330_/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_188_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19240_ _18213_/X _18734_/X _19240_/S vssd1 vssd1 vccd1 vccd1 _19240_/X sky130_fd_sc_hd__mux2_1
X_16452_ _16453_/A _17780_/B vssd1 vssd1 vccd1 vccd1 _19322_/A sky130_fd_sc_hd__and2_1
X_13664_ _13664_/A vssd1 vssd1 vccd1 vccd1 _15588_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_232_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15403_ _26508_/Q _26380_/Q _16256_/B vssd1 vssd1 vccd1 vccd1 _15404_/B sky130_fd_sc_hd__mux2_1
X_19171_ _17308_/X _18810_/X _19168_/X _19170_/X _18832_/X vssd1 vssd1 vccd1 vccd1
+ _19171_/X sky130_fd_sc_hd__o221a_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16383_ _14661_/A _16378_/X _16382_/X _14623_/A vssd1 vssd1 vccd1 vccd1 _16383_/X
+ sky130_fd_sc_hd__o211a_1
X_13595_ _13410_/X _13589_/X _13594_/X _13159_/A vssd1 vssd1 vccd1 vccd1 _13595_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18122_ _18823_/A vssd1 vssd1 vccd1 vccd1 _19066_/A sky130_fd_sc_hd__buf_2
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15334_ _15313_/A _15330_/X _15332_/X _15333_/X vssd1 vssd1 vccd1 vccd1 _15334_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_61_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18053_ _18051_/X _18052_/X _18254_/A vssd1 vssd1 vccd1 vccd1 _18053_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15265_ _15633_/S vssd1 vssd1 vccd1 vccd1 _15265_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_184_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17004_ _16784_/X _17001_/X _16841_/B _17003_/X input215/X vssd1 vssd1 vccd1 vccd1
+ _17004_/X sky130_fd_sc_hd__a32o_4
X_14216_ _14214_/X _14215_/X _14223_/S vssd1 vssd1 vccd1 vccd1 _14216_/X sky130_fd_sc_hd__mux2_1
X_15196_ _15758_/S vssd1 vssd1 vccd1 vccd1 _15197_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14147_ _14147_/A _14147_/B vssd1 vssd1 vccd1 vccd1 _23523_/A sky130_fd_sc_hd__nand2_4
XFILLER_258_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18955_ _26957_/Q _18569_/A _18570_/A _26989_/Q vssd1 vssd1 vccd1 vccd1 _18955_/X
+ sky130_fd_sc_hd__a22o_1
X_14078_ _13976_/X _14059_/X _14077_/X _13509_/A vssd1 vssd1 vccd1 vccd1 _14078_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_239_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13029_ _13029_/A vssd1 vssd1 vccd1 vccd1 _15885_/A sky130_fd_sc_hd__buf_2
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17906_ _17819_/B _15342_/B _17954_/S vssd1 vssd1 vccd1 vccd1 _17906_/X sky130_fd_sc_hd__mux2_1
X_18886_ _18967_/A _18886_/B vssd1 vssd1 vccd1 vccd1 _18886_/Y sky130_fd_sc_hd__nand2_2
XFILLER_267_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17837_ _17837_/A _15701_/B vssd1 vssd1 vccd1 vccd1 _17837_/X sky130_fd_sc_hd__or2b_1
XFILLER_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17768_ _17673_/X _17764_/X _17767_/X vssd1 vssd1 vccd1 vccd1 _17768_/X sky130_fd_sc_hd__a21o_1
XFILLER_242_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19507_ _19499_/X _18524_/X _19506_/X _19502_/X vssd1 vssd1 vccd1 vccd1 _25637_/D
+ sky130_fd_sc_hd__o211a_1
X_16719_ _25666_/Q vssd1 vssd1 vccd1 vccd1 _22483_/A sky130_fd_sc_hd__buf_4
XFILLER_212_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17699_ _17745_/A vssd1 vssd1 vccd1 vccd1 _17750_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_430 _26234_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_441 _25730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19438_ _26971_/Q _18764_/X _18765_/X _27003_/Q vssd1 vssd1 vccd1 vccd1 _19438_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_211_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_452 _17059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_463 _19072_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_474 _12846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_485 _21195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_496 _16951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19369_ _27065_/Q _18811_/X _19366_/X _19368_/X _18823_/X vssd1 vssd1 vccd1 vccd1
+ _19369_/X sky130_fd_sc_hd__o221a_2
X_21400_ _21597_/A vssd1 vssd1 vccd1 vccd1 _21400_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22380_ _22472_/B vssd1 vssd1 vccd1 vccd1 _22380_/X sky130_fd_sc_hd__buf_8
XFILLER_176_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21331_ _25942_/Q _21310_/X _21329_/Y _21330_/X vssd1 vssd1 vccd1 vccd1 _25942_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_24050_ _24061_/A vssd1 vssd1 vccd1 vccd1 _24059_/S sky130_fd_sc_hd__buf_4
X_21262_ _24871_/A vssd1 vssd1 vccd1 vccd1 _21262_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23001_ _23001_/A vssd1 vssd1 vccd1 vccd1 _26472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20213_ _27121_/Q _20079_/X _20112_/X _20212_/X vssd1 vssd1 vccd1 vccd1 _20213_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21193_ input9/X _16641_/A _21191_/X _21192_/X vssd1 vssd1 vccd1 vccd1 _21194_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_278_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20144_ _20144_/A _20144_/B vssd1 vssd1 vccd1 vccd1 _20200_/A sky130_fd_sc_hd__xnor2_1
XFILLER_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24952_ _27150_/Q _24930_/X _24951_/Y _24949_/X vssd1 vssd1 vccd1 vccd1 _27150_/D
+ sky130_fd_sc_hd__o211a_1
X_20075_ _19894_/X _20074_/X _19902_/X vssd1 vssd1 vccd1 vccd1 _20075_/X sky130_fd_sc_hd__a21o_1
XFILLER_246_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23903_ _23903_/A vssd1 vssd1 vccd1 vccd1 _26830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24883_ _24881_/Y _24882_/X _24871_/X vssd1 vssd1 vccd1 vccd1 _27127_/D sky130_fd_sc_hd__a21oi_1
XFILLER_73_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26622_ _26813_/CLK _26622_/D vssd1 vssd1 vccd1 vccd1 _26622_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23834_ _23845_/A vssd1 vssd1 vccd1 vccd1 _23843_/S sky130_fd_sc_hd__clkbuf_8
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26553_ _27297_/CLK _26553_/D vssd1 vssd1 vccd1 vccd1 _26553_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20977_ _20977_/A _16668_/B vssd1 vssd1 vccd1 vccd1 _21870_/A sky130_fd_sc_hd__or2b_2
X_23765_ _23765_/A vssd1 vssd1 vccd1 vccd1 _26772_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25504_ _27014_/CLK _25504_/D vssd1 vssd1 vccd1 vccd1 _25504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22716_ _22716_/A vssd1 vssd1 vccd1 vccd1 _26350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_281_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26484_ _27291_/CLK _26484_/D vssd1 vssd1 vccd1 vccd1 _26484_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_14_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_23696_ _23696_/A vssd1 vssd1 vccd1 vccd1 _23696_/X sky130_fd_sc_hd__buf_2
XFILLER_202_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25435_ _23744_/X _27313_/Q _25437_/S vssd1 vssd1 vccd1 vccd1 _25436_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22647_ _23690_/A vssd1 vssd1 vccd1 vccd1 _22647_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_198_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13380_ _17824_/B vssd1 vssd1 vccd1 vccd1 _13380_/Y sky130_fd_sc_hd__inv_2
X_22578_ _26307_/Q _22578_/B vssd1 vssd1 vccd1 vccd1 _22578_/Y sky130_fd_sc_hd__nand2_1
X_25366_ _25366_/A vssd1 vssd1 vccd1 vccd1 _27282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27105_ _27110_/CLK _27105_/D vssd1 vssd1 vccd1 vccd1 _27105_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24317_ _26996_/Q _24318_/C _26997_/Q vssd1 vssd1 vccd1 vccd1 _24319_/B sky130_fd_sc_hd__a21oi_1
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21529_ _21488_/X _25864_/Q _21528_/Y _21518_/X vssd1 vssd1 vccd1 vccd1 _21529_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_126_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25297_ _25297_/A vssd1 vssd1 vccd1 vccd1 _27251_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_163_wb_clk_i clkbuf_4_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _25673_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_182_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27036_ _27133_/CLK _27036_/D vssd1 vssd1 vccd1 vccd1 _27036_/Q sky130_fd_sc_hd__dfxtp_1
X_15050_ _15044_/X _15045_/X _15049_/X vssd1 vssd1 vccd1 vccd1 _15050_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24248_ _24291_/A vssd1 vssd1 vccd1 vccd1 _24285_/A sky130_fd_sc_hd__buf_2
XFILLER_154_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14001_ _26914_/Q _14001_/B vssd1 vssd1 vccd1 vccd1 _14001_/X sky130_fd_sc_hd__or2_1
XFILLER_5_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24179_ _24188_/A _24184_/C vssd1 vssd1 vccd1 vccd1 _24179_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18740_ _18805_/A vssd1 vssd1 vccd1 vccd1 _18740_/X sky130_fd_sc_hd__clkbuf_2
XTAP_5330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15952_ _17816_/C vssd1 vssd1 vccd1 vccd1 _18838_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput130 dout1[30] vssd1 vssd1 vccd1 vccd1 input130/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_5352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput141 dout1[40] vssd1 vssd1 vccd1 vccd1 input141/X sky130_fd_sc_hd__clkbuf_2
Xinput152 dout1[50] vssd1 vssd1 vccd1 vccd1 input152/X sky130_fd_sc_hd__clkbuf_2
XTAP_5363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14903_ _14766_/A _14901_/X _14902_/X _12757_/A vssd1 vssd1 vccd1 vccd1 _14904_/C
+ sky130_fd_sc_hd__o211a_1
Xinput163 dout1[60] vssd1 vssd1 vccd1 vccd1 input163/X sky130_fd_sc_hd__clkbuf_2
XTAP_5374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18671_ _13549_/X _18285_/A _18669_/X _18973_/A _25608_/Q vssd1 vssd1 vccd1 vccd1
+ _18672_/B sky130_fd_sc_hd__a32o_1
XFILLER_264_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _13890_/X _26889_/Q _26761_/Q _13706_/A _13049_/A vssd1 vssd1 vccd1 vccd1
+ _15883_/X sky130_fd_sc_hd__a221o_1
XFILLER_237_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput174 irq[12] vssd1 vssd1 vccd1 vccd1 _19611_/C sky130_fd_sc_hd__clkbuf_8
XTAP_5396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput185 irq[8] vssd1 vssd1 vccd1 vccd1 input185/X sky130_fd_sc_hd__buf_4
Xinput196 localMemory_wb_adr_i[15] vssd1 vssd1 vccd1 vccd1 input196/X sky130_fd_sc_hd__clkbuf_1
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17622_ _17633_/A _17622_/B vssd1 vssd1 vccd1 vccd1 _25587_/D sky130_fd_sc_hd__nor2_1
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834_ _14834_/A _14834_/B _14834_/C vssd1 vssd1 vccd1 vccd1 _15873_/C sky130_fd_sc_hd__nor3_1
XFILLER_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_251_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ _17608_/A vssd1 vssd1 vccd1 vccd1 _17553_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14765_ _14765_/A vssd1 vssd1 vccd1 vccd1 _14766_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16504_ _14650_/X _16499_/X _16503_/X _14679_/X vssd1 vssd1 vccd1 vccd1 _16504_/X
+ sky130_fd_sc_hd__o211a_1
X_13716_ _16071_/S _13713_/X _13715_/X _14362_/A _15646_/A vssd1 vssd1 vccd1 vccd1
+ _13717_/C sky130_fd_sc_hd__o2111a_1
XFILLER_204_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17484_ _26246_/Q _17455_/A _21206_/A _25974_/Q vssd1 vssd1 vccd1 vccd1 _21219_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_60_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14696_ _16221_/S vssd1 vssd1 vccd1 vccd1 _16476_/S sky130_fd_sc_hd__buf_4
XFILLER_189_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19223_ _27125_/Q _18504_/A _19221_/X _19222_/X vssd1 vssd1 vccd1 vccd1 _19223_/X
+ sky130_fd_sc_hd__o22a_2
X_16435_ _16336_/X _16433_/X _16434_/X _12755_/A vssd1 vssd1 vccd1 vccd1 _16439_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13647_ _26497_/Q _26369_/Q _15923_/S vssd1 vssd1 vccd1 vccd1 _13647_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19154_ _19121_/B _19122_/B _17792_/X vssd1 vssd1 vccd1 vccd1 _19155_/B sky130_fd_sc_hd__o21ai_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16366_ _16350_/X _16365_/X _14724_/A vssd1 vssd1 vccd1 vccd1 _16366_/Y sky130_fd_sc_hd__a21oi_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _13578_/A vssd1 vssd1 vccd1 vccd1 _13578_/X sky130_fd_sc_hd__clkbuf_2
X_18105_ _18234_/A vssd1 vssd1 vccd1 vccd1 _18949_/B sky130_fd_sc_hd__clkbuf_2
X_15317_ _15317_/A vssd1 vssd1 vccd1 vccd1 _15318_/A sky130_fd_sc_hd__buf_2
XFILLER_9_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19085_ _17444_/D _18972_/X _18973_/X _19084_/Y vssd1 vssd1 vccd1 vccd1 _19085_/X
+ sky130_fd_sc_hd__a211o_1
X_16297_ _27320_/Q _26577_/Q _16301_/S vssd1 vssd1 vccd1 vccd1 _16297_/X sky130_fd_sc_hd__mux2_1
XFILLER_258_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18036_ _18036_/A _18182_/B vssd1 vssd1 vccd1 vccd1 _18358_/A sky130_fd_sc_hd__nor2_2
X_15248_ _14600_/A _15246_/Y _15247_/X _15135_/X vssd1 vssd1 vccd1 vccd1 _15248_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_173_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15179_ _16143_/S vssd1 vssd1 vccd1 vccd1 _16400_/S sky130_fd_sc_hd__buf_4
XFILLER_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19987_ _19657_/X _19985_/X _19986_/Y _19941_/A vssd1 vssd1 vccd1 vccd1 _19987_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18938_ _19192_/B _18686_/B _18938_/S vssd1 vssd1 vccd1 vccd1 _18938_/X sky130_fd_sc_hd__mux2_1
.ends

