VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Video
  CLASS BLOCK ;
  FOREIGN Video ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN sram0_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 20.440 500.000 21.040 ;
    END
  END sram0_csb0
  PIN sram0_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 23.160 500.000 23.760 ;
    END
  END sram0_csb1
  PIN sram0_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 38.120 500.000 38.720 ;
    END
  END sram0_dout0[0]
  PIN sram0_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 221.040 500.000 221.640 ;
    END
  END sram0_dout0[10]
  PIN sram0_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 233.960 500.000 234.560 ;
    END
  END sram0_dout0[11]
  PIN sram0_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 246.200 500.000 246.800 ;
    END
  END sram0_dout0[12]
  PIN sram0_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 259.120 500.000 259.720 ;
    END
  END sram0_dout0[13]
  PIN sram0_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 272.040 500.000 272.640 ;
    END
  END sram0_dout0[14]
  PIN sram0_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 284.280 500.000 284.880 ;
    END
  END sram0_dout0[15]
  PIN sram0_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 297.200 500.000 297.800 ;
    END
  END sram0_dout0[16]
  PIN sram0_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 310.120 500.000 310.720 ;
    END
  END sram0_dout0[17]
  PIN sram0_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 322.360 500.000 322.960 ;
    END
  END sram0_dout0[18]
  PIN sram0_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 335.280 500.000 335.880 ;
    END
  END sram0_dout0[19]
  PIN sram0_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 58.520 500.000 59.120 ;
    END
  END sram0_dout0[1]
  PIN sram0_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 348.200 500.000 348.800 ;
    END
  END sram0_dout0[20]
  PIN sram0_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 360.440 500.000 361.040 ;
    END
  END sram0_dout0[21]
  PIN sram0_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 373.360 500.000 373.960 ;
    END
  END sram0_dout0[22]
  PIN sram0_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 386.280 500.000 386.880 ;
    END
  END sram0_dout0[23]
  PIN sram0_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 398.520 500.000 399.120 ;
    END
  END sram0_dout0[24]
  PIN sram0_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 411.440 500.000 412.040 ;
    END
  END sram0_dout0[25]
  PIN sram0_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 424.360 500.000 424.960 ;
    END
  END sram0_dout0[26]
  PIN sram0_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 436.600 500.000 437.200 ;
    END
  END sram0_dout0[27]
  PIN sram0_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 449.520 500.000 450.120 ;
    END
  END sram0_dout0[28]
  PIN sram0_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 462.440 500.000 463.040 ;
    END
  END sram0_dout0[29]
  PIN sram0_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 78.920 500.000 79.520 ;
    END
  END sram0_dout0[2]
  PIN sram0_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 474.680 500.000 475.280 ;
    END
  END sram0_dout0[30]
  PIN sram0_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 487.600 500.000 488.200 ;
    END
  END sram0_dout0[31]
  PIN sram0_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 99.320 500.000 99.920 ;
    END
  END sram0_dout0[3]
  PIN sram0_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 119.720 500.000 120.320 ;
    END
  END sram0_dout0[4]
  PIN sram0_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 137.400 500.000 138.000 ;
    END
  END sram0_dout0[5]
  PIN sram0_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 155.080 500.000 155.680 ;
    END
  END sram0_dout0[6]
  PIN sram0_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 172.760 500.000 173.360 ;
    END
  END sram0_dout0[7]
  PIN sram0_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 190.440 500.000 191.040 ;
    END
  END sram0_dout0[8]
  PIN sram0_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 208.120 500.000 208.720 ;
    END
  END sram0_dout0[9]
  PIN sram0_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 40.840 500.000 41.440 ;
    END
  END sram0_dout1[0]
  PIN sram0_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 223.760 500.000 224.360 ;
    END
  END sram0_dout1[10]
  PIN sram0_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 236.000 500.000 236.600 ;
    END
  END sram0_dout1[11]
  PIN sram0_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 248.920 500.000 249.520 ;
    END
  END sram0_dout1[12]
  PIN sram0_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 261.840 500.000 262.440 ;
    END
  END sram0_dout1[13]
  PIN sram0_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 274.080 500.000 274.680 ;
    END
  END sram0_dout1[14]
  PIN sram0_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 287.000 500.000 287.600 ;
    END
  END sram0_dout1[15]
  PIN sram0_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 299.920 500.000 300.520 ;
    END
  END sram0_dout1[16]
  PIN sram0_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 312.160 500.000 312.760 ;
    END
  END sram0_dout1[17]
  PIN sram0_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 325.080 500.000 325.680 ;
    END
  END sram0_dout1[18]
  PIN sram0_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 338.000 500.000 338.600 ;
    END
  END sram0_dout1[19]
  PIN sram0_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 61.240 500.000 61.840 ;
    END
  END sram0_dout1[1]
  PIN sram0_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 350.240 500.000 350.840 ;
    END
  END sram0_dout1[20]
  PIN sram0_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 363.160 500.000 363.760 ;
    END
  END sram0_dout1[21]
  PIN sram0_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 376.080 500.000 376.680 ;
    END
  END sram0_dout1[22]
  PIN sram0_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 388.320 500.000 388.920 ;
    END
  END sram0_dout1[23]
  PIN sram0_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 401.240 500.000 401.840 ;
    END
  END sram0_dout1[24]
  PIN sram0_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 414.160 500.000 414.760 ;
    END
  END sram0_dout1[25]
  PIN sram0_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 426.400 500.000 427.000 ;
    END
  END sram0_dout1[26]
  PIN sram0_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 439.320 500.000 439.920 ;
    END
  END sram0_dout1[27]
  PIN sram0_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 452.240 500.000 452.840 ;
    END
  END sram0_dout1[28]
  PIN sram0_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 464.480 500.000 465.080 ;
    END
  END sram0_dout1[29]
  PIN sram0_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 81.640 500.000 82.240 ;
    END
  END sram0_dout1[2]
  PIN sram0_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 477.400 500.000 478.000 ;
    END
  END sram0_dout1[30]
  PIN sram0_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 490.320 500.000 490.920 ;
    END
  END sram0_dout1[31]
  PIN sram0_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 102.040 500.000 102.640 ;
    END
  END sram0_dout1[3]
  PIN sram0_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 122.440 500.000 123.040 ;
    END
  END sram0_dout1[4]
  PIN sram0_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 140.120 500.000 140.720 ;
    END
  END sram0_dout1[5]
  PIN sram0_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 157.800 500.000 158.400 ;
    END
  END sram0_dout1[6]
  PIN sram0_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 175.480 500.000 176.080 ;
    END
  END sram0_dout1[7]
  PIN sram0_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 193.160 500.000 193.760 ;
    END
  END sram0_dout1[8]
  PIN sram0_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 210.840 500.000 211.440 ;
    END
  END sram0_dout1[9]
  PIN sram1_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 25.880 500.000 26.480 ;
    END
  END sram1_csb0
  PIN sram1_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 28.600 500.000 29.200 ;
    END
  END sram1_csb1
  PIN sram1_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 43.560 500.000 44.160 ;
    END
  END sram1_dout0[0]
  PIN sram1_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 226.480 500.000 227.080 ;
    END
  END sram1_dout0[10]
  PIN sram1_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 238.720 500.000 239.320 ;
    END
  END sram1_dout0[11]
  PIN sram1_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 251.640 500.000 252.240 ;
    END
  END sram1_dout0[12]
  PIN sram1_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 264.560 500.000 265.160 ;
    END
  END sram1_dout0[13]
  PIN sram1_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 276.800 500.000 277.400 ;
    END
  END sram1_dout0[14]
  PIN sram1_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 289.720 500.000 290.320 ;
    END
  END sram1_dout0[15]
  PIN sram1_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 301.960 500.000 302.560 ;
    END
  END sram1_dout0[16]
  PIN sram1_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 314.880 500.000 315.480 ;
    END
  END sram1_dout0[17]
  PIN sram1_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 327.800 500.000 328.400 ;
    END
  END sram1_dout0[18]
  PIN sram1_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 340.040 500.000 340.640 ;
    END
  END sram1_dout0[19]
  PIN sram1_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 63.960 500.000 64.560 ;
    END
  END sram1_dout0[1]
  PIN sram1_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 352.960 500.000 353.560 ;
    END
  END sram1_dout0[20]
  PIN sram1_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 365.880 500.000 366.480 ;
    END
  END sram1_dout0[21]
  PIN sram1_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 378.120 500.000 378.720 ;
    END
  END sram1_dout0[22]
  PIN sram1_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 391.040 500.000 391.640 ;
    END
  END sram1_dout0[23]
  PIN sram1_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 403.960 500.000 404.560 ;
    END
  END sram1_dout0[24]
  PIN sram1_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 416.200 500.000 416.800 ;
    END
  END sram1_dout0[25]
  PIN sram1_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 429.120 500.000 429.720 ;
    END
  END sram1_dout0[26]
  PIN sram1_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 442.040 500.000 442.640 ;
    END
  END sram1_dout0[27]
  PIN sram1_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 454.280 500.000 454.880 ;
    END
  END sram1_dout0[28]
  PIN sram1_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 467.200 500.000 467.800 ;
    END
  END sram1_dout0[29]
  PIN sram1_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 84.360 500.000 84.960 ;
    END
  END sram1_dout0[2]
  PIN sram1_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 480.120 500.000 480.720 ;
    END
  END sram1_dout0[30]
  PIN sram1_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 492.360 500.000 492.960 ;
    END
  END sram1_dout0[31]
  PIN sram1_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 104.080 500.000 104.680 ;
    END
  END sram1_dout0[3]
  PIN sram1_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 124.480 500.000 125.080 ;
    END
  END sram1_dout0[4]
  PIN sram1_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 142.160 500.000 142.760 ;
    END
  END sram1_dout0[5]
  PIN sram1_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 160.520 500.000 161.120 ;
    END
  END sram1_dout0[6]
  PIN sram1_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 178.200 500.000 178.800 ;
    END
  END sram1_dout0[7]
  PIN sram1_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 195.880 500.000 196.480 ;
    END
  END sram1_dout0[8]
  PIN sram1_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 213.560 500.000 214.160 ;
    END
  END sram1_dout0[9]
  PIN sram1_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 46.280 500.000 46.880 ;
    END
  END sram1_dout1[0]
  PIN sram1_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 228.520 500.000 229.120 ;
    END
  END sram1_dout1[10]
  PIN sram1_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 241.440 500.000 242.040 ;
    END
  END sram1_dout1[11]
  PIN sram1_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 254.360 500.000 254.960 ;
    END
  END sram1_dout1[12]
  PIN sram1_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 266.600 500.000 267.200 ;
    END
  END sram1_dout1[13]
  PIN sram1_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 279.520 500.000 280.120 ;
    END
  END sram1_dout1[14]
  PIN sram1_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 292.440 500.000 293.040 ;
    END
  END sram1_dout1[15]
  PIN sram1_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 304.680 500.000 305.280 ;
    END
  END sram1_dout1[16]
  PIN sram1_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 317.600 500.000 318.200 ;
    END
  END sram1_dout1[17]
  PIN sram1_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 330.520 500.000 331.120 ;
    END
  END sram1_dout1[18]
  PIN sram1_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 342.760 500.000 343.360 ;
    END
  END sram1_dout1[19]
  PIN sram1_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 66.680 500.000 67.280 ;
    END
  END sram1_dout1[1]
  PIN sram1_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 355.680 500.000 356.280 ;
    END
  END sram1_dout1[20]
  PIN sram1_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 367.920 500.000 368.520 ;
    END
  END sram1_dout1[21]
  PIN sram1_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 380.840 500.000 381.440 ;
    END
  END sram1_dout1[22]
  PIN sram1_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 393.760 500.000 394.360 ;
    END
  END sram1_dout1[23]
  PIN sram1_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 406.000 500.000 406.600 ;
    END
  END sram1_dout1[24]
  PIN sram1_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 418.920 500.000 419.520 ;
    END
  END sram1_dout1[25]
  PIN sram1_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 431.840 500.000 432.440 ;
    END
  END sram1_dout1[26]
  PIN sram1_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 444.080 500.000 444.680 ;
    END
  END sram1_dout1[27]
  PIN sram1_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 457.000 500.000 457.600 ;
    END
  END sram1_dout1[28]
  PIN sram1_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 469.920 500.000 470.520 ;
    END
  END sram1_dout1[29]
  PIN sram1_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 86.400 500.000 87.000 ;
    END
  END sram1_dout1[2]
  PIN sram1_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 482.160 500.000 482.760 ;
    END
  END sram1_dout1[30]
  PIN sram1_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 495.080 500.000 495.680 ;
    END
  END sram1_dout1[31]
  PIN sram1_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 106.800 500.000 107.400 ;
    END
  END sram1_dout1[3]
  PIN sram1_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 127.200 500.000 127.800 ;
    END
  END sram1_dout1[4]
  PIN sram1_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 144.880 500.000 145.480 ;
    END
  END sram1_dout1[5]
  PIN sram1_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 162.560 500.000 163.160 ;
    END
  END sram1_dout1[6]
  PIN sram1_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 180.240 500.000 180.840 ;
    END
  END sram1_dout1[7]
  PIN sram1_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 198.600 500.000 199.200 ;
    END
  END sram1_dout1[8]
  PIN sram1_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 216.280 500.000 216.880 ;
    END
  END sram1_dout1[9]
  PIN sram_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 48.320 500.000 48.920 ;
    END
  END sram_addr0[0]
  PIN sram_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 68.720 500.000 69.320 ;
    END
  END sram_addr0[1]
  PIN sram_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 89.120 500.000 89.720 ;
    END
  END sram_addr0[2]
  PIN sram_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 109.520 500.000 110.120 ;
    END
  END sram_addr0[3]
  PIN sram_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 129.920 500.000 130.520 ;
    END
  END sram_addr0[4]
  PIN sram_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 147.600 500.000 148.200 ;
    END
  END sram_addr0[5]
  PIN sram_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 165.280 500.000 165.880 ;
    END
  END sram_addr0[6]
  PIN sram_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 182.960 500.000 183.560 ;
    END
  END sram_addr0[7]
  PIN sram_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 200.640 500.000 201.240 ;
    END
  END sram_addr0[8]
  PIN sram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 51.040 500.000 51.640 ;
    END
  END sram_addr1[0]
  PIN sram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 71.440 500.000 72.040 ;
    END
  END sram_addr1[1]
  PIN sram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 91.840 500.000 92.440 ;
    END
  END sram_addr1[2]
  PIN sram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 112.240 500.000 112.840 ;
    END
  END sram_addr1[3]
  PIN sram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 132.640 500.000 133.240 ;
    END
  END sram_addr1[4]
  PIN sram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 150.320 500.000 150.920 ;
    END
  END sram_addr1[5]
  PIN sram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 168.000 500.000 168.600 ;
    END
  END sram_addr1[6]
  PIN sram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 185.680 500.000 186.280 ;
    END
  END sram_addr1[7]
  PIN sram_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 203.360 500.000 203.960 ;
    END
  END sram_addr1[8]
  PIN sram_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 30.640 500.000 31.240 ;
    END
  END sram_clk0
  PIN sram_clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 33.360 500.000 33.960 ;
    END
  END sram_clk1
  PIN sram_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 53.760 500.000 54.360 ;
    END
  END sram_din0[0]
  PIN sram_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 231.240 500.000 231.840 ;
    END
  END sram_din0[10]
  PIN sram_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 244.160 500.000 244.760 ;
    END
  END sram_din0[11]
  PIN sram_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 256.400 500.000 257.000 ;
    END
  END sram_din0[12]
  PIN sram_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 269.320 500.000 269.920 ;
    END
  END sram_din0[13]
  PIN sram_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 282.240 500.000 282.840 ;
    END
  END sram_din0[14]
  PIN sram_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 294.480 500.000 295.080 ;
    END
  END sram_din0[15]
  PIN sram_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 307.400 500.000 308.000 ;
    END
  END sram_din0[16]
  PIN sram_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 320.320 500.000 320.920 ;
    END
  END sram_din0[17]
  PIN sram_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 332.560 500.000 333.160 ;
    END
  END sram_din0[18]
  PIN sram_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 345.480 500.000 346.080 ;
    END
  END sram_din0[19]
  PIN sram_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 74.160 500.000 74.760 ;
    END
  END sram_din0[1]
  PIN sram_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 358.400 500.000 359.000 ;
    END
  END sram_din0[20]
  PIN sram_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 370.640 500.000 371.240 ;
    END
  END sram_din0[21]
  PIN sram_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 383.560 500.000 384.160 ;
    END
  END sram_din0[22]
  PIN sram_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 396.480 500.000 397.080 ;
    END
  END sram_din0[23]
  PIN sram_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 408.720 500.000 409.320 ;
    END
  END sram_din0[24]
  PIN sram_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 421.640 500.000 422.240 ;
    END
  END sram_din0[25]
  PIN sram_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 433.880 500.000 434.480 ;
    END
  END sram_din0[26]
  PIN sram_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 446.800 500.000 447.400 ;
    END
  END sram_din0[27]
  PIN sram_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 459.720 500.000 460.320 ;
    END
  END sram_din0[28]
  PIN sram_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 471.960 500.000 472.560 ;
    END
  END sram_din0[29]
  PIN sram_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 94.560 500.000 95.160 ;
    END
  END sram_din0[2]
  PIN sram_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 484.880 500.000 485.480 ;
    END
  END sram_din0[30]
  PIN sram_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 497.800 500.000 498.400 ;
    END
  END sram_din0[31]
  PIN sram_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 114.280 500.000 114.880 ;
    END
  END sram_din0[3]
  PIN sram_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 134.680 500.000 135.280 ;
    END
  END sram_din0[4]
  PIN sram_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 152.360 500.000 152.960 ;
    END
  END sram_din0[5]
  PIN sram_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 170.040 500.000 170.640 ;
    END
  END sram_din0[6]
  PIN sram_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 188.400 500.000 189.000 ;
    END
  END sram_din0[7]
  PIN sram_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 206.080 500.000 206.680 ;
    END
  END sram_din0[8]
  PIN sram_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 218.320 500.000 218.920 ;
    END
  END sram_din0[9]
  PIN sram_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 36.080 500.000 36.680 ;
    END
  END sram_web0
  PIN sram_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 56.480 500.000 57.080 ;
    END
  END sram_wmask0[0]
  PIN sram_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 76.200 500.000 76.800 ;
    END
  END sram_wmask0[1]
  PIN sram_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 96.600 500.000 97.200 ;
    END
  END sram_wmask0[2]
  PIN sram_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 117.000 500.000 117.600 ;
    END
  END sram_wmask0[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vga_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 5.480 500.000 6.080 ;
    END
  END vga_b[0]
  PIN vga_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 12.960 500.000 13.560 ;
    END
  END vga_b[1]
  PIN vga_g[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 8.200 500.000 8.800 ;
    END
  END vga_g[0]
  PIN vga_g[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 15.680 500.000 16.280 ;
    END
  END vga_g[1]
  PIN vga_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 0.720 500.000 1.320 ;
    END
  END vga_hsync
  PIN vga_r[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 10.240 500.000 10.840 ;
    END
  END vga_r[0]
  PIN vga_r[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 18.400 500.000 19.000 ;
    END
  END vga_r[1]
  PIN vga_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 2.760 500.000 3.360 ;
    END
  END vga_vsync
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END wb_cyc_i
  PIN wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END wb_data_i[0]
  PIN wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END wb_data_i[10]
  PIN wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END wb_data_i[11]
  PIN wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END wb_data_i[12]
  PIN wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END wb_data_i[13]
  PIN wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END wb_data_i[14]
  PIN wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END wb_data_i[15]
  PIN wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END wb_data_i[16]
  PIN wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END wb_data_i[17]
  PIN wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END wb_data_i[18]
  PIN wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END wb_data_i[19]
  PIN wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END wb_data_i[1]
  PIN wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END wb_data_i[20]
  PIN wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END wb_data_i[21]
  PIN wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END wb_data_i[22]
  PIN wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END wb_data_i[23]
  PIN wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END wb_data_i[24]
  PIN wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END wb_data_i[25]
  PIN wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END wb_data_i[26]
  PIN wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END wb_data_i[27]
  PIN wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END wb_data_i[28]
  PIN wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END wb_data_i[29]
  PIN wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wb_data_i[2]
  PIN wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END wb_data_i[30]
  PIN wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END wb_data_i[31]
  PIN wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END wb_data_i[3]
  PIN wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END wb_data_i[4]
  PIN wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END wb_data_i[5]
  PIN wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END wb_data_i[6]
  PIN wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END wb_data_i[7]
  PIN wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END wb_data_i[8]
  PIN wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END wb_data_i[9]
  PIN wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END wb_data_o[0]
  PIN wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END wb_data_o[10]
  PIN wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END wb_data_o[11]
  PIN wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END wb_data_o[12]
  PIN wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END wb_data_o[13]
  PIN wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END wb_data_o[14]
  PIN wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END wb_data_o[15]
  PIN wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END wb_data_o[16]
  PIN wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END wb_data_o[17]
  PIN wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END wb_data_o[18]
  PIN wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END wb_data_o[19]
  PIN wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END wb_data_o[1]
  PIN wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END wb_data_o[20]
  PIN wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END wb_data_o[21]
  PIN wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END wb_data_o[22]
  PIN wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END wb_data_o[23]
  PIN wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 4.000 ;
    END
  END wb_data_o[24]
  PIN wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END wb_data_o[25]
  PIN wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END wb_data_o[26]
  PIN wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END wb_data_o[27]
  PIN wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END wb_data_o[28]
  PIN wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 0.000 477.390 4.000 ;
    END
  END wb_data_o[29]
  PIN wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END wb_data_o[2]
  PIN wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END wb_data_o[30]
  PIN wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END wb_data_o[31]
  PIN wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END wb_data_o[3]
  PIN wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END wb_data_o[4]
  PIN wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END wb_data_o[5]
  PIN wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END wb_data_o[6]
  PIN wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wb_data_o[7]
  PIN wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END wb_data_o[8]
  PIN wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END wb_data_o[9]
  PIN wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END wb_error_o
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END wb_sel_i[3]
  PIN wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END wb_stall_o
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 2.370 6.840 499.950 487.120 ;
      LAYER met2 ;
        RECT 2.400 4.280 499.930 498.285 ;
        RECT 2.950 0.835 6.710 4.280 ;
        RECT 7.550 0.835 11.770 4.280 ;
        RECT 12.610 0.835 16.830 4.280 ;
        RECT 17.670 0.835 21.890 4.280 ;
        RECT 22.730 0.835 26.950 4.280 ;
        RECT 27.790 0.835 32.010 4.280 ;
        RECT 32.850 0.835 37.070 4.280 ;
        RECT 37.910 0.835 41.670 4.280 ;
        RECT 42.510 0.835 46.730 4.280 ;
        RECT 47.570 0.835 51.790 4.280 ;
        RECT 52.630 0.835 56.850 4.280 ;
        RECT 57.690 0.835 61.910 4.280 ;
        RECT 62.750 0.835 66.970 4.280 ;
        RECT 67.810 0.835 72.030 4.280 ;
        RECT 72.870 0.835 77.090 4.280 ;
        RECT 77.930 0.835 81.690 4.280 ;
        RECT 82.530 0.835 86.750 4.280 ;
        RECT 87.590 0.835 91.810 4.280 ;
        RECT 92.650 0.835 96.870 4.280 ;
        RECT 97.710 0.835 101.930 4.280 ;
        RECT 102.770 0.835 106.990 4.280 ;
        RECT 107.830 0.835 112.050 4.280 ;
        RECT 112.890 0.835 117.110 4.280 ;
        RECT 117.950 0.835 121.710 4.280 ;
        RECT 122.550 0.835 126.770 4.280 ;
        RECT 127.610 0.835 131.830 4.280 ;
        RECT 132.670 0.835 136.890 4.280 ;
        RECT 137.730 0.835 141.950 4.280 ;
        RECT 142.790 0.835 147.010 4.280 ;
        RECT 147.850 0.835 152.070 4.280 ;
        RECT 152.910 0.835 156.670 4.280 ;
        RECT 157.510 0.835 161.730 4.280 ;
        RECT 162.570 0.835 166.790 4.280 ;
        RECT 167.630 0.835 171.850 4.280 ;
        RECT 172.690 0.835 176.910 4.280 ;
        RECT 177.750 0.835 181.970 4.280 ;
        RECT 182.810 0.835 187.030 4.280 ;
        RECT 187.870 0.835 192.090 4.280 ;
        RECT 192.930 0.835 196.690 4.280 ;
        RECT 197.530 0.835 201.750 4.280 ;
        RECT 202.590 0.835 206.810 4.280 ;
        RECT 207.650 0.835 211.870 4.280 ;
        RECT 212.710 0.835 216.930 4.280 ;
        RECT 217.770 0.835 221.990 4.280 ;
        RECT 222.830 0.835 227.050 4.280 ;
        RECT 227.890 0.835 232.110 4.280 ;
        RECT 232.950 0.835 236.710 4.280 ;
        RECT 237.550 0.835 241.770 4.280 ;
        RECT 242.610 0.835 246.830 4.280 ;
        RECT 247.670 0.835 251.890 4.280 ;
        RECT 252.730 0.835 256.950 4.280 ;
        RECT 257.790 0.835 262.010 4.280 ;
        RECT 262.850 0.835 267.070 4.280 ;
        RECT 267.910 0.835 271.670 4.280 ;
        RECT 272.510 0.835 276.730 4.280 ;
        RECT 277.570 0.835 281.790 4.280 ;
        RECT 282.630 0.835 286.850 4.280 ;
        RECT 287.690 0.835 291.910 4.280 ;
        RECT 292.750 0.835 296.970 4.280 ;
        RECT 297.810 0.835 302.030 4.280 ;
        RECT 302.870 0.835 307.090 4.280 ;
        RECT 307.930 0.835 311.690 4.280 ;
        RECT 312.530 0.835 316.750 4.280 ;
        RECT 317.590 0.835 321.810 4.280 ;
        RECT 322.650 0.835 326.870 4.280 ;
        RECT 327.710 0.835 331.930 4.280 ;
        RECT 332.770 0.835 336.990 4.280 ;
        RECT 337.830 0.835 342.050 4.280 ;
        RECT 342.890 0.835 347.110 4.280 ;
        RECT 347.950 0.835 351.710 4.280 ;
        RECT 352.550 0.835 356.770 4.280 ;
        RECT 357.610 0.835 361.830 4.280 ;
        RECT 362.670 0.835 366.890 4.280 ;
        RECT 367.730 0.835 371.950 4.280 ;
        RECT 372.790 0.835 377.010 4.280 ;
        RECT 377.850 0.835 382.070 4.280 ;
        RECT 382.910 0.835 386.670 4.280 ;
        RECT 387.510 0.835 391.730 4.280 ;
        RECT 392.570 0.835 396.790 4.280 ;
        RECT 397.630 0.835 401.850 4.280 ;
        RECT 402.690 0.835 406.910 4.280 ;
        RECT 407.750 0.835 411.970 4.280 ;
        RECT 412.810 0.835 417.030 4.280 ;
        RECT 417.870 0.835 422.090 4.280 ;
        RECT 422.930 0.835 426.690 4.280 ;
        RECT 427.530 0.835 431.750 4.280 ;
        RECT 432.590 0.835 436.810 4.280 ;
        RECT 437.650 0.835 441.870 4.280 ;
        RECT 442.710 0.835 446.930 4.280 ;
        RECT 447.770 0.835 451.990 4.280 ;
        RECT 452.830 0.835 457.050 4.280 ;
        RECT 457.890 0.835 462.110 4.280 ;
        RECT 462.950 0.835 466.710 4.280 ;
        RECT 467.550 0.835 471.770 4.280 ;
        RECT 472.610 0.835 476.830 4.280 ;
        RECT 477.670 0.835 481.890 4.280 ;
        RECT 482.730 0.835 486.950 4.280 ;
        RECT 487.790 0.835 492.010 4.280 ;
        RECT 492.850 0.835 497.070 4.280 ;
        RECT 497.910 0.835 499.930 4.280 ;
      LAYER met3 ;
        RECT 9.265 497.400 495.600 498.265 ;
        RECT 9.265 496.080 499.955 497.400 ;
        RECT 9.265 494.680 495.600 496.080 ;
        RECT 9.265 493.360 499.955 494.680 ;
        RECT 9.265 491.960 495.600 493.360 ;
        RECT 9.265 491.320 499.955 491.960 ;
        RECT 9.265 489.920 495.600 491.320 ;
        RECT 9.265 488.600 499.955 489.920 ;
        RECT 9.265 487.200 495.600 488.600 ;
        RECT 9.265 485.880 499.955 487.200 ;
        RECT 9.265 484.480 495.600 485.880 ;
        RECT 9.265 483.160 499.955 484.480 ;
        RECT 9.265 481.760 495.600 483.160 ;
        RECT 9.265 481.120 499.955 481.760 ;
        RECT 9.265 479.720 495.600 481.120 ;
        RECT 9.265 478.400 499.955 479.720 ;
        RECT 9.265 477.000 495.600 478.400 ;
        RECT 9.265 475.680 499.955 477.000 ;
        RECT 9.265 474.280 495.600 475.680 ;
        RECT 9.265 472.960 499.955 474.280 ;
        RECT 9.265 471.560 495.600 472.960 ;
        RECT 9.265 470.920 499.955 471.560 ;
        RECT 9.265 469.520 495.600 470.920 ;
        RECT 9.265 468.200 499.955 469.520 ;
        RECT 9.265 466.800 495.600 468.200 ;
        RECT 9.265 465.480 499.955 466.800 ;
        RECT 9.265 464.080 495.600 465.480 ;
        RECT 9.265 463.440 499.955 464.080 ;
        RECT 9.265 462.040 495.600 463.440 ;
        RECT 9.265 460.720 499.955 462.040 ;
        RECT 9.265 459.320 495.600 460.720 ;
        RECT 9.265 458.000 499.955 459.320 ;
        RECT 9.265 456.600 495.600 458.000 ;
        RECT 9.265 455.280 499.955 456.600 ;
        RECT 9.265 453.880 495.600 455.280 ;
        RECT 9.265 453.240 499.955 453.880 ;
        RECT 9.265 451.840 495.600 453.240 ;
        RECT 9.265 450.520 499.955 451.840 ;
        RECT 9.265 449.120 495.600 450.520 ;
        RECT 9.265 447.800 499.955 449.120 ;
        RECT 9.265 446.400 495.600 447.800 ;
        RECT 9.265 445.080 499.955 446.400 ;
        RECT 9.265 443.680 495.600 445.080 ;
        RECT 9.265 443.040 499.955 443.680 ;
        RECT 9.265 441.640 495.600 443.040 ;
        RECT 9.265 440.320 499.955 441.640 ;
        RECT 9.265 438.920 495.600 440.320 ;
        RECT 9.265 437.600 499.955 438.920 ;
        RECT 9.265 436.200 495.600 437.600 ;
        RECT 9.265 434.880 499.955 436.200 ;
        RECT 9.265 433.480 495.600 434.880 ;
        RECT 9.265 432.840 499.955 433.480 ;
        RECT 9.265 431.440 495.600 432.840 ;
        RECT 9.265 430.120 499.955 431.440 ;
        RECT 9.265 428.720 495.600 430.120 ;
        RECT 9.265 427.400 499.955 428.720 ;
        RECT 9.265 426.000 495.600 427.400 ;
        RECT 9.265 425.360 499.955 426.000 ;
        RECT 9.265 423.960 495.600 425.360 ;
        RECT 9.265 422.640 499.955 423.960 ;
        RECT 9.265 421.240 495.600 422.640 ;
        RECT 9.265 419.920 499.955 421.240 ;
        RECT 9.265 418.520 495.600 419.920 ;
        RECT 9.265 417.200 499.955 418.520 ;
        RECT 9.265 415.800 495.600 417.200 ;
        RECT 9.265 415.160 499.955 415.800 ;
        RECT 9.265 413.760 495.600 415.160 ;
        RECT 9.265 412.440 499.955 413.760 ;
        RECT 9.265 411.040 495.600 412.440 ;
        RECT 9.265 409.720 499.955 411.040 ;
        RECT 9.265 408.320 495.600 409.720 ;
        RECT 9.265 407.000 499.955 408.320 ;
        RECT 9.265 405.600 495.600 407.000 ;
        RECT 9.265 404.960 499.955 405.600 ;
        RECT 9.265 403.560 495.600 404.960 ;
        RECT 9.265 402.240 499.955 403.560 ;
        RECT 9.265 400.840 495.600 402.240 ;
        RECT 9.265 399.520 499.955 400.840 ;
        RECT 9.265 398.120 495.600 399.520 ;
        RECT 9.265 397.480 499.955 398.120 ;
        RECT 9.265 396.080 495.600 397.480 ;
        RECT 9.265 394.760 499.955 396.080 ;
        RECT 9.265 393.360 495.600 394.760 ;
        RECT 9.265 392.040 499.955 393.360 ;
        RECT 9.265 390.640 495.600 392.040 ;
        RECT 9.265 389.320 499.955 390.640 ;
        RECT 9.265 387.920 495.600 389.320 ;
        RECT 9.265 387.280 499.955 387.920 ;
        RECT 9.265 385.880 495.600 387.280 ;
        RECT 9.265 384.560 499.955 385.880 ;
        RECT 9.265 383.160 495.600 384.560 ;
        RECT 9.265 381.840 499.955 383.160 ;
        RECT 9.265 380.440 495.600 381.840 ;
        RECT 9.265 379.120 499.955 380.440 ;
        RECT 9.265 377.720 495.600 379.120 ;
        RECT 9.265 377.080 499.955 377.720 ;
        RECT 9.265 375.680 495.600 377.080 ;
        RECT 9.265 374.360 499.955 375.680 ;
        RECT 9.265 372.960 495.600 374.360 ;
        RECT 9.265 371.640 499.955 372.960 ;
        RECT 9.265 370.240 495.600 371.640 ;
        RECT 9.265 368.920 499.955 370.240 ;
        RECT 9.265 367.520 495.600 368.920 ;
        RECT 9.265 366.880 499.955 367.520 ;
        RECT 9.265 365.480 495.600 366.880 ;
        RECT 9.265 364.160 499.955 365.480 ;
        RECT 9.265 362.760 495.600 364.160 ;
        RECT 9.265 361.440 499.955 362.760 ;
        RECT 9.265 360.040 495.600 361.440 ;
        RECT 9.265 359.400 499.955 360.040 ;
        RECT 9.265 358.000 495.600 359.400 ;
        RECT 9.265 356.680 499.955 358.000 ;
        RECT 9.265 355.280 495.600 356.680 ;
        RECT 9.265 353.960 499.955 355.280 ;
        RECT 9.265 352.560 495.600 353.960 ;
        RECT 9.265 351.240 499.955 352.560 ;
        RECT 9.265 349.840 495.600 351.240 ;
        RECT 9.265 349.200 499.955 349.840 ;
        RECT 9.265 347.800 495.600 349.200 ;
        RECT 9.265 346.480 499.955 347.800 ;
        RECT 9.265 345.080 495.600 346.480 ;
        RECT 9.265 343.760 499.955 345.080 ;
        RECT 9.265 342.360 495.600 343.760 ;
        RECT 9.265 341.040 499.955 342.360 ;
        RECT 9.265 339.640 495.600 341.040 ;
        RECT 9.265 339.000 499.955 339.640 ;
        RECT 9.265 337.600 495.600 339.000 ;
        RECT 9.265 336.280 499.955 337.600 ;
        RECT 9.265 334.880 495.600 336.280 ;
        RECT 9.265 333.560 499.955 334.880 ;
        RECT 9.265 332.160 495.600 333.560 ;
        RECT 9.265 331.520 499.955 332.160 ;
        RECT 9.265 330.120 495.600 331.520 ;
        RECT 9.265 328.800 499.955 330.120 ;
        RECT 9.265 327.400 495.600 328.800 ;
        RECT 9.265 326.080 499.955 327.400 ;
        RECT 9.265 324.680 495.600 326.080 ;
        RECT 9.265 323.360 499.955 324.680 ;
        RECT 9.265 321.960 495.600 323.360 ;
        RECT 9.265 321.320 499.955 321.960 ;
        RECT 9.265 319.920 495.600 321.320 ;
        RECT 9.265 318.600 499.955 319.920 ;
        RECT 9.265 317.200 495.600 318.600 ;
        RECT 9.265 315.880 499.955 317.200 ;
        RECT 9.265 314.480 495.600 315.880 ;
        RECT 9.265 313.160 499.955 314.480 ;
        RECT 9.265 311.760 495.600 313.160 ;
        RECT 9.265 311.120 499.955 311.760 ;
        RECT 9.265 309.720 495.600 311.120 ;
        RECT 9.265 308.400 499.955 309.720 ;
        RECT 9.265 307.000 495.600 308.400 ;
        RECT 9.265 305.680 499.955 307.000 ;
        RECT 9.265 304.280 495.600 305.680 ;
        RECT 9.265 302.960 499.955 304.280 ;
        RECT 9.265 301.560 495.600 302.960 ;
        RECT 9.265 300.920 499.955 301.560 ;
        RECT 9.265 299.520 495.600 300.920 ;
        RECT 9.265 298.200 499.955 299.520 ;
        RECT 9.265 296.800 495.600 298.200 ;
        RECT 9.265 295.480 499.955 296.800 ;
        RECT 9.265 294.080 495.600 295.480 ;
        RECT 9.265 293.440 499.955 294.080 ;
        RECT 9.265 292.040 495.600 293.440 ;
        RECT 9.265 290.720 499.955 292.040 ;
        RECT 9.265 289.320 495.600 290.720 ;
        RECT 9.265 288.000 499.955 289.320 ;
        RECT 9.265 286.600 495.600 288.000 ;
        RECT 9.265 285.280 499.955 286.600 ;
        RECT 9.265 283.880 495.600 285.280 ;
        RECT 9.265 283.240 499.955 283.880 ;
        RECT 9.265 281.840 495.600 283.240 ;
        RECT 9.265 280.520 499.955 281.840 ;
        RECT 9.265 279.120 495.600 280.520 ;
        RECT 9.265 277.800 499.955 279.120 ;
        RECT 9.265 276.400 495.600 277.800 ;
        RECT 9.265 275.080 499.955 276.400 ;
        RECT 9.265 273.680 495.600 275.080 ;
        RECT 9.265 273.040 499.955 273.680 ;
        RECT 9.265 271.640 495.600 273.040 ;
        RECT 9.265 270.320 499.955 271.640 ;
        RECT 9.265 268.920 495.600 270.320 ;
        RECT 9.265 267.600 499.955 268.920 ;
        RECT 9.265 266.200 495.600 267.600 ;
        RECT 9.265 265.560 499.955 266.200 ;
        RECT 9.265 264.160 495.600 265.560 ;
        RECT 9.265 262.840 499.955 264.160 ;
        RECT 9.265 261.440 495.600 262.840 ;
        RECT 9.265 260.120 499.955 261.440 ;
        RECT 9.265 258.720 495.600 260.120 ;
        RECT 9.265 257.400 499.955 258.720 ;
        RECT 9.265 256.000 495.600 257.400 ;
        RECT 9.265 255.360 499.955 256.000 ;
        RECT 9.265 253.960 495.600 255.360 ;
        RECT 9.265 252.640 499.955 253.960 ;
        RECT 9.265 251.240 495.600 252.640 ;
        RECT 9.265 249.920 499.955 251.240 ;
        RECT 9.265 248.520 495.600 249.920 ;
        RECT 9.265 247.200 499.955 248.520 ;
        RECT 9.265 245.800 495.600 247.200 ;
        RECT 9.265 245.160 499.955 245.800 ;
        RECT 9.265 243.760 495.600 245.160 ;
        RECT 9.265 242.440 499.955 243.760 ;
        RECT 9.265 241.040 495.600 242.440 ;
        RECT 9.265 239.720 499.955 241.040 ;
        RECT 9.265 238.320 495.600 239.720 ;
        RECT 9.265 237.000 499.955 238.320 ;
        RECT 9.265 235.600 495.600 237.000 ;
        RECT 9.265 234.960 499.955 235.600 ;
        RECT 9.265 233.560 495.600 234.960 ;
        RECT 9.265 232.240 499.955 233.560 ;
        RECT 9.265 230.840 495.600 232.240 ;
        RECT 9.265 229.520 499.955 230.840 ;
        RECT 9.265 228.120 495.600 229.520 ;
        RECT 9.265 227.480 499.955 228.120 ;
        RECT 9.265 226.080 495.600 227.480 ;
        RECT 9.265 224.760 499.955 226.080 ;
        RECT 9.265 223.360 495.600 224.760 ;
        RECT 9.265 222.040 499.955 223.360 ;
        RECT 9.265 220.640 495.600 222.040 ;
        RECT 9.265 219.320 499.955 220.640 ;
        RECT 9.265 217.920 495.600 219.320 ;
        RECT 9.265 217.280 499.955 217.920 ;
        RECT 9.265 215.880 495.600 217.280 ;
        RECT 9.265 214.560 499.955 215.880 ;
        RECT 9.265 213.160 495.600 214.560 ;
        RECT 9.265 211.840 499.955 213.160 ;
        RECT 9.265 210.440 495.600 211.840 ;
        RECT 9.265 209.120 499.955 210.440 ;
        RECT 9.265 207.720 495.600 209.120 ;
        RECT 9.265 207.080 499.955 207.720 ;
        RECT 9.265 205.680 495.600 207.080 ;
        RECT 9.265 204.360 499.955 205.680 ;
        RECT 9.265 202.960 495.600 204.360 ;
        RECT 9.265 201.640 499.955 202.960 ;
        RECT 9.265 200.240 495.600 201.640 ;
        RECT 9.265 199.600 499.955 200.240 ;
        RECT 9.265 198.200 495.600 199.600 ;
        RECT 9.265 196.880 499.955 198.200 ;
        RECT 9.265 195.480 495.600 196.880 ;
        RECT 9.265 194.160 499.955 195.480 ;
        RECT 9.265 192.760 495.600 194.160 ;
        RECT 9.265 191.440 499.955 192.760 ;
        RECT 9.265 190.040 495.600 191.440 ;
        RECT 9.265 189.400 499.955 190.040 ;
        RECT 9.265 188.000 495.600 189.400 ;
        RECT 9.265 186.680 499.955 188.000 ;
        RECT 9.265 185.280 495.600 186.680 ;
        RECT 9.265 183.960 499.955 185.280 ;
        RECT 9.265 182.560 495.600 183.960 ;
        RECT 9.265 181.240 499.955 182.560 ;
        RECT 9.265 179.840 495.600 181.240 ;
        RECT 9.265 179.200 499.955 179.840 ;
        RECT 9.265 177.800 495.600 179.200 ;
        RECT 9.265 176.480 499.955 177.800 ;
        RECT 9.265 175.080 495.600 176.480 ;
        RECT 9.265 173.760 499.955 175.080 ;
        RECT 9.265 172.360 495.600 173.760 ;
        RECT 9.265 171.040 499.955 172.360 ;
        RECT 9.265 169.640 495.600 171.040 ;
        RECT 9.265 169.000 499.955 169.640 ;
        RECT 9.265 167.600 495.600 169.000 ;
        RECT 9.265 166.280 499.955 167.600 ;
        RECT 9.265 164.880 495.600 166.280 ;
        RECT 9.265 163.560 499.955 164.880 ;
        RECT 9.265 162.160 495.600 163.560 ;
        RECT 9.265 161.520 499.955 162.160 ;
        RECT 9.265 160.120 495.600 161.520 ;
        RECT 9.265 158.800 499.955 160.120 ;
        RECT 9.265 157.400 495.600 158.800 ;
        RECT 9.265 156.080 499.955 157.400 ;
        RECT 9.265 154.680 495.600 156.080 ;
        RECT 9.265 153.360 499.955 154.680 ;
        RECT 9.265 151.960 495.600 153.360 ;
        RECT 9.265 151.320 499.955 151.960 ;
        RECT 9.265 149.920 495.600 151.320 ;
        RECT 9.265 148.600 499.955 149.920 ;
        RECT 9.265 147.200 495.600 148.600 ;
        RECT 9.265 145.880 499.955 147.200 ;
        RECT 9.265 144.480 495.600 145.880 ;
        RECT 9.265 143.160 499.955 144.480 ;
        RECT 9.265 141.760 495.600 143.160 ;
        RECT 9.265 141.120 499.955 141.760 ;
        RECT 9.265 139.720 495.600 141.120 ;
        RECT 9.265 138.400 499.955 139.720 ;
        RECT 9.265 137.000 495.600 138.400 ;
        RECT 9.265 135.680 499.955 137.000 ;
        RECT 9.265 134.280 495.600 135.680 ;
        RECT 9.265 133.640 499.955 134.280 ;
        RECT 9.265 132.240 495.600 133.640 ;
        RECT 9.265 130.920 499.955 132.240 ;
        RECT 9.265 129.520 495.600 130.920 ;
        RECT 9.265 128.200 499.955 129.520 ;
        RECT 9.265 126.800 495.600 128.200 ;
        RECT 9.265 125.480 499.955 126.800 ;
        RECT 9.265 124.080 495.600 125.480 ;
        RECT 9.265 123.440 499.955 124.080 ;
        RECT 9.265 122.040 495.600 123.440 ;
        RECT 9.265 120.720 499.955 122.040 ;
        RECT 9.265 119.320 495.600 120.720 ;
        RECT 9.265 118.000 499.955 119.320 ;
        RECT 9.265 116.600 495.600 118.000 ;
        RECT 9.265 115.280 499.955 116.600 ;
        RECT 9.265 113.880 495.600 115.280 ;
        RECT 9.265 113.240 499.955 113.880 ;
        RECT 9.265 111.840 495.600 113.240 ;
        RECT 9.265 110.520 499.955 111.840 ;
        RECT 9.265 109.120 495.600 110.520 ;
        RECT 9.265 107.800 499.955 109.120 ;
        RECT 9.265 106.400 495.600 107.800 ;
        RECT 9.265 105.080 499.955 106.400 ;
        RECT 9.265 103.680 495.600 105.080 ;
        RECT 9.265 103.040 499.955 103.680 ;
        RECT 9.265 101.640 495.600 103.040 ;
        RECT 9.265 100.320 499.955 101.640 ;
        RECT 9.265 98.920 495.600 100.320 ;
        RECT 9.265 97.600 499.955 98.920 ;
        RECT 9.265 96.200 495.600 97.600 ;
        RECT 9.265 95.560 499.955 96.200 ;
        RECT 9.265 94.160 495.600 95.560 ;
        RECT 9.265 92.840 499.955 94.160 ;
        RECT 9.265 91.440 495.600 92.840 ;
        RECT 9.265 90.120 499.955 91.440 ;
        RECT 9.265 88.720 495.600 90.120 ;
        RECT 9.265 87.400 499.955 88.720 ;
        RECT 9.265 86.000 495.600 87.400 ;
        RECT 9.265 85.360 499.955 86.000 ;
        RECT 9.265 83.960 495.600 85.360 ;
        RECT 9.265 82.640 499.955 83.960 ;
        RECT 9.265 81.240 495.600 82.640 ;
        RECT 9.265 79.920 499.955 81.240 ;
        RECT 9.265 78.520 495.600 79.920 ;
        RECT 9.265 77.200 499.955 78.520 ;
        RECT 9.265 75.800 495.600 77.200 ;
        RECT 9.265 75.160 499.955 75.800 ;
        RECT 9.265 73.760 495.600 75.160 ;
        RECT 9.265 72.440 499.955 73.760 ;
        RECT 9.265 71.040 495.600 72.440 ;
        RECT 9.265 69.720 499.955 71.040 ;
        RECT 9.265 68.320 495.600 69.720 ;
        RECT 9.265 67.680 499.955 68.320 ;
        RECT 9.265 66.280 495.600 67.680 ;
        RECT 9.265 64.960 499.955 66.280 ;
        RECT 9.265 63.560 495.600 64.960 ;
        RECT 9.265 62.240 499.955 63.560 ;
        RECT 9.265 60.840 495.600 62.240 ;
        RECT 9.265 59.520 499.955 60.840 ;
        RECT 9.265 58.120 495.600 59.520 ;
        RECT 9.265 57.480 499.955 58.120 ;
        RECT 9.265 56.080 495.600 57.480 ;
        RECT 9.265 54.760 499.955 56.080 ;
        RECT 9.265 53.360 495.600 54.760 ;
        RECT 9.265 52.040 499.955 53.360 ;
        RECT 9.265 50.640 495.600 52.040 ;
        RECT 9.265 49.320 499.955 50.640 ;
        RECT 9.265 47.920 495.600 49.320 ;
        RECT 9.265 47.280 499.955 47.920 ;
        RECT 9.265 45.880 495.600 47.280 ;
        RECT 9.265 44.560 499.955 45.880 ;
        RECT 9.265 43.160 495.600 44.560 ;
        RECT 9.265 41.840 499.955 43.160 ;
        RECT 9.265 40.440 495.600 41.840 ;
        RECT 9.265 39.120 499.955 40.440 ;
        RECT 9.265 37.720 495.600 39.120 ;
        RECT 9.265 37.080 499.955 37.720 ;
        RECT 9.265 35.680 495.600 37.080 ;
        RECT 9.265 34.360 499.955 35.680 ;
        RECT 9.265 32.960 495.600 34.360 ;
        RECT 9.265 31.640 499.955 32.960 ;
        RECT 9.265 30.240 495.600 31.640 ;
        RECT 9.265 29.600 499.955 30.240 ;
        RECT 9.265 28.200 495.600 29.600 ;
        RECT 9.265 26.880 499.955 28.200 ;
        RECT 9.265 25.480 495.600 26.880 ;
        RECT 9.265 24.160 499.955 25.480 ;
        RECT 9.265 22.760 495.600 24.160 ;
        RECT 9.265 21.440 499.955 22.760 ;
        RECT 9.265 20.040 495.600 21.440 ;
        RECT 9.265 19.400 499.955 20.040 ;
        RECT 9.265 18.000 495.600 19.400 ;
        RECT 9.265 16.680 499.955 18.000 ;
        RECT 9.265 15.280 495.600 16.680 ;
        RECT 9.265 13.960 499.955 15.280 ;
        RECT 9.265 12.560 495.600 13.960 ;
        RECT 9.265 11.240 499.955 12.560 ;
        RECT 9.265 9.840 495.600 11.240 ;
        RECT 9.265 9.200 499.955 9.840 ;
        RECT 9.265 7.800 495.600 9.200 ;
        RECT 9.265 6.480 499.955 7.800 ;
        RECT 9.265 5.080 495.600 6.480 ;
        RECT 9.265 3.760 499.955 5.080 ;
        RECT 9.265 2.360 495.600 3.760 ;
        RECT 9.265 1.720 499.955 2.360 ;
        RECT 9.265 0.855 495.600 1.720 ;
      LAYER met4 ;
        RECT 454.775 17.855 481.440 379.265 ;
        RECT 483.840 17.855 495.585 379.265 ;
  END
END Video
END LIBRARY

