VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Configuration
  CLASS BLOCK ;
  FOREIGN Configuration ;
  ORIGIN 0.000 0.000 ;
  SIZE 50.000 BY 125.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END clk
  PIN core0Index[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 0.720 50.000 1.320 ;
    END
  END core0Index[0]
  PIN core0Index[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 2.760 50.000 3.360 ;
    END
  END core0Index[1]
  PIN core0Index[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 5.480 50.000 6.080 ;
    END
  END core0Index[2]
  PIN core0Index[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 8.200 50.000 8.800 ;
    END
  END core0Index[3]
  PIN core0Index[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 10.920 50.000 11.520 ;
    END
  END core0Index[4]
  PIN core0Index[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 13.640 50.000 14.240 ;
    END
  END core0Index[5]
  PIN core0Index[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 16.360 50.000 16.960 ;
    END
  END core0Index[6]
  PIN core0Index[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 19.080 50.000 19.680 ;
    END
  END core0Index[7]
  PIN core1Index[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 21.800 50.000 22.400 ;
    END
  END core1Index[0]
  PIN core1Index[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 24.520 50.000 25.120 ;
    END
  END core1Index[1]
  PIN core1Index[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 27.240 50.000 27.840 ;
    END
  END core1Index[2]
  PIN core1Index[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 29.960 50.000 30.560 ;
    END
  END core1Index[3]
  PIN core1Index[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 32.000 50.000 32.600 ;
    END
  END core1Index[4]
  PIN core1Index[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 34.720 50.000 35.320 ;
    END
  END core1Index[5]
  PIN core1Index[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 37.440 50.000 38.040 ;
    END
  END core1Index[6]
  PIN core1Index[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 40.160 50.000 40.760 ;
    END
  END core1Index[7]
  PIN manufacturerID[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 42.880 50.000 43.480 ;
    END
  END manufacturerID[0]
  PIN manufacturerID[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 69.400 50.000 70.000 ;
    END
  END manufacturerID[10]
  PIN manufacturerID[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 45.600 50.000 46.200 ;
    END
  END manufacturerID[1]
  PIN manufacturerID[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 48.320 50.000 48.920 ;
    END
  END manufacturerID[2]
  PIN manufacturerID[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 51.040 50.000 51.640 ;
    END
  END manufacturerID[3]
  PIN manufacturerID[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 53.760 50.000 54.360 ;
    END
  END manufacturerID[4]
  PIN manufacturerID[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 56.480 50.000 57.080 ;
    END
  END manufacturerID[5]
  PIN manufacturerID[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 59.200 50.000 59.800 ;
    END
  END manufacturerID[6]
  PIN manufacturerID[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 61.920 50.000 62.520 ;
    END
  END manufacturerID[7]
  PIN manufacturerID[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 63.960 50.000 64.560 ;
    END
  END manufacturerID[8]
  PIN manufacturerID[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 66.680 50.000 67.280 ;
    END
  END manufacturerID[9]
  PIN partID[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 72.120 50.000 72.720 ;
    END
  END partID[0]
  PIN partID[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 98.640 50.000 99.240 ;
    END
  END partID[10]
  PIN partID[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 101.360 50.000 101.960 ;
    END
  END partID[11]
  PIN partID[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 104.080 50.000 104.680 ;
    END
  END partID[12]
  PIN partID[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 106.800 50.000 107.400 ;
    END
  END partID[13]
  PIN partID[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 109.520 50.000 110.120 ;
    END
  END partID[14]
  PIN partID[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 112.240 50.000 112.840 ;
    END
  END partID[15]
  PIN partID[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 74.840 50.000 75.440 ;
    END
  END partID[1]
  PIN partID[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 77.560 50.000 78.160 ;
    END
  END partID[2]
  PIN partID[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 80.280 50.000 80.880 ;
    END
  END partID[3]
  PIN partID[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 83.000 50.000 83.600 ;
    END
  END partID[4]
  PIN partID[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 85.720 50.000 86.320 ;
    END
  END partID[5]
  PIN partID[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 88.440 50.000 89.040 ;
    END
  END partID[6]
  PIN partID[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 91.160 50.000 91.760 ;
    END
  END partID[7]
  PIN partID[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 93.880 50.000 94.480 ;
    END
  END partID[8]
  PIN partID[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 95.920 50.000 96.520 ;
    END
  END partID[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 11.210 10.640 12.810 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.200 10.640 25.800 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.185 10.640 38.785 111.760 ;
    END
  END vccd1
  PIN versionID[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 114.960 50.000 115.560 ;
    END
  END versionID[0]
  PIN versionID[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 117.680 50.000 118.280 ;
    END
  END versionID[1]
  PIN versionID[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 120.400 50.000 121.000 ;
    END
  END versionID[2]
  PIN versionID[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 123.120 50.000 123.720 ;
    END
  END versionID[3]
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 17.710 10.640 19.310 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 30.695 10.640 32.295 111.760 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 110.105 44.350 111.710 ;
        RECT 5.330 104.665 44.350 107.495 ;
        RECT 5.330 99.225 44.350 102.055 ;
        RECT 5.330 93.785 44.350 96.615 ;
        RECT 5.330 88.345 44.350 91.175 ;
        RECT 5.330 82.905 44.350 85.735 ;
        RECT 5.330 77.465 44.350 80.295 ;
        RECT 5.330 72.025 44.350 74.855 ;
        RECT 5.330 66.585 44.350 69.415 ;
        RECT 5.330 61.145 44.350 63.975 ;
        RECT 5.330 55.705 44.350 58.535 ;
        RECT 5.330 50.265 44.350 53.095 ;
        RECT 5.330 44.825 44.350 47.655 ;
        RECT 5.330 39.385 44.350 42.215 ;
        RECT 5.330 33.945 44.350 36.775 ;
        RECT 5.330 28.505 44.350 31.335 ;
        RECT 5.330 23.065 44.350 25.895 ;
        RECT 5.330 17.625 44.350 20.455 ;
        RECT 5.330 12.185 44.350 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 44.160 111.605 ;
      LAYER met1 ;
        RECT 5.520 10.640 44.160 111.760 ;
      LAYER met2 ;
        RECT 11.240 4.280 41.310 123.605 ;
        RECT 11.240 0.835 24.650 4.280 ;
        RECT 25.490 0.835 41.310 4.280 ;
      LAYER met3 ;
        RECT 11.210 122.720 45.600 123.585 ;
        RECT 11.210 121.400 46.000 122.720 ;
        RECT 11.210 120.000 45.600 121.400 ;
        RECT 11.210 118.680 46.000 120.000 ;
        RECT 11.210 117.280 45.600 118.680 ;
        RECT 11.210 115.960 46.000 117.280 ;
        RECT 11.210 114.560 45.600 115.960 ;
        RECT 11.210 113.240 46.000 114.560 ;
        RECT 11.210 111.840 45.600 113.240 ;
        RECT 11.210 110.520 46.000 111.840 ;
        RECT 11.210 109.120 45.600 110.520 ;
        RECT 11.210 107.800 46.000 109.120 ;
        RECT 11.210 106.400 45.600 107.800 ;
        RECT 11.210 105.080 46.000 106.400 ;
        RECT 11.210 103.680 45.600 105.080 ;
        RECT 11.210 102.360 46.000 103.680 ;
        RECT 11.210 100.960 45.600 102.360 ;
        RECT 11.210 99.640 46.000 100.960 ;
        RECT 11.210 98.240 45.600 99.640 ;
        RECT 11.210 96.920 46.000 98.240 ;
        RECT 11.210 95.520 45.600 96.920 ;
        RECT 11.210 94.880 46.000 95.520 ;
        RECT 11.210 93.480 45.600 94.880 ;
        RECT 11.210 92.160 46.000 93.480 ;
        RECT 11.210 90.760 45.600 92.160 ;
        RECT 11.210 89.440 46.000 90.760 ;
        RECT 11.210 88.040 45.600 89.440 ;
        RECT 11.210 86.720 46.000 88.040 ;
        RECT 11.210 85.320 45.600 86.720 ;
        RECT 11.210 84.000 46.000 85.320 ;
        RECT 11.210 82.600 45.600 84.000 ;
        RECT 11.210 81.280 46.000 82.600 ;
        RECT 11.210 79.880 45.600 81.280 ;
        RECT 11.210 78.560 46.000 79.880 ;
        RECT 11.210 77.160 45.600 78.560 ;
        RECT 11.210 75.840 46.000 77.160 ;
        RECT 11.210 74.440 45.600 75.840 ;
        RECT 11.210 73.120 46.000 74.440 ;
        RECT 11.210 71.720 45.600 73.120 ;
        RECT 11.210 70.400 46.000 71.720 ;
        RECT 11.210 69.000 45.600 70.400 ;
        RECT 11.210 67.680 46.000 69.000 ;
        RECT 11.210 66.280 45.600 67.680 ;
        RECT 11.210 64.960 46.000 66.280 ;
        RECT 11.210 63.560 45.600 64.960 ;
        RECT 11.210 62.920 46.000 63.560 ;
        RECT 11.210 61.520 45.600 62.920 ;
        RECT 11.210 60.200 46.000 61.520 ;
        RECT 11.210 58.800 45.600 60.200 ;
        RECT 11.210 57.480 46.000 58.800 ;
        RECT 11.210 56.080 45.600 57.480 ;
        RECT 11.210 54.760 46.000 56.080 ;
        RECT 11.210 53.360 45.600 54.760 ;
        RECT 11.210 52.040 46.000 53.360 ;
        RECT 11.210 50.640 45.600 52.040 ;
        RECT 11.210 49.320 46.000 50.640 ;
        RECT 11.210 47.920 45.600 49.320 ;
        RECT 11.210 46.600 46.000 47.920 ;
        RECT 11.210 45.200 45.600 46.600 ;
        RECT 11.210 43.880 46.000 45.200 ;
        RECT 11.210 42.480 45.600 43.880 ;
        RECT 11.210 41.160 46.000 42.480 ;
        RECT 11.210 39.760 45.600 41.160 ;
        RECT 11.210 38.440 46.000 39.760 ;
        RECT 11.210 37.040 45.600 38.440 ;
        RECT 11.210 35.720 46.000 37.040 ;
        RECT 11.210 34.320 45.600 35.720 ;
        RECT 11.210 33.000 46.000 34.320 ;
        RECT 11.210 31.600 45.600 33.000 ;
        RECT 11.210 30.960 46.000 31.600 ;
        RECT 11.210 29.560 45.600 30.960 ;
        RECT 11.210 28.240 46.000 29.560 ;
        RECT 11.210 26.840 45.600 28.240 ;
        RECT 11.210 25.520 46.000 26.840 ;
        RECT 11.210 24.120 45.600 25.520 ;
        RECT 11.210 22.800 46.000 24.120 ;
        RECT 11.210 21.400 45.600 22.800 ;
        RECT 11.210 20.080 46.000 21.400 ;
        RECT 11.210 18.680 45.600 20.080 ;
        RECT 11.210 17.360 46.000 18.680 ;
        RECT 11.210 15.960 45.600 17.360 ;
        RECT 11.210 14.640 46.000 15.960 ;
        RECT 11.210 13.240 45.600 14.640 ;
        RECT 11.210 11.920 46.000 13.240 ;
        RECT 11.210 10.520 45.600 11.920 ;
        RECT 11.210 9.200 46.000 10.520 ;
        RECT 11.210 7.800 45.600 9.200 ;
        RECT 11.210 6.480 46.000 7.800 ;
        RECT 11.210 5.080 45.600 6.480 ;
        RECT 11.210 3.760 46.000 5.080 ;
        RECT 11.210 2.360 45.600 3.760 ;
        RECT 11.210 1.720 46.000 2.360 ;
        RECT 11.210 0.855 45.600 1.720 ;
      LAYER met4 ;
        RECT 19.710 10.640 23.800 111.760 ;
        RECT 26.200 10.640 30.295 111.760 ;
  END
END Configuration
END LIBRARY

