magic
tech sky130A
magscale 1 2
timestamp 1653084941
<< obsli1 >>
rect 1104 2159 158884 97393
<< obsm1 >>
rect 382 1300 158884 98048
<< metal2 >>
rect 386 99200 442 100000
rect 1214 99200 1270 100000
rect 2042 99200 2098 100000
rect 2870 99200 2926 100000
rect 3698 99200 3754 100000
rect 4618 99200 4674 100000
rect 5446 99200 5502 100000
rect 6274 99200 6330 100000
rect 7102 99200 7158 100000
rect 7930 99200 7986 100000
rect 8850 99200 8906 100000
rect 9678 99200 9734 100000
rect 10506 99200 10562 100000
rect 11334 99200 11390 100000
rect 12162 99200 12218 100000
rect 13082 99200 13138 100000
rect 13910 99200 13966 100000
rect 14738 99200 14794 100000
rect 15566 99200 15622 100000
rect 16394 99200 16450 100000
rect 17314 99200 17370 100000
rect 18142 99200 18198 100000
rect 18970 99200 19026 100000
rect 19798 99200 19854 100000
rect 20626 99200 20682 100000
rect 21546 99200 21602 100000
rect 22374 99200 22430 100000
rect 23202 99200 23258 100000
rect 24030 99200 24086 100000
rect 24858 99200 24914 100000
rect 25778 99200 25834 100000
rect 26606 99200 26662 100000
rect 27434 99200 27490 100000
rect 28262 99200 28318 100000
rect 29090 99200 29146 100000
rect 30010 99200 30066 100000
rect 30838 99200 30894 100000
rect 31666 99200 31722 100000
rect 32494 99200 32550 100000
rect 33322 99200 33378 100000
rect 34242 99200 34298 100000
rect 35070 99200 35126 100000
rect 35898 99200 35954 100000
rect 36726 99200 36782 100000
rect 37554 99200 37610 100000
rect 38474 99200 38530 100000
rect 39302 99200 39358 100000
rect 40130 99200 40186 100000
rect 40958 99200 41014 100000
rect 41786 99200 41842 100000
rect 42706 99200 42762 100000
rect 43534 99200 43590 100000
rect 44362 99200 44418 100000
rect 45190 99200 45246 100000
rect 46018 99200 46074 100000
rect 46938 99200 46994 100000
rect 47766 99200 47822 100000
rect 48594 99200 48650 100000
rect 49422 99200 49478 100000
rect 50250 99200 50306 100000
rect 51170 99200 51226 100000
rect 51998 99200 52054 100000
rect 52826 99200 52882 100000
rect 53654 99200 53710 100000
rect 54482 99200 54538 100000
rect 55402 99200 55458 100000
rect 56230 99200 56286 100000
rect 57058 99200 57114 100000
rect 57886 99200 57942 100000
rect 58714 99200 58770 100000
rect 59634 99200 59690 100000
rect 60462 99200 60518 100000
rect 61290 99200 61346 100000
rect 62118 99200 62174 100000
rect 62946 99200 63002 100000
rect 63866 99200 63922 100000
rect 64694 99200 64750 100000
rect 65522 99200 65578 100000
rect 66350 99200 66406 100000
rect 67178 99200 67234 100000
rect 68098 99200 68154 100000
rect 68926 99200 68982 100000
rect 69754 99200 69810 100000
rect 70582 99200 70638 100000
rect 71410 99200 71466 100000
rect 72330 99200 72386 100000
rect 73158 99200 73214 100000
rect 73986 99200 74042 100000
rect 74814 99200 74870 100000
rect 75642 99200 75698 100000
rect 76562 99200 76618 100000
rect 77390 99200 77446 100000
rect 78218 99200 78274 100000
rect 79046 99200 79102 100000
rect 79874 99200 79930 100000
rect 80794 99200 80850 100000
rect 81622 99200 81678 100000
rect 82450 99200 82506 100000
rect 83278 99200 83334 100000
rect 84106 99200 84162 100000
rect 85026 99200 85082 100000
rect 85854 99200 85910 100000
rect 86682 99200 86738 100000
rect 87510 99200 87566 100000
rect 88338 99200 88394 100000
rect 89258 99200 89314 100000
rect 90086 99200 90142 100000
rect 90914 99200 90970 100000
rect 91742 99200 91798 100000
rect 92570 99200 92626 100000
rect 93490 99200 93546 100000
rect 94318 99200 94374 100000
rect 95146 99200 95202 100000
rect 95974 99200 96030 100000
rect 96802 99200 96858 100000
rect 97722 99200 97778 100000
rect 98550 99200 98606 100000
rect 99378 99200 99434 100000
rect 100206 99200 100262 100000
rect 101034 99200 101090 100000
rect 101954 99200 102010 100000
rect 102782 99200 102838 100000
rect 103610 99200 103666 100000
rect 104438 99200 104494 100000
rect 105266 99200 105322 100000
rect 106186 99200 106242 100000
rect 107014 99200 107070 100000
rect 107842 99200 107898 100000
rect 108670 99200 108726 100000
rect 109498 99200 109554 100000
rect 110418 99200 110474 100000
rect 111246 99200 111302 100000
rect 112074 99200 112130 100000
rect 112902 99200 112958 100000
rect 113730 99200 113786 100000
rect 114650 99200 114706 100000
rect 115478 99200 115534 100000
rect 116306 99200 116362 100000
rect 117134 99200 117190 100000
rect 117962 99200 118018 100000
rect 118882 99200 118938 100000
rect 119710 99200 119766 100000
rect 120538 99200 120594 100000
rect 121366 99200 121422 100000
rect 122194 99200 122250 100000
rect 123114 99200 123170 100000
rect 123942 99200 123998 100000
rect 124770 99200 124826 100000
rect 125598 99200 125654 100000
rect 126426 99200 126482 100000
rect 127346 99200 127402 100000
rect 128174 99200 128230 100000
rect 129002 99200 129058 100000
rect 129830 99200 129886 100000
rect 130658 99200 130714 100000
rect 131578 99200 131634 100000
rect 132406 99200 132462 100000
rect 133234 99200 133290 100000
rect 134062 99200 134118 100000
rect 134890 99200 134946 100000
rect 135810 99200 135866 100000
rect 136638 99200 136694 100000
rect 137466 99200 137522 100000
rect 138294 99200 138350 100000
rect 139122 99200 139178 100000
rect 140042 99200 140098 100000
rect 140870 99200 140926 100000
rect 141698 99200 141754 100000
rect 142526 99200 142582 100000
rect 143354 99200 143410 100000
rect 144274 99200 144330 100000
rect 145102 99200 145158 100000
rect 145930 99200 145986 100000
rect 146758 99200 146814 100000
rect 147586 99200 147642 100000
rect 148506 99200 148562 100000
rect 149334 99200 149390 100000
rect 150162 99200 150218 100000
rect 150990 99200 151046 100000
rect 151818 99200 151874 100000
rect 152738 99200 152794 100000
rect 153566 99200 153622 100000
rect 154394 99200 154450 100000
rect 155222 99200 155278 100000
rect 156050 99200 156106 100000
rect 156970 99200 157026 100000
rect 157798 99200 157854 100000
rect 158626 99200 158682 100000
rect 159454 99200 159510 100000
rect 2042 0 2098 800
rect 6090 0 6146 800
rect 10230 0 10286 800
rect 14278 0 14334 800
rect 18418 0 18474 800
rect 22466 0 22522 800
rect 26606 0 26662 800
rect 30746 0 30802 800
rect 34794 0 34850 800
rect 38934 0 38990 800
rect 42982 0 43038 800
rect 47122 0 47178 800
rect 51262 0 51318 800
rect 55310 0 55366 800
rect 59450 0 59506 800
rect 63498 0 63554 800
rect 67638 0 67694 800
rect 71778 0 71834 800
rect 75826 0 75882 800
rect 79966 0 80022 800
rect 84014 0 84070 800
rect 88154 0 88210 800
rect 92202 0 92258 800
rect 96342 0 96398 800
rect 100482 0 100538 800
rect 104530 0 104586 800
rect 108670 0 108726 800
rect 112718 0 112774 800
rect 116858 0 116914 800
rect 120998 0 121054 800
rect 125046 0 125102 800
rect 129186 0 129242 800
rect 133234 0 133290 800
rect 137374 0 137430 800
rect 141514 0 141570 800
rect 145562 0 145618 800
rect 149702 0 149758 800
rect 153750 0 153806 800
rect 157890 0 157946 800
<< obsm2 >>
rect 498 99144 1158 99657
rect 1326 99144 1986 99657
rect 2154 99144 2814 99657
rect 2982 99144 3642 99657
rect 3810 99144 4562 99657
rect 4730 99144 5390 99657
rect 5558 99144 6218 99657
rect 6386 99144 7046 99657
rect 7214 99144 7874 99657
rect 8042 99144 8794 99657
rect 8962 99144 9622 99657
rect 9790 99144 10450 99657
rect 10618 99144 11278 99657
rect 11446 99144 12106 99657
rect 12274 99144 13026 99657
rect 13194 99144 13854 99657
rect 14022 99144 14682 99657
rect 14850 99144 15510 99657
rect 15678 99144 16338 99657
rect 16506 99144 17258 99657
rect 17426 99144 18086 99657
rect 18254 99144 18914 99657
rect 19082 99144 19742 99657
rect 19910 99144 20570 99657
rect 20738 99144 21490 99657
rect 21658 99144 22318 99657
rect 22486 99144 23146 99657
rect 23314 99144 23974 99657
rect 24142 99144 24802 99657
rect 24970 99144 25722 99657
rect 25890 99144 26550 99657
rect 26718 99144 27378 99657
rect 27546 99144 28206 99657
rect 28374 99144 29034 99657
rect 29202 99144 29954 99657
rect 30122 99144 30782 99657
rect 30950 99144 31610 99657
rect 31778 99144 32438 99657
rect 32606 99144 33266 99657
rect 33434 99144 34186 99657
rect 34354 99144 35014 99657
rect 35182 99144 35842 99657
rect 36010 99144 36670 99657
rect 36838 99144 37498 99657
rect 37666 99144 38418 99657
rect 38586 99144 39246 99657
rect 39414 99144 40074 99657
rect 40242 99144 40902 99657
rect 41070 99144 41730 99657
rect 41898 99144 42650 99657
rect 42818 99144 43478 99657
rect 43646 99144 44306 99657
rect 44474 99144 45134 99657
rect 45302 99144 45962 99657
rect 46130 99144 46882 99657
rect 47050 99144 47710 99657
rect 47878 99144 48538 99657
rect 48706 99144 49366 99657
rect 49534 99144 50194 99657
rect 50362 99144 51114 99657
rect 51282 99144 51942 99657
rect 52110 99144 52770 99657
rect 52938 99144 53598 99657
rect 53766 99144 54426 99657
rect 54594 99144 55346 99657
rect 55514 99144 56174 99657
rect 56342 99144 57002 99657
rect 57170 99144 57830 99657
rect 57998 99144 58658 99657
rect 58826 99144 59578 99657
rect 59746 99144 60406 99657
rect 60574 99144 61234 99657
rect 61402 99144 62062 99657
rect 62230 99144 62890 99657
rect 63058 99144 63810 99657
rect 63978 99144 64638 99657
rect 64806 99144 65466 99657
rect 65634 99144 66294 99657
rect 66462 99144 67122 99657
rect 67290 99144 68042 99657
rect 68210 99144 68870 99657
rect 69038 99144 69698 99657
rect 69866 99144 70526 99657
rect 70694 99144 71354 99657
rect 71522 99144 72274 99657
rect 72442 99144 73102 99657
rect 73270 99144 73930 99657
rect 74098 99144 74758 99657
rect 74926 99144 75586 99657
rect 75754 99144 76506 99657
rect 76674 99144 77334 99657
rect 77502 99144 78162 99657
rect 78330 99144 78990 99657
rect 79158 99144 79818 99657
rect 79986 99144 80738 99657
rect 80906 99144 81566 99657
rect 81734 99144 82394 99657
rect 82562 99144 83222 99657
rect 83390 99144 84050 99657
rect 84218 99144 84970 99657
rect 85138 99144 85798 99657
rect 85966 99144 86626 99657
rect 86794 99144 87454 99657
rect 87622 99144 88282 99657
rect 88450 99144 89202 99657
rect 89370 99144 90030 99657
rect 90198 99144 90858 99657
rect 91026 99144 91686 99657
rect 91854 99144 92514 99657
rect 92682 99144 93434 99657
rect 93602 99144 94262 99657
rect 94430 99144 95090 99657
rect 95258 99144 95918 99657
rect 96086 99144 96746 99657
rect 96914 99144 97666 99657
rect 97834 99144 98494 99657
rect 98662 99144 99322 99657
rect 99490 99144 100150 99657
rect 100318 99144 100978 99657
rect 101146 99144 101898 99657
rect 102066 99144 102726 99657
rect 102894 99144 103554 99657
rect 103722 99144 104382 99657
rect 104550 99144 105210 99657
rect 105378 99144 106130 99657
rect 106298 99144 106958 99657
rect 107126 99144 107786 99657
rect 107954 99144 108614 99657
rect 108782 99144 109442 99657
rect 109610 99144 110362 99657
rect 110530 99144 111190 99657
rect 111358 99144 112018 99657
rect 112186 99144 112846 99657
rect 113014 99144 113674 99657
rect 113842 99144 114594 99657
rect 114762 99144 115422 99657
rect 115590 99144 116250 99657
rect 116418 99144 117078 99657
rect 117246 99144 117906 99657
rect 118074 99144 118826 99657
rect 118994 99144 119654 99657
rect 119822 99144 120482 99657
rect 120650 99144 121310 99657
rect 121478 99144 122138 99657
rect 122306 99144 123058 99657
rect 123226 99144 123886 99657
rect 124054 99144 124714 99657
rect 124882 99144 125542 99657
rect 125710 99144 126370 99657
rect 126538 99144 127290 99657
rect 127458 99144 128118 99657
rect 128286 99144 128946 99657
rect 129114 99144 129774 99657
rect 129942 99144 130602 99657
rect 130770 99144 131522 99657
rect 131690 99144 132350 99657
rect 132518 99144 133178 99657
rect 133346 99144 134006 99657
rect 134174 99144 134834 99657
rect 135002 99144 135754 99657
rect 135922 99144 136582 99657
rect 136750 99144 137410 99657
rect 137578 99144 138238 99657
rect 138406 99144 139066 99657
rect 139234 99144 139986 99657
rect 140154 99144 140814 99657
rect 140982 99144 141642 99657
rect 141810 99144 142470 99657
rect 142638 99144 143298 99657
rect 143466 99144 144218 99657
rect 144386 99144 145046 99657
rect 145214 99144 145874 99657
rect 146042 99144 146702 99657
rect 146870 99144 147530 99657
rect 147698 99144 148450 99657
rect 148618 99144 149278 99657
rect 149446 99144 150106 99657
rect 150274 99144 150934 99657
rect 151102 99144 151762 99657
rect 151930 99144 152682 99657
rect 152850 99144 153510 99657
rect 153678 99144 154338 99657
rect 154506 99144 155166 99657
rect 155334 99144 155994 99657
rect 156162 99144 156914 99657
rect 157082 99144 157742 99657
rect 157910 99144 158498 99657
rect 388 856 158498 99144
rect 388 167 1986 856
rect 2154 167 6034 856
rect 6202 167 10174 856
rect 10342 167 14222 856
rect 14390 167 18362 856
rect 18530 167 22410 856
rect 22578 167 26550 856
rect 26718 167 30690 856
rect 30858 167 34738 856
rect 34906 167 38878 856
rect 39046 167 42926 856
rect 43094 167 47066 856
rect 47234 167 51206 856
rect 51374 167 55254 856
rect 55422 167 59394 856
rect 59562 167 63442 856
rect 63610 167 67582 856
rect 67750 167 71722 856
rect 71890 167 75770 856
rect 75938 167 79910 856
rect 80078 167 83958 856
rect 84126 167 88098 856
rect 88266 167 92146 856
rect 92314 167 96286 856
rect 96454 167 100426 856
rect 100594 167 104474 856
rect 104642 167 108614 856
rect 108782 167 112662 856
rect 112830 167 116802 856
rect 116970 167 120942 856
rect 121110 167 124990 856
rect 125158 167 129130 856
rect 129298 167 133178 856
rect 133346 167 137318 856
rect 137486 167 141458 856
rect 141626 167 145506 856
rect 145674 167 149646 856
rect 149814 167 153694 856
rect 153862 167 157834 856
rect 158002 167 158498 856
<< metal3 >>
rect 159200 99560 160000 99680
rect 0 99016 800 99136
rect 159200 99016 160000 99136
rect 159200 98608 160000 98728
rect 159200 98064 160000 98184
rect 0 97384 800 97504
rect 159200 97520 160000 97640
rect 159200 97112 160000 97232
rect 159200 96568 160000 96688
rect 159200 96024 160000 96144
rect 0 95616 800 95736
rect 159200 95616 160000 95736
rect 159200 95072 160000 95192
rect 159200 94528 160000 94648
rect 0 93984 800 94104
rect 159200 94120 160000 94240
rect 159200 93576 160000 93696
rect 159200 93168 160000 93288
rect 159200 92624 160000 92744
rect 0 92216 800 92336
rect 159200 92080 160000 92200
rect 159200 91672 160000 91792
rect 159200 91128 160000 91248
rect 0 90584 800 90704
rect 159200 90584 160000 90704
rect 159200 90176 160000 90296
rect 159200 89632 160000 89752
rect 159200 89088 160000 89208
rect 0 88816 800 88936
rect 159200 88680 160000 88800
rect 159200 88136 160000 88256
rect 159200 87728 160000 87848
rect 0 87184 800 87304
rect 159200 87184 160000 87304
rect 159200 86640 160000 86760
rect 159200 86232 160000 86352
rect 159200 85688 160000 85808
rect 0 85416 800 85536
rect 159200 85144 160000 85264
rect 159200 84736 160000 84856
rect 159200 84192 160000 84312
rect 0 83784 800 83904
rect 159200 83648 160000 83768
rect 159200 83240 160000 83360
rect 159200 82696 160000 82816
rect 159200 82288 160000 82408
rect 0 82016 800 82136
rect 159200 81744 160000 81864
rect 159200 81200 160000 81320
rect 159200 80792 160000 80912
rect 0 80384 800 80504
rect 159200 80248 160000 80368
rect 159200 79704 160000 79824
rect 159200 79296 160000 79416
rect 0 78752 800 78872
rect 159200 78752 160000 78872
rect 159200 78208 160000 78328
rect 159200 77800 160000 77920
rect 159200 77256 160000 77376
rect 0 76984 800 77104
rect 159200 76712 160000 76832
rect 159200 76304 160000 76424
rect 159200 75760 160000 75880
rect 0 75352 800 75472
rect 159200 75352 160000 75472
rect 159200 74808 160000 74928
rect 159200 74264 160000 74384
rect 159200 73856 160000 73976
rect 0 73584 800 73704
rect 159200 73312 160000 73432
rect 159200 72768 160000 72888
rect 159200 72360 160000 72480
rect 0 71952 800 72072
rect 159200 71816 160000 71936
rect 159200 71272 160000 71392
rect 159200 70864 160000 70984
rect 0 70184 800 70304
rect 159200 70320 160000 70440
rect 159200 69912 160000 70032
rect 159200 69368 160000 69488
rect 159200 68824 160000 68944
rect 0 68552 800 68672
rect 159200 68416 160000 68536
rect 159200 67872 160000 67992
rect 159200 67328 160000 67448
rect 0 66784 800 66904
rect 159200 66920 160000 67040
rect 159200 66376 160000 66496
rect 159200 65832 160000 65952
rect 159200 65424 160000 65544
rect 0 65152 800 65272
rect 159200 64880 160000 65000
rect 159200 64472 160000 64592
rect 159200 63928 160000 64048
rect 0 63384 800 63504
rect 159200 63384 160000 63504
rect 159200 62976 160000 63096
rect 159200 62432 160000 62552
rect 0 61752 800 61872
rect 159200 61888 160000 62008
rect 159200 61480 160000 61600
rect 159200 60936 160000 61056
rect 159200 60392 160000 60512
rect 0 60120 800 60240
rect 159200 59984 160000 60104
rect 159200 59440 160000 59560
rect 159200 58896 160000 59016
rect 0 58352 800 58472
rect 159200 58488 160000 58608
rect 159200 57944 160000 58064
rect 159200 57536 160000 57656
rect 159200 56992 160000 57112
rect 0 56720 800 56840
rect 159200 56448 160000 56568
rect 159200 56040 160000 56160
rect 159200 55496 160000 55616
rect 0 54952 800 55072
rect 159200 54952 160000 55072
rect 159200 54544 160000 54664
rect 159200 54000 160000 54120
rect 0 53320 800 53440
rect 159200 53456 160000 53576
rect 159200 53048 160000 53168
rect 159200 52504 160000 52624
rect 159200 52096 160000 52216
rect 0 51552 800 51672
rect 159200 51552 160000 51672
rect 159200 51008 160000 51128
rect 159200 50600 160000 50720
rect 0 49920 800 50040
rect 159200 50056 160000 50176
rect 159200 49512 160000 49632
rect 159200 49104 160000 49224
rect 159200 48560 160000 48680
rect 0 48152 800 48272
rect 159200 48016 160000 48136
rect 159200 47608 160000 47728
rect 159200 47064 160000 47184
rect 0 46520 800 46640
rect 159200 46656 160000 46776
rect 159200 46112 160000 46232
rect 159200 45568 160000 45688
rect 159200 45160 160000 45280
rect 0 44752 800 44872
rect 159200 44616 160000 44736
rect 159200 44072 160000 44192
rect 159200 43664 160000 43784
rect 0 43120 800 43240
rect 159200 43120 160000 43240
rect 159200 42576 160000 42696
rect 159200 42168 160000 42288
rect 159200 41624 160000 41744
rect 0 41352 800 41472
rect 159200 41216 160000 41336
rect 159200 40672 160000 40792
rect 159200 40128 160000 40248
rect 0 39720 800 39840
rect 159200 39720 160000 39840
rect 159200 39176 160000 39296
rect 159200 38632 160000 38752
rect 0 38088 800 38208
rect 159200 38224 160000 38344
rect 159200 37680 160000 37800
rect 159200 37136 160000 37256
rect 159200 36728 160000 36848
rect 0 36320 800 36440
rect 159200 36184 160000 36304
rect 159200 35640 160000 35760
rect 159200 35232 160000 35352
rect 0 34688 800 34808
rect 159200 34688 160000 34808
rect 159200 34280 160000 34400
rect 159200 33736 160000 33856
rect 159200 33192 160000 33312
rect 0 32920 800 33040
rect 159200 32784 160000 32904
rect 159200 32240 160000 32360
rect 159200 31696 160000 31816
rect 0 31288 800 31408
rect 159200 31288 160000 31408
rect 159200 30744 160000 30864
rect 159200 30200 160000 30320
rect 159200 29792 160000 29912
rect 0 29520 800 29640
rect 159200 29248 160000 29368
rect 159200 28840 160000 28960
rect 159200 28296 160000 28416
rect 0 27888 800 28008
rect 159200 27752 160000 27872
rect 159200 27344 160000 27464
rect 159200 26800 160000 26920
rect 0 26120 800 26240
rect 159200 26256 160000 26376
rect 159200 25848 160000 25968
rect 159200 25304 160000 25424
rect 159200 24760 160000 24880
rect 0 24488 800 24608
rect 159200 24352 160000 24472
rect 159200 23808 160000 23928
rect 159200 23400 160000 23520
rect 0 22720 800 22840
rect 159200 22856 160000 22976
rect 159200 22312 160000 22432
rect 159200 21904 160000 22024
rect 159200 21360 160000 21480
rect 0 21088 800 21208
rect 159200 20816 160000 20936
rect 159200 20408 160000 20528
rect 159200 19864 160000 19984
rect 0 19456 800 19576
rect 159200 19320 160000 19440
rect 159200 18912 160000 19032
rect 159200 18368 160000 18488
rect 0 17688 800 17808
rect 159200 17824 160000 17944
rect 159200 17416 160000 17536
rect 159200 16872 160000 16992
rect 159200 16464 160000 16584
rect 0 16056 800 16176
rect 159200 15920 160000 16040
rect 159200 15376 160000 15496
rect 159200 14968 160000 15088
rect 0 14288 800 14408
rect 159200 14424 160000 14544
rect 159200 13880 160000 14000
rect 159200 13472 160000 13592
rect 159200 12928 160000 13048
rect 0 12656 800 12776
rect 159200 12384 160000 12504
rect 159200 11976 160000 12096
rect 159200 11432 160000 11552
rect 0 10888 800 11008
rect 159200 11024 160000 11144
rect 159200 10480 160000 10600
rect 159200 9936 160000 10056
rect 159200 9528 160000 9648
rect 0 9256 800 9376
rect 159200 8984 160000 9104
rect 159200 8440 160000 8560
rect 159200 8032 160000 8152
rect 0 7488 800 7608
rect 159200 7488 160000 7608
rect 159200 6944 160000 7064
rect 159200 6536 160000 6656
rect 0 5856 800 5976
rect 159200 5992 160000 6112
rect 159200 5584 160000 5704
rect 159200 5040 160000 5160
rect 159200 4496 160000 4616
rect 0 4088 800 4208
rect 159200 4088 160000 4208
rect 159200 3544 160000 3664
rect 159200 3000 160000 3120
rect 0 2456 800 2576
rect 159200 2592 160000 2712
rect 159200 2048 160000 2168
rect 159200 1504 160000 1624
rect 159200 1096 160000 1216
rect 0 824 800 944
rect 159200 552 160000 672
rect 159200 144 160000 264
<< obsm3 >>
rect 800 99480 159120 99653
rect 800 99216 159200 99480
rect 880 98936 159120 99216
rect 800 98808 159200 98936
rect 800 98528 159120 98808
rect 800 98264 159200 98528
rect 800 97984 159120 98264
rect 800 97720 159200 97984
rect 800 97584 159120 97720
rect 880 97440 159120 97584
rect 880 97312 159200 97440
rect 880 97304 159120 97312
rect 800 97032 159120 97304
rect 800 96768 159200 97032
rect 800 96488 159120 96768
rect 800 96224 159200 96488
rect 800 95944 159120 96224
rect 800 95816 159200 95944
rect 880 95536 159120 95816
rect 800 95272 159200 95536
rect 800 94992 159120 95272
rect 800 94728 159200 94992
rect 800 94448 159120 94728
rect 800 94320 159200 94448
rect 800 94184 159120 94320
rect 880 94040 159120 94184
rect 880 93904 159200 94040
rect 800 93776 159200 93904
rect 800 93496 159120 93776
rect 800 93368 159200 93496
rect 800 93088 159120 93368
rect 800 92824 159200 93088
rect 800 92544 159120 92824
rect 800 92416 159200 92544
rect 880 92280 159200 92416
rect 880 92136 159120 92280
rect 800 92000 159120 92136
rect 800 91872 159200 92000
rect 800 91592 159120 91872
rect 800 91328 159200 91592
rect 800 91048 159120 91328
rect 800 90784 159200 91048
rect 880 90504 159120 90784
rect 800 90376 159200 90504
rect 800 90096 159120 90376
rect 800 89832 159200 90096
rect 800 89552 159120 89832
rect 800 89288 159200 89552
rect 800 89016 159120 89288
rect 880 89008 159120 89016
rect 880 88880 159200 89008
rect 880 88736 159120 88880
rect 800 88600 159120 88736
rect 800 88336 159200 88600
rect 800 88056 159120 88336
rect 800 87928 159200 88056
rect 800 87648 159120 87928
rect 800 87384 159200 87648
rect 880 87104 159120 87384
rect 800 86840 159200 87104
rect 800 86560 159120 86840
rect 800 86432 159200 86560
rect 800 86152 159120 86432
rect 800 85888 159200 86152
rect 800 85616 159120 85888
rect 880 85608 159120 85616
rect 880 85344 159200 85608
rect 880 85336 159120 85344
rect 800 85064 159120 85336
rect 800 84936 159200 85064
rect 800 84656 159120 84936
rect 800 84392 159200 84656
rect 800 84112 159120 84392
rect 800 83984 159200 84112
rect 880 83848 159200 83984
rect 880 83704 159120 83848
rect 800 83568 159120 83704
rect 800 83440 159200 83568
rect 800 83160 159120 83440
rect 800 82896 159200 83160
rect 800 82616 159120 82896
rect 800 82488 159200 82616
rect 800 82216 159120 82488
rect 880 82208 159120 82216
rect 880 81944 159200 82208
rect 880 81936 159120 81944
rect 800 81664 159120 81936
rect 800 81400 159200 81664
rect 800 81120 159120 81400
rect 800 80992 159200 81120
rect 800 80712 159120 80992
rect 800 80584 159200 80712
rect 880 80448 159200 80584
rect 880 80304 159120 80448
rect 800 80168 159120 80304
rect 800 79904 159200 80168
rect 800 79624 159120 79904
rect 800 79496 159200 79624
rect 800 79216 159120 79496
rect 800 78952 159200 79216
rect 880 78672 159120 78952
rect 800 78408 159200 78672
rect 800 78128 159120 78408
rect 800 78000 159200 78128
rect 800 77720 159120 78000
rect 800 77456 159200 77720
rect 800 77184 159120 77456
rect 880 77176 159120 77184
rect 880 76912 159200 77176
rect 880 76904 159120 76912
rect 800 76632 159120 76904
rect 800 76504 159200 76632
rect 800 76224 159120 76504
rect 800 75960 159200 76224
rect 800 75680 159120 75960
rect 800 75552 159200 75680
rect 880 75272 159120 75552
rect 800 75008 159200 75272
rect 800 74728 159120 75008
rect 800 74464 159200 74728
rect 800 74184 159120 74464
rect 800 74056 159200 74184
rect 800 73784 159120 74056
rect 880 73776 159120 73784
rect 880 73512 159200 73776
rect 880 73504 159120 73512
rect 800 73232 159120 73504
rect 800 72968 159200 73232
rect 800 72688 159120 72968
rect 800 72560 159200 72688
rect 800 72280 159120 72560
rect 800 72152 159200 72280
rect 880 72016 159200 72152
rect 880 71872 159120 72016
rect 800 71736 159120 71872
rect 800 71472 159200 71736
rect 800 71192 159120 71472
rect 800 71064 159200 71192
rect 800 70784 159120 71064
rect 800 70520 159200 70784
rect 800 70384 159120 70520
rect 880 70240 159120 70384
rect 880 70112 159200 70240
rect 880 70104 159120 70112
rect 800 69832 159120 70104
rect 800 69568 159200 69832
rect 800 69288 159120 69568
rect 800 69024 159200 69288
rect 800 68752 159120 69024
rect 880 68744 159120 68752
rect 880 68616 159200 68744
rect 880 68472 159120 68616
rect 800 68336 159120 68472
rect 800 68072 159200 68336
rect 800 67792 159120 68072
rect 800 67528 159200 67792
rect 800 67248 159120 67528
rect 800 67120 159200 67248
rect 800 66984 159120 67120
rect 880 66840 159120 66984
rect 880 66704 159200 66840
rect 800 66576 159200 66704
rect 800 66296 159120 66576
rect 800 66032 159200 66296
rect 800 65752 159120 66032
rect 800 65624 159200 65752
rect 800 65352 159120 65624
rect 880 65344 159120 65352
rect 880 65080 159200 65344
rect 880 65072 159120 65080
rect 800 64800 159120 65072
rect 800 64672 159200 64800
rect 800 64392 159120 64672
rect 800 64128 159200 64392
rect 800 63848 159120 64128
rect 800 63584 159200 63848
rect 880 63304 159120 63584
rect 800 63176 159200 63304
rect 800 62896 159120 63176
rect 800 62632 159200 62896
rect 800 62352 159120 62632
rect 800 62088 159200 62352
rect 800 61952 159120 62088
rect 880 61808 159120 61952
rect 880 61680 159200 61808
rect 880 61672 159120 61680
rect 800 61400 159120 61672
rect 800 61136 159200 61400
rect 800 60856 159120 61136
rect 800 60592 159200 60856
rect 800 60320 159120 60592
rect 880 60312 159120 60320
rect 880 60184 159200 60312
rect 880 60040 159120 60184
rect 800 59904 159120 60040
rect 800 59640 159200 59904
rect 800 59360 159120 59640
rect 800 59096 159200 59360
rect 800 58816 159120 59096
rect 800 58688 159200 58816
rect 800 58552 159120 58688
rect 880 58408 159120 58552
rect 880 58272 159200 58408
rect 800 58144 159200 58272
rect 800 57864 159120 58144
rect 800 57736 159200 57864
rect 800 57456 159120 57736
rect 800 57192 159200 57456
rect 800 56920 159120 57192
rect 880 56912 159120 56920
rect 880 56648 159200 56912
rect 880 56640 159120 56648
rect 800 56368 159120 56640
rect 800 56240 159200 56368
rect 800 55960 159120 56240
rect 800 55696 159200 55960
rect 800 55416 159120 55696
rect 800 55152 159200 55416
rect 880 54872 159120 55152
rect 800 54744 159200 54872
rect 800 54464 159120 54744
rect 800 54200 159200 54464
rect 800 53920 159120 54200
rect 800 53656 159200 53920
rect 800 53520 159120 53656
rect 880 53376 159120 53520
rect 880 53248 159200 53376
rect 880 53240 159120 53248
rect 800 52968 159120 53240
rect 800 52704 159200 52968
rect 800 52424 159120 52704
rect 800 52296 159200 52424
rect 800 52016 159120 52296
rect 800 51752 159200 52016
rect 880 51472 159120 51752
rect 800 51208 159200 51472
rect 800 50928 159120 51208
rect 800 50800 159200 50928
rect 800 50520 159120 50800
rect 800 50256 159200 50520
rect 800 50120 159120 50256
rect 880 49976 159120 50120
rect 880 49840 159200 49976
rect 800 49712 159200 49840
rect 800 49432 159120 49712
rect 800 49304 159200 49432
rect 800 49024 159120 49304
rect 800 48760 159200 49024
rect 800 48480 159120 48760
rect 800 48352 159200 48480
rect 880 48216 159200 48352
rect 880 48072 159120 48216
rect 800 47936 159120 48072
rect 800 47808 159200 47936
rect 800 47528 159120 47808
rect 800 47264 159200 47528
rect 800 46984 159120 47264
rect 800 46856 159200 46984
rect 800 46720 159120 46856
rect 880 46576 159120 46720
rect 880 46440 159200 46576
rect 800 46312 159200 46440
rect 800 46032 159120 46312
rect 800 45768 159200 46032
rect 800 45488 159120 45768
rect 800 45360 159200 45488
rect 800 45080 159120 45360
rect 800 44952 159200 45080
rect 880 44816 159200 44952
rect 880 44672 159120 44816
rect 800 44536 159120 44672
rect 800 44272 159200 44536
rect 800 43992 159120 44272
rect 800 43864 159200 43992
rect 800 43584 159120 43864
rect 800 43320 159200 43584
rect 880 43040 159120 43320
rect 800 42776 159200 43040
rect 800 42496 159120 42776
rect 800 42368 159200 42496
rect 800 42088 159120 42368
rect 800 41824 159200 42088
rect 800 41552 159120 41824
rect 880 41544 159120 41552
rect 880 41416 159200 41544
rect 880 41272 159120 41416
rect 800 41136 159120 41272
rect 800 40872 159200 41136
rect 800 40592 159120 40872
rect 800 40328 159200 40592
rect 800 40048 159120 40328
rect 800 39920 159200 40048
rect 880 39640 159120 39920
rect 800 39376 159200 39640
rect 800 39096 159120 39376
rect 800 38832 159200 39096
rect 800 38552 159120 38832
rect 800 38424 159200 38552
rect 800 38288 159120 38424
rect 880 38144 159120 38288
rect 880 38008 159200 38144
rect 800 37880 159200 38008
rect 800 37600 159120 37880
rect 800 37336 159200 37600
rect 800 37056 159120 37336
rect 800 36928 159200 37056
rect 800 36648 159120 36928
rect 800 36520 159200 36648
rect 880 36384 159200 36520
rect 880 36240 159120 36384
rect 800 36104 159120 36240
rect 800 35840 159200 36104
rect 800 35560 159120 35840
rect 800 35432 159200 35560
rect 800 35152 159120 35432
rect 800 34888 159200 35152
rect 880 34608 159120 34888
rect 800 34480 159200 34608
rect 800 34200 159120 34480
rect 800 33936 159200 34200
rect 800 33656 159120 33936
rect 800 33392 159200 33656
rect 800 33120 159120 33392
rect 880 33112 159120 33120
rect 880 32984 159200 33112
rect 880 32840 159120 32984
rect 800 32704 159120 32840
rect 800 32440 159200 32704
rect 800 32160 159120 32440
rect 800 31896 159200 32160
rect 800 31616 159120 31896
rect 800 31488 159200 31616
rect 880 31208 159120 31488
rect 800 30944 159200 31208
rect 800 30664 159120 30944
rect 800 30400 159200 30664
rect 800 30120 159120 30400
rect 800 29992 159200 30120
rect 800 29720 159120 29992
rect 880 29712 159120 29720
rect 880 29448 159200 29712
rect 880 29440 159120 29448
rect 800 29168 159120 29440
rect 800 29040 159200 29168
rect 800 28760 159120 29040
rect 800 28496 159200 28760
rect 800 28216 159120 28496
rect 800 28088 159200 28216
rect 880 27952 159200 28088
rect 880 27808 159120 27952
rect 800 27672 159120 27808
rect 800 27544 159200 27672
rect 800 27264 159120 27544
rect 800 27000 159200 27264
rect 800 26720 159120 27000
rect 800 26456 159200 26720
rect 800 26320 159120 26456
rect 880 26176 159120 26320
rect 880 26048 159200 26176
rect 880 26040 159120 26048
rect 800 25768 159120 26040
rect 800 25504 159200 25768
rect 800 25224 159120 25504
rect 800 24960 159200 25224
rect 800 24688 159120 24960
rect 880 24680 159120 24688
rect 880 24552 159200 24680
rect 880 24408 159120 24552
rect 800 24272 159120 24408
rect 800 24008 159200 24272
rect 800 23728 159120 24008
rect 800 23600 159200 23728
rect 800 23320 159120 23600
rect 800 23056 159200 23320
rect 800 22920 159120 23056
rect 880 22776 159120 22920
rect 880 22640 159200 22776
rect 800 22512 159200 22640
rect 800 22232 159120 22512
rect 800 22104 159200 22232
rect 800 21824 159120 22104
rect 800 21560 159200 21824
rect 800 21288 159120 21560
rect 880 21280 159120 21288
rect 880 21016 159200 21280
rect 880 21008 159120 21016
rect 800 20736 159120 21008
rect 800 20608 159200 20736
rect 800 20328 159120 20608
rect 800 20064 159200 20328
rect 800 19784 159120 20064
rect 800 19656 159200 19784
rect 880 19520 159200 19656
rect 880 19376 159120 19520
rect 800 19240 159120 19376
rect 800 19112 159200 19240
rect 800 18832 159120 19112
rect 800 18568 159200 18832
rect 800 18288 159120 18568
rect 800 18024 159200 18288
rect 800 17888 159120 18024
rect 880 17744 159120 17888
rect 880 17616 159200 17744
rect 880 17608 159120 17616
rect 800 17336 159120 17608
rect 800 17072 159200 17336
rect 800 16792 159120 17072
rect 800 16664 159200 16792
rect 800 16384 159120 16664
rect 800 16256 159200 16384
rect 880 16120 159200 16256
rect 880 15976 159120 16120
rect 800 15840 159120 15976
rect 800 15576 159200 15840
rect 800 15296 159120 15576
rect 800 15168 159200 15296
rect 800 14888 159120 15168
rect 800 14624 159200 14888
rect 800 14488 159120 14624
rect 880 14344 159120 14488
rect 880 14208 159200 14344
rect 800 14080 159200 14208
rect 800 13800 159120 14080
rect 800 13672 159200 13800
rect 800 13392 159120 13672
rect 800 13128 159200 13392
rect 800 12856 159120 13128
rect 880 12848 159120 12856
rect 880 12584 159200 12848
rect 880 12576 159120 12584
rect 800 12304 159120 12576
rect 800 12176 159200 12304
rect 800 11896 159120 12176
rect 800 11632 159200 11896
rect 800 11352 159120 11632
rect 800 11224 159200 11352
rect 800 11088 159120 11224
rect 880 10944 159120 11088
rect 880 10808 159200 10944
rect 800 10680 159200 10808
rect 800 10400 159120 10680
rect 800 10136 159200 10400
rect 800 9856 159120 10136
rect 800 9728 159200 9856
rect 800 9456 159120 9728
rect 880 9448 159120 9456
rect 880 9184 159200 9448
rect 880 9176 159120 9184
rect 800 8904 159120 9176
rect 800 8640 159200 8904
rect 800 8360 159120 8640
rect 800 8232 159200 8360
rect 800 7952 159120 8232
rect 800 7688 159200 7952
rect 880 7408 159120 7688
rect 800 7144 159200 7408
rect 800 6864 159120 7144
rect 800 6736 159200 6864
rect 800 6456 159120 6736
rect 800 6192 159200 6456
rect 800 6056 159120 6192
rect 880 5912 159120 6056
rect 880 5784 159200 5912
rect 880 5776 159120 5784
rect 800 5504 159120 5776
rect 800 5240 159200 5504
rect 800 4960 159120 5240
rect 800 4696 159200 4960
rect 800 4416 159120 4696
rect 800 4288 159200 4416
rect 880 4008 159120 4288
rect 800 3744 159200 4008
rect 800 3464 159120 3744
rect 800 3200 159200 3464
rect 800 2920 159120 3200
rect 800 2792 159200 2920
rect 800 2656 159120 2792
rect 880 2512 159120 2656
rect 880 2376 159200 2512
rect 800 2248 159200 2376
rect 800 1968 159120 2248
rect 800 1704 159200 1968
rect 800 1424 159120 1704
rect 800 1296 159200 1424
rect 800 1024 159120 1296
rect 880 1016 159120 1024
rect 880 752 159200 1016
rect 880 744 159120 752
rect 800 472 159120 744
rect 800 344 159200 472
rect 800 171 159120 344
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
rect 111728 2128 112048 97424
rect 127088 2128 127408 97424
rect 142448 2128 142768 97424
rect 157808 2128 158128 97424
<< obsm4 >>
rect 155723 88163 155789 92581
<< labels >>
rlabel metal2 s 7102 99200 7158 100000 6 addr0[0]
port 1 nsew signal output
rlabel metal2 s 7930 99200 7986 100000 6 addr0[1]
port 2 nsew signal output
rlabel metal2 s 8850 99200 8906 100000 6 addr0[2]
port 3 nsew signal output
rlabel metal2 s 9678 99200 9734 100000 6 addr0[3]
port 4 nsew signal output
rlabel metal2 s 10506 99200 10562 100000 6 addr0[4]
port 5 nsew signal output
rlabel metal2 s 11334 99200 11390 100000 6 addr0[5]
port 6 nsew signal output
rlabel metal2 s 12162 99200 12218 100000 6 addr0[6]
port 7 nsew signal output
rlabel metal2 s 13082 99200 13138 100000 6 addr0[7]
port 8 nsew signal output
rlabel metal2 s 13910 99200 13966 100000 6 addr0[8]
port 9 nsew signal output
rlabel metal2 s 98550 99200 98606 100000 6 addr1[0]
port 10 nsew signal output
rlabel metal2 s 99378 99200 99434 100000 6 addr1[1]
port 11 nsew signal output
rlabel metal2 s 100206 99200 100262 100000 6 addr1[2]
port 12 nsew signal output
rlabel metal2 s 101034 99200 101090 100000 6 addr1[3]
port 13 nsew signal output
rlabel metal2 s 101954 99200 102010 100000 6 addr1[4]
port 14 nsew signal output
rlabel metal2 s 102782 99200 102838 100000 6 addr1[5]
port 15 nsew signal output
rlabel metal2 s 103610 99200 103666 100000 6 addr1[6]
port 16 nsew signal output
rlabel metal2 s 104438 99200 104494 100000 6 addr1[7]
port 17 nsew signal output
rlabel metal2 s 105266 99200 105322 100000 6 addr1[8]
port 18 nsew signal output
rlabel metal2 s 386 99200 442 100000 6 clk0
port 19 nsew signal output
rlabel metal2 s 95974 99200 96030 100000 6 clk1
port 20 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 coreIndex[0]
port 21 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 coreIndex[1]
port 22 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 coreIndex[2]
port 23 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 coreIndex[3]
port 24 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 coreIndex[4]
port 25 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 coreIndex[5]
port 26 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 coreIndex[6]
port 27 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 coreIndex[7]
port 28 nsew signal input
rlabel metal3 s 159200 1096 160000 1216 6 core_wb_ack_i
port 29 nsew signal input
rlabel metal3 s 159200 4088 160000 4208 6 core_wb_adr_o[0]
port 30 nsew signal output
rlabel metal3 s 159200 20816 160000 20936 6 core_wb_adr_o[10]
port 31 nsew signal output
rlabel metal3 s 159200 22312 160000 22432 6 core_wb_adr_o[11]
port 32 nsew signal output
rlabel metal3 s 159200 23808 160000 23928 6 core_wb_adr_o[12]
port 33 nsew signal output
rlabel metal3 s 159200 25304 160000 25424 6 core_wb_adr_o[13]
port 34 nsew signal output
rlabel metal3 s 159200 26800 160000 26920 6 core_wb_adr_o[14]
port 35 nsew signal output
rlabel metal3 s 159200 28296 160000 28416 6 core_wb_adr_o[15]
port 36 nsew signal output
rlabel metal3 s 159200 29792 160000 29912 6 core_wb_adr_o[16]
port 37 nsew signal output
rlabel metal3 s 159200 31288 160000 31408 6 core_wb_adr_o[17]
port 38 nsew signal output
rlabel metal3 s 159200 32784 160000 32904 6 core_wb_adr_o[18]
port 39 nsew signal output
rlabel metal3 s 159200 34280 160000 34400 6 core_wb_adr_o[19]
port 40 nsew signal output
rlabel metal3 s 159200 5992 160000 6112 6 core_wb_adr_o[1]
port 41 nsew signal output
rlabel metal3 s 159200 35640 160000 35760 6 core_wb_adr_o[20]
port 42 nsew signal output
rlabel metal3 s 159200 37136 160000 37256 6 core_wb_adr_o[21]
port 43 nsew signal output
rlabel metal3 s 159200 38632 160000 38752 6 core_wb_adr_o[22]
port 44 nsew signal output
rlabel metal3 s 159200 40128 160000 40248 6 core_wb_adr_o[23]
port 45 nsew signal output
rlabel metal3 s 159200 41624 160000 41744 6 core_wb_adr_o[24]
port 46 nsew signal output
rlabel metal3 s 159200 43120 160000 43240 6 core_wb_adr_o[25]
port 47 nsew signal output
rlabel metal3 s 159200 44616 160000 44736 6 core_wb_adr_o[26]
port 48 nsew signal output
rlabel metal3 s 159200 46112 160000 46232 6 core_wb_adr_o[27]
port 49 nsew signal output
rlabel metal3 s 159200 8032 160000 8152 6 core_wb_adr_o[2]
port 50 nsew signal output
rlabel metal3 s 159200 9936 160000 10056 6 core_wb_adr_o[3]
port 51 nsew signal output
rlabel metal3 s 159200 11976 160000 12096 6 core_wb_adr_o[4]
port 52 nsew signal output
rlabel metal3 s 159200 13472 160000 13592 6 core_wb_adr_o[5]
port 53 nsew signal output
rlabel metal3 s 159200 14968 160000 15088 6 core_wb_adr_o[6]
port 54 nsew signal output
rlabel metal3 s 159200 16464 160000 16584 6 core_wb_adr_o[7]
port 55 nsew signal output
rlabel metal3 s 159200 17824 160000 17944 6 core_wb_adr_o[8]
port 56 nsew signal output
rlabel metal3 s 159200 19320 160000 19440 6 core_wb_adr_o[9]
port 57 nsew signal output
rlabel metal3 s 159200 1504 160000 1624 6 core_wb_cyc_o
port 58 nsew signal output
rlabel metal3 s 159200 4496 160000 4616 6 core_wb_data_i[0]
port 59 nsew signal input
rlabel metal3 s 159200 21360 160000 21480 6 core_wb_data_i[10]
port 60 nsew signal input
rlabel metal3 s 159200 22856 160000 22976 6 core_wb_data_i[11]
port 61 nsew signal input
rlabel metal3 s 159200 24352 160000 24472 6 core_wb_data_i[12]
port 62 nsew signal input
rlabel metal3 s 159200 25848 160000 25968 6 core_wb_data_i[13]
port 63 nsew signal input
rlabel metal3 s 159200 27344 160000 27464 6 core_wb_data_i[14]
port 64 nsew signal input
rlabel metal3 s 159200 28840 160000 28960 6 core_wb_data_i[15]
port 65 nsew signal input
rlabel metal3 s 159200 30200 160000 30320 6 core_wb_data_i[16]
port 66 nsew signal input
rlabel metal3 s 159200 31696 160000 31816 6 core_wb_data_i[17]
port 67 nsew signal input
rlabel metal3 s 159200 33192 160000 33312 6 core_wb_data_i[18]
port 68 nsew signal input
rlabel metal3 s 159200 34688 160000 34808 6 core_wb_data_i[19]
port 69 nsew signal input
rlabel metal3 s 159200 6536 160000 6656 6 core_wb_data_i[1]
port 70 nsew signal input
rlabel metal3 s 159200 36184 160000 36304 6 core_wb_data_i[20]
port 71 nsew signal input
rlabel metal3 s 159200 37680 160000 37800 6 core_wb_data_i[21]
port 72 nsew signal input
rlabel metal3 s 159200 39176 160000 39296 6 core_wb_data_i[22]
port 73 nsew signal input
rlabel metal3 s 159200 40672 160000 40792 6 core_wb_data_i[23]
port 74 nsew signal input
rlabel metal3 s 159200 42168 160000 42288 6 core_wb_data_i[24]
port 75 nsew signal input
rlabel metal3 s 159200 43664 160000 43784 6 core_wb_data_i[25]
port 76 nsew signal input
rlabel metal3 s 159200 45160 160000 45280 6 core_wb_data_i[26]
port 77 nsew signal input
rlabel metal3 s 159200 46656 160000 46776 6 core_wb_data_i[27]
port 78 nsew signal input
rlabel metal3 s 159200 47608 160000 47728 6 core_wb_data_i[28]
port 79 nsew signal input
rlabel metal3 s 159200 48560 160000 48680 6 core_wb_data_i[29]
port 80 nsew signal input
rlabel metal3 s 159200 8440 160000 8560 6 core_wb_data_i[2]
port 81 nsew signal input
rlabel metal3 s 159200 49512 160000 49632 6 core_wb_data_i[30]
port 82 nsew signal input
rlabel metal3 s 159200 50600 160000 50720 6 core_wb_data_i[31]
port 83 nsew signal input
rlabel metal3 s 159200 10480 160000 10600 6 core_wb_data_i[3]
port 84 nsew signal input
rlabel metal3 s 159200 12384 160000 12504 6 core_wb_data_i[4]
port 85 nsew signal input
rlabel metal3 s 159200 13880 160000 14000 6 core_wb_data_i[5]
port 86 nsew signal input
rlabel metal3 s 159200 15376 160000 15496 6 core_wb_data_i[6]
port 87 nsew signal input
rlabel metal3 s 159200 16872 160000 16992 6 core_wb_data_i[7]
port 88 nsew signal input
rlabel metal3 s 159200 18368 160000 18488 6 core_wb_data_i[8]
port 89 nsew signal input
rlabel metal3 s 159200 19864 160000 19984 6 core_wb_data_i[9]
port 90 nsew signal input
rlabel metal3 s 159200 5040 160000 5160 6 core_wb_data_o[0]
port 91 nsew signal output
rlabel metal3 s 159200 21904 160000 22024 6 core_wb_data_o[10]
port 92 nsew signal output
rlabel metal3 s 159200 23400 160000 23520 6 core_wb_data_o[11]
port 93 nsew signal output
rlabel metal3 s 159200 24760 160000 24880 6 core_wb_data_o[12]
port 94 nsew signal output
rlabel metal3 s 159200 26256 160000 26376 6 core_wb_data_o[13]
port 95 nsew signal output
rlabel metal3 s 159200 27752 160000 27872 6 core_wb_data_o[14]
port 96 nsew signal output
rlabel metal3 s 159200 29248 160000 29368 6 core_wb_data_o[15]
port 97 nsew signal output
rlabel metal3 s 159200 30744 160000 30864 6 core_wb_data_o[16]
port 98 nsew signal output
rlabel metal3 s 159200 32240 160000 32360 6 core_wb_data_o[17]
port 99 nsew signal output
rlabel metal3 s 159200 33736 160000 33856 6 core_wb_data_o[18]
port 100 nsew signal output
rlabel metal3 s 159200 35232 160000 35352 6 core_wb_data_o[19]
port 101 nsew signal output
rlabel metal3 s 159200 6944 160000 7064 6 core_wb_data_o[1]
port 102 nsew signal output
rlabel metal3 s 159200 36728 160000 36848 6 core_wb_data_o[20]
port 103 nsew signal output
rlabel metal3 s 159200 38224 160000 38344 6 core_wb_data_o[21]
port 104 nsew signal output
rlabel metal3 s 159200 39720 160000 39840 6 core_wb_data_o[22]
port 105 nsew signal output
rlabel metal3 s 159200 41216 160000 41336 6 core_wb_data_o[23]
port 106 nsew signal output
rlabel metal3 s 159200 42576 160000 42696 6 core_wb_data_o[24]
port 107 nsew signal output
rlabel metal3 s 159200 44072 160000 44192 6 core_wb_data_o[25]
port 108 nsew signal output
rlabel metal3 s 159200 45568 160000 45688 6 core_wb_data_o[26]
port 109 nsew signal output
rlabel metal3 s 159200 47064 160000 47184 6 core_wb_data_o[27]
port 110 nsew signal output
rlabel metal3 s 159200 48016 160000 48136 6 core_wb_data_o[28]
port 111 nsew signal output
rlabel metal3 s 159200 49104 160000 49224 6 core_wb_data_o[29]
port 112 nsew signal output
rlabel metal3 s 159200 8984 160000 9104 6 core_wb_data_o[2]
port 113 nsew signal output
rlabel metal3 s 159200 50056 160000 50176 6 core_wb_data_o[30]
port 114 nsew signal output
rlabel metal3 s 159200 51008 160000 51128 6 core_wb_data_o[31]
port 115 nsew signal output
rlabel metal3 s 159200 11024 160000 11144 6 core_wb_data_o[3]
port 116 nsew signal output
rlabel metal3 s 159200 12928 160000 13048 6 core_wb_data_o[4]
port 117 nsew signal output
rlabel metal3 s 159200 14424 160000 14544 6 core_wb_data_o[5]
port 118 nsew signal output
rlabel metal3 s 159200 15920 160000 16040 6 core_wb_data_o[6]
port 119 nsew signal output
rlabel metal3 s 159200 17416 160000 17536 6 core_wb_data_o[7]
port 120 nsew signal output
rlabel metal3 s 159200 18912 160000 19032 6 core_wb_data_o[8]
port 121 nsew signal output
rlabel metal3 s 159200 20408 160000 20528 6 core_wb_data_o[9]
port 122 nsew signal output
rlabel metal3 s 159200 2048 160000 2168 6 core_wb_error_i
port 123 nsew signal input
rlabel metal3 s 159200 5584 160000 5704 6 core_wb_sel_o[0]
port 124 nsew signal output
rlabel metal3 s 159200 7488 160000 7608 6 core_wb_sel_o[1]
port 125 nsew signal output
rlabel metal3 s 159200 9528 160000 9648 6 core_wb_sel_o[2]
port 126 nsew signal output
rlabel metal3 s 159200 11432 160000 11552 6 core_wb_sel_o[3]
port 127 nsew signal output
rlabel metal3 s 159200 2592 160000 2712 6 core_wb_stall_i
port 128 nsew signal input
rlabel metal3 s 159200 3000 160000 3120 6 core_wb_stb_o
port 129 nsew signal output
rlabel metal3 s 159200 3544 160000 3664 6 core_wb_we_o
port 130 nsew signal output
rlabel metal2 s 1214 99200 1270 100000 6 csb0[0]
port 131 nsew signal output
rlabel metal2 s 2042 99200 2098 100000 6 csb0[1]
port 132 nsew signal output
rlabel metal2 s 96802 99200 96858 100000 6 csb1[0]
port 133 nsew signal output
rlabel metal2 s 97722 99200 97778 100000 6 csb1[1]
port 134 nsew signal output
rlabel metal2 s 14738 99200 14794 100000 6 din0[0]
port 135 nsew signal output
rlabel metal2 s 23202 99200 23258 100000 6 din0[10]
port 136 nsew signal output
rlabel metal2 s 24030 99200 24086 100000 6 din0[11]
port 137 nsew signal output
rlabel metal2 s 24858 99200 24914 100000 6 din0[12]
port 138 nsew signal output
rlabel metal2 s 25778 99200 25834 100000 6 din0[13]
port 139 nsew signal output
rlabel metal2 s 26606 99200 26662 100000 6 din0[14]
port 140 nsew signal output
rlabel metal2 s 27434 99200 27490 100000 6 din0[15]
port 141 nsew signal output
rlabel metal2 s 28262 99200 28318 100000 6 din0[16]
port 142 nsew signal output
rlabel metal2 s 29090 99200 29146 100000 6 din0[17]
port 143 nsew signal output
rlabel metal2 s 30010 99200 30066 100000 6 din0[18]
port 144 nsew signal output
rlabel metal2 s 30838 99200 30894 100000 6 din0[19]
port 145 nsew signal output
rlabel metal2 s 15566 99200 15622 100000 6 din0[1]
port 146 nsew signal output
rlabel metal2 s 31666 99200 31722 100000 6 din0[20]
port 147 nsew signal output
rlabel metal2 s 32494 99200 32550 100000 6 din0[21]
port 148 nsew signal output
rlabel metal2 s 33322 99200 33378 100000 6 din0[22]
port 149 nsew signal output
rlabel metal2 s 34242 99200 34298 100000 6 din0[23]
port 150 nsew signal output
rlabel metal2 s 35070 99200 35126 100000 6 din0[24]
port 151 nsew signal output
rlabel metal2 s 35898 99200 35954 100000 6 din0[25]
port 152 nsew signal output
rlabel metal2 s 36726 99200 36782 100000 6 din0[26]
port 153 nsew signal output
rlabel metal2 s 37554 99200 37610 100000 6 din0[27]
port 154 nsew signal output
rlabel metal2 s 38474 99200 38530 100000 6 din0[28]
port 155 nsew signal output
rlabel metal2 s 39302 99200 39358 100000 6 din0[29]
port 156 nsew signal output
rlabel metal2 s 16394 99200 16450 100000 6 din0[2]
port 157 nsew signal output
rlabel metal2 s 40130 99200 40186 100000 6 din0[30]
port 158 nsew signal output
rlabel metal2 s 40958 99200 41014 100000 6 din0[31]
port 159 nsew signal output
rlabel metal2 s 17314 99200 17370 100000 6 din0[3]
port 160 nsew signal output
rlabel metal2 s 18142 99200 18198 100000 6 din0[4]
port 161 nsew signal output
rlabel metal2 s 18970 99200 19026 100000 6 din0[5]
port 162 nsew signal output
rlabel metal2 s 19798 99200 19854 100000 6 din0[6]
port 163 nsew signal output
rlabel metal2 s 20626 99200 20682 100000 6 din0[7]
port 164 nsew signal output
rlabel metal2 s 21546 99200 21602 100000 6 din0[8]
port 165 nsew signal output
rlabel metal2 s 22374 99200 22430 100000 6 din0[9]
port 166 nsew signal output
rlabel metal2 s 41786 99200 41842 100000 6 dout0[0]
port 167 nsew signal input
rlabel metal2 s 50250 99200 50306 100000 6 dout0[10]
port 168 nsew signal input
rlabel metal2 s 51170 99200 51226 100000 6 dout0[11]
port 169 nsew signal input
rlabel metal2 s 51998 99200 52054 100000 6 dout0[12]
port 170 nsew signal input
rlabel metal2 s 52826 99200 52882 100000 6 dout0[13]
port 171 nsew signal input
rlabel metal2 s 53654 99200 53710 100000 6 dout0[14]
port 172 nsew signal input
rlabel metal2 s 54482 99200 54538 100000 6 dout0[15]
port 173 nsew signal input
rlabel metal2 s 55402 99200 55458 100000 6 dout0[16]
port 174 nsew signal input
rlabel metal2 s 56230 99200 56286 100000 6 dout0[17]
port 175 nsew signal input
rlabel metal2 s 57058 99200 57114 100000 6 dout0[18]
port 176 nsew signal input
rlabel metal2 s 57886 99200 57942 100000 6 dout0[19]
port 177 nsew signal input
rlabel metal2 s 42706 99200 42762 100000 6 dout0[1]
port 178 nsew signal input
rlabel metal2 s 58714 99200 58770 100000 6 dout0[20]
port 179 nsew signal input
rlabel metal2 s 59634 99200 59690 100000 6 dout0[21]
port 180 nsew signal input
rlabel metal2 s 60462 99200 60518 100000 6 dout0[22]
port 181 nsew signal input
rlabel metal2 s 61290 99200 61346 100000 6 dout0[23]
port 182 nsew signal input
rlabel metal2 s 62118 99200 62174 100000 6 dout0[24]
port 183 nsew signal input
rlabel metal2 s 62946 99200 63002 100000 6 dout0[25]
port 184 nsew signal input
rlabel metal2 s 63866 99200 63922 100000 6 dout0[26]
port 185 nsew signal input
rlabel metal2 s 64694 99200 64750 100000 6 dout0[27]
port 186 nsew signal input
rlabel metal2 s 65522 99200 65578 100000 6 dout0[28]
port 187 nsew signal input
rlabel metal2 s 66350 99200 66406 100000 6 dout0[29]
port 188 nsew signal input
rlabel metal2 s 43534 99200 43590 100000 6 dout0[2]
port 189 nsew signal input
rlabel metal2 s 67178 99200 67234 100000 6 dout0[30]
port 190 nsew signal input
rlabel metal2 s 68098 99200 68154 100000 6 dout0[31]
port 191 nsew signal input
rlabel metal2 s 68926 99200 68982 100000 6 dout0[32]
port 192 nsew signal input
rlabel metal2 s 69754 99200 69810 100000 6 dout0[33]
port 193 nsew signal input
rlabel metal2 s 70582 99200 70638 100000 6 dout0[34]
port 194 nsew signal input
rlabel metal2 s 71410 99200 71466 100000 6 dout0[35]
port 195 nsew signal input
rlabel metal2 s 72330 99200 72386 100000 6 dout0[36]
port 196 nsew signal input
rlabel metal2 s 73158 99200 73214 100000 6 dout0[37]
port 197 nsew signal input
rlabel metal2 s 73986 99200 74042 100000 6 dout0[38]
port 198 nsew signal input
rlabel metal2 s 74814 99200 74870 100000 6 dout0[39]
port 199 nsew signal input
rlabel metal2 s 44362 99200 44418 100000 6 dout0[3]
port 200 nsew signal input
rlabel metal2 s 75642 99200 75698 100000 6 dout0[40]
port 201 nsew signal input
rlabel metal2 s 76562 99200 76618 100000 6 dout0[41]
port 202 nsew signal input
rlabel metal2 s 77390 99200 77446 100000 6 dout0[42]
port 203 nsew signal input
rlabel metal2 s 78218 99200 78274 100000 6 dout0[43]
port 204 nsew signal input
rlabel metal2 s 79046 99200 79102 100000 6 dout0[44]
port 205 nsew signal input
rlabel metal2 s 79874 99200 79930 100000 6 dout0[45]
port 206 nsew signal input
rlabel metal2 s 80794 99200 80850 100000 6 dout0[46]
port 207 nsew signal input
rlabel metal2 s 81622 99200 81678 100000 6 dout0[47]
port 208 nsew signal input
rlabel metal2 s 82450 99200 82506 100000 6 dout0[48]
port 209 nsew signal input
rlabel metal2 s 83278 99200 83334 100000 6 dout0[49]
port 210 nsew signal input
rlabel metal2 s 45190 99200 45246 100000 6 dout0[4]
port 211 nsew signal input
rlabel metal2 s 84106 99200 84162 100000 6 dout0[50]
port 212 nsew signal input
rlabel metal2 s 85026 99200 85082 100000 6 dout0[51]
port 213 nsew signal input
rlabel metal2 s 85854 99200 85910 100000 6 dout0[52]
port 214 nsew signal input
rlabel metal2 s 86682 99200 86738 100000 6 dout0[53]
port 215 nsew signal input
rlabel metal2 s 87510 99200 87566 100000 6 dout0[54]
port 216 nsew signal input
rlabel metal2 s 88338 99200 88394 100000 6 dout0[55]
port 217 nsew signal input
rlabel metal2 s 89258 99200 89314 100000 6 dout0[56]
port 218 nsew signal input
rlabel metal2 s 90086 99200 90142 100000 6 dout0[57]
port 219 nsew signal input
rlabel metal2 s 90914 99200 90970 100000 6 dout0[58]
port 220 nsew signal input
rlabel metal2 s 91742 99200 91798 100000 6 dout0[59]
port 221 nsew signal input
rlabel metal2 s 46018 99200 46074 100000 6 dout0[5]
port 222 nsew signal input
rlabel metal2 s 92570 99200 92626 100000 6 dout0[60]
port 223 nsew signal input
rlabel metal2 s 93490 99200 93546 100000 6 dout0[61]
port 224 nsew signal input
rlabel metal2 s 94318 99200 94374 100000 6 dout0[62]
port 225 nsew signal input
rlabel metal2 s 95146 99200 95202 100000 6 dout0[63]
port 226 nsew signal input
rlabel metal2 s 46938 99200 46994 100000 6 dout0[6]
port 227 nsew signal input
rlabel metal2 s 47766 99200 47822 100000 6 dout0[7]
port 228 nsew signal input
rlabel metal2 s 48594 99200 48650 100000 6 dout0[8]
port 229 nsew signal input
rlabel metal2 s 49422 99200 49478 100000 6 dout0[9]
port 230 nsew signal input
rlabel metal2 s 106186 99200 106242 100000 6 dout1[0]
port 231 nsew signal input
rlabel metal2 s 114650 99200 114706 100000 6 dout1[10]
port 232 nsew signal input
rlabel metal2 s 115478 99200 115534 100000 6 dout1[11]
port 233 nsew signal input
rlabel metal2 s 116306 99200 116362 100000 6 dout1[12]
port 234 nsew signal input
rlabel metal2 s 117134 99200 117190 100000 6 dout1[13]
port 235 nsew signal input
rlabel metal2 s 117962 99200 118018 100000 6 dout1[14]
port 236 nsew signal input
rlabel metal2 s 118882 99200 118938 100000 6 dout1[15]
port 237 nsew signal input
rlabel metal2 s 119710 99200 119766 100000 6 dout1[16]
port 238 nsew signal input
rlabel metal2 s 120538 99200 120594 100000 6 dout1[17]
port 239 nsew signal input
rlabel metal2 s 121366 99200 121422 100000 6 dout1[18]
port 240 nsew signal input
rlabel metal2 s 122194 99200 122250 100000 6 dout1[19]
port 241 nsew signal input
rlabel metal2 s 107014 99200 107070 100000 6 dout1[1]
port 242 nsew signal input
rlabel metal2 s 123114 99200 123170 100000 6 dout1[20]
port 243 nsew signal input
rlabel metal2 s 123942 99200 123998 100000 6 dout1[21]
port 244 nsew signal input
rlabel metal2 s 124770 99200 124826 100000 6 dout1[22]
port 245 nsew signal input
rlabel metal2 s 125598 99200 125654 100000 6 dout1[23]
port 246 nsew signal input
rlabel metal2 s 126426 99200 126482 100000 6 dout1[24]
port 247 nsew signal input
rlabel metal2 s 127346 99200 127402 100000 6 dout1[25]
port 248 nsew signal input
rlabel metal2 s 128174 99200 128230 100000 6 dout1[26]
port 249 nsew signal input
rlabel metal2 s 129002 99200 129058 100000 6 dout1[27]
port 250 nsew signal input
rlabel metal2 s 129830 99200 129886 100000 6 dout1[28]
port 251 nsew signal input
rlabel metal2 s 130658 99200 130714 100000 6 dout1[29]
port 252 nsew signal input
rlabel metal2 s 107842 99200 107898 100000 6 dout1[2]
port 253 nsew signal input
rlabel metal2 s 131578 99200 131634 100000 6 dout1[30]
port 254 nsew signal input
rlabel metal2 s 132406 99200 132462 100000 6 dout1[31]
port 255 nsew signal input
rlabel metal2 s 133234 99200 133290 100000 6 dout1[32]
port 256 nsew signal input
rlabel metal2 s 134062 99200 134118 100000 6 dout1[33]
port 257 nsew signal input
rlabel metal2 s 134890 99200 134946 100000 6 dout1[34]
port 258 nsew signal input
rlabel metal2 s 135810 99200 135866 100000 6 dout1[35]
port 259 nsew signal input
rlabel metal2 s 136638 99200 136694 100000 6 dout1[36]
port 260 nsew signal input
rlabel metal2 s 137466 99200 137522 100000 6 dout1[37]
port 261 nsew signal input
rlabel metal2 s 138294 99200 138350 100000 6 dout1[38]
port 262 nsew signal input
rlabel metal2 s 139122 99200 139178 100000 6 dout1[39]
port 263 nsew signal input
rlabel metal2 s 108670 99200 108726 100000 6 dout1[3]
port 264 nsew signal input
rlabel metal2 s 140042 99200 140098 100000 6 dout1[40]
port 265 nsew signal input
rlabel metal2 s 140870 99200 140926 100000 6 dout1[41]
port 266 nsew signal input
rlabel metal2 s 141698 99200 141754 100000 6 dout1[42]
port 267 nsew signal input
rlabel metal2 s 142526 99200 142582 100000 6 dout1[43]
port 268 nsew signal input
rlabel metal2 s 143354 99200 143410 100000 6 dout1[44]
port 269 nsew signal input
rlabel metal2 s 144274 99200 144330 100000 6 dout1[45]
port 270 nsew signal input
rlabel metal2 s 145102 99200 145158 100000 6 dout1[46]
port 271 nsew signal input
rlabel metal2 s 145930 99200 145986 100000 6 dout1[47]
port 272 nsew signal input
rlabel metal2 s 146758 99200 146814 100000 6 dout1[48]
port 273 nsew signal input
rlabel metal2 s 147586 99200 147642 100000 6 dout1[49]
port 274 nsew signal input
rlabel metal2 s 109498 99200 109554 100000 6 dout1[4]
port 275 nsew signal input
rlabel metal2 s 148506 99200 148562 100000 6 dout1[50]
port 276 nsew signal input
rlabel metal2 s 149334 99200 149390 100000 6 dout1[51]
port 277 nsew signal input
rlabel metal2 s 150162 99200 150218 100000 6 dout1[52]
port 278 nsew signal input
rlabel metal2 s 150990 99200 151046 100000 6 dout1[53]
port 279 nsew signal input
rlabel metal2 s 151818 99200 151874 100000 6 dout1[54]
port 280 nsew signal input
rlabel metal2 s 152738 99200 152794 100000 6 dout1[55]
port 281 nsew signal input
rlabel metal2 s 153566 99200 153622 100000 6 dout1[56]
port 282 nsew signal input
rlabel metal2 s 154394 99200 154450 100000 6 dout1[57]
port 283 nsew signal input
rlabel metal2 s 155222 99200 155278 100000 6 dout1[58]
port 284 nsew signal input
rlabel metal2 s 156050 99200 156106 100000 6 dout1[59]
port 285 nsew signal input
rlabel metal2 s 110418 99200 110474 100000 6 dout1[5]
port 286 nsew signal input
rlabel metal2 s 156970 99200 157026 100000 6 dout1[60]
port 287 nsew signal input
rlabel metal2 s 157798 99200 157854 100000 6 dout1[61]
port 288 nsew signal input
rlabel metal2 s 158626 99200 158682 100000 6 dout1[62]
port 289 nsew signal input
rlabel metal2 s 159454 99200 159510 100000 6 dout1[63]
port 290 nsew signal input
rlabel metal2 s 111246 99200 111302 100000 6 dout1[6]
port 291 nsew signal input
rlabel metal2 s 112074 99200 112130 100000 6 dout1[7]
port 292 nsew signal input
rlabel metal2 s 112902 99200 112958 100000 6 dout1[8]
port 293 nsew signal input
rlabel metal2 s 113730 99200 113786 100000 6 dout1[9]
port 294 nsew signal input
rlabel metal3 s 0 824 800 944 6 jtag_tck
port 295 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 jtag_tdi
port 296 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 jtag_tdo
port 297 nsew signal output
rlabel metal3 s 0 5856 800 5976 6 jtag_tms
port 298 nsew signal input
rlabel metal3 s 159200 51552 160000 51672 6 localMemory_wb_ack_o
port 299 nsew signal output
rlabel metal3 s 159200 54544 160000 54664 6 localMemory_wb_adr_i[0]
port 300 nsew signal input
rlabel metal3 s 159200 71272 160000 71392 6 localMemory_wb_adr_i[10]
port 301 nsew signal input
rlabel metal3 s 159200 72768 160000 72888 6 localMemory_wb_adr_i[11]
port 302 nsew signal input
rlabel metal3 s 159200 74264 160000 74384 6 localMemory_wb_adr_i[12]
port 303 nsew signal input
rlabel metal3 s 159200 75760 160000 75880 6 localMemory_wb_adr_i[13]
port 304 nsew signal input
rlabel metal3 s 159200 77256 160000 77376 6 localMemory_wb_adr_i[14]
port 305 nsew signal input
rlabel metal3 s 159200 78752 160000 78872 6 localMemory_wb_adr_i[15]
port 306 nsew signal input
rlabel metal3 s 159200 80248 160000 80368 6 localMemory_wb_adr_i[16]
port 307 nsew signal input
rlabel metal3 s 159200 81744 160000 81864 6 localMemory_wb_adr_i[17]
port 308 nsew signal input
rlabel metal3 s 159200 83240 160000 83360 6 localMemory_wb_adr_i[18]
port 309 nsew signal input
rlabel metal3 s 159200 84736 160000 84856 6 localMemory_wb_adr_i[19]
port 310 nsew signal input
rlabel metal3 s 159200 56448 160000 56568 6 localMemory_wb_adr_i[1]
port 311 nsew signal input
rlabel metal3 s 159200 86232 160000 86352 6 localMemory_wb_adr_i[20]
port 312 nsew signal input
rlabel metal3 s 159200 87728 160000 87848 6 localMemory_wb_adr_i[21]
port 313 nsew signal input
rlabel metal3 s 159200 89088 160000 89208 6 localMemory_wb_adr_i[22]
port 314 nsew signal input
rlabel metal3 s 159200 90584 160000 90704 6 localMemory_wb_adr_i[23]
port 315 nsew signal input
rlabel metal3 s 159200 58488 160000 58608 6 localMemory_wb_adr_i[2]
port 316 nsew signal input
rlabel metal3 s 159200 60392 160000 60512 6 localMemory_wb_adr_i[3]
port 317 nsew signal input
rlabel metal3 s 159200 62432 160000 62552 6 localMemory_wb_adr_i[4]
port 318 nsew signal input
rlabel metal3 s 159200 63928 160000 64048 6 localMemory_wb_adr_i[5]
port 319 nsew signal input
rlabel metal3 s 159200 65424 160000 65544 6 localMemory_wb_adr_i[6]
port 320 nsew signal input
rlabel metal3 s 159200 66920 160000 67040 6 localMemory_wb_adr_i[7]
port 321 nsew signal input
rlabel metal3 s 159200 68416 160000 68536 6 localMemory_wb_adr_i[8]
port 322 nsew signal input
rlabel metal3 s 159200 69912 160000 70032 6 localMemory_wb_adr_i[9]
port 323 nsew signal input
rlabel metal3 s 159200 52096 160000 52216 6 localMemory_wb_cyc_i
port 324 nsew signal input
rlabel metal3 s 159200 54952 160000 55072 6 localMemory_wb_data_i[0]
port 325 nsew signal input
rlabel metal3 s 159200 71816 160000 71936 6 localMemory_wb_data_i[10]
port 326 nsew signal input
rlabel metal3 s 159200 73312 160000 73432 6 localMemory_wb_data_i[11]
port 327 nsew signal input
rlabel metal3 s 159200 74808 160000 74928 6 localMemory_wb_data_i[12]
port 328 nsew signal input
rlabel metal3 s 159200 76304 160000 76424 6 localMemory_wb_data_i[13]
port 329 nsew signal input
rlabel metal3 s 159200 77800 160000 77920 6 localMemory_wb_data_i[14]
port 330 nsew signal input
rlabel metal3 s 159200 79296 160000 79416 6 localMemory_wb_data_i[15]
port 331 nsew signal input
rlabel metal3 s 159200 80792 160000 80912 6 localMemory_wb_data_i[16]
port 332 nsew signal input
rlabel metal3 s 159200 82288 160000 82408 6 localMemory_wb_data_i[17]
port 333 nsew signal input
rlabel metal3 s 159200 83648 160000 83768 6 localMemory_wb_data_i[18]
port 334 nsew signal input
rlabel metal3 s 159200 85144 160000 85264 6 localMemory_wb_data_i[19]
port 335 nsew signal input
rlabel metal3 s 159200 56992 160000 57112 6 localMemory_wb_data_i[1]
port 336 nsew signal input
rlabel metal3 s 159200 86640 160000 86760 6 localMemory_wb_data_i[20]
port 337 nsew signal input
rlabel metal3 s 159200 88136 160000 88256 6 localMemory_wb_data_i[21]
port 338 nsew signal input
rlabel metal3 s 159200 89632 160000 89752 6 localMemory_wb_data_i[22]
port 339 nsew signal input
rlabel metal3 s 159200 91128 160000 91248 6 localMemory_wb_data_i[23]
port 340 nsew signal input
rlabel metal3 s 159200 92080 160000 92200 6 localMemory_wb_data_i[24]
port 341 nsew signal input
rlabel metal3 s 159200 93168 160000 93288 6 localMemory_wb_data_i[25]
port 342 nsew signal input
rlabel metal3 s 159200 94120 160000 94240 6 localMemory_wb_data_i[26]
port 343 nsew signal input
rlabel metal3 s 159200 95072 160000 95192 6 localMemory_wb_data_i[27]
port 344 nsew signal input
rlabel metal3 s 159200 96024 160000 96144 6 localMemory_wb_data_i[28]
port 345 nsew signal input
rlabel metal3 s 159200 97112 160000 97232 6 localMemory_wb_data_i[29]
port 346 nsew signal input
rlabel metal3 s 159200 58896 160000 59016 6 localMemory_wb_data_i[2]
port 347 nsew signal input
rlabel metal3 s 159200 98064 160000 98184 6 localMemory_wb_data_i[30]
port 348 nsew signal input
rlabel metal3 s 159200 99016 160000 99136 6 localMemory_wb_data_i[31]
port 349 nsew signal input
rlabel metal3 s 159200 60936 160000 61056 6 localMemory_wb_data_i[3]
port 350 nsew signal input
rlabel metal3 s 159200 62976 160000 63096 6 localMemory_wb_data_i[4]
port 351 nsew signal input
rlabel metal3 s 159200 64472 160000 64592 6 localMemory_wb_data_i[5]
port 352 nsew signal input
rlabel metal3 s 159200 65832 160000 65952 6 localMemory_wb_data_i[6]
port 353 nsew signal input
rlabel metal3 s 159200 67328 160000 67448 6 localMemory_wb_data_i[7]
port 354 nsew signal input
rlabel metal3 s 159200 68824 160000 68944 6 localMemory_wb_data_i[8]
port 355 nsew signal input
rlabel metal3 s 159200 70320 160000 70440 6 localMemory_wb_data_i[9]
port 356 nsew signal input
rlabel metal3 s 159200 55496 160000 55616 6 localMemory_wb_data_o[0]
port 357 nsew signal output
rlabel metal3 s 159200 72360 160000 72480 6 localMemory_wb_data_o[10]
port 358 nsew signal output
rlabel metal3 s 159200 73856 160000 73976 6 localMemory_wb_data_o[11]
port 359 nsew signal output
rlabel metal3 s 159200 75352 160000 75472 6 localMemory_wb_data_o[12]
port 360 nsew signal output
rlabel metal3 s 159200 76712 160000 76832 6 localMemory_wb_data_o[13]
port 361 nsew signal output
rlabel metal3 s 159200 78208 160000 78328 6 localMemory_wb_data_o[14]
port 362 nsew signal output
rlabel metal3 s 159200 79704 160000 79824 6 localMemory_wb_data_o[15]
port 363 nsew signal output
rlabel metal3 s 159200 81200 160000 81320 6 localMemory_wb_data_o[16]
port 364 nsew signal output
rlabel metal3 s 159200 82696 160000 82816 6 localMemory_wb_data_o[17]
port 365 nsew signal output
rlabel metal3 s 159200 84192 160000 84312 6 localMemory_wb_data_o[18]
port 366 nsew signal output
rlabel metal3 s 159200 85688 160000 85808 6 localMemory_wb_data_o[19]
port 367 nsew signal output
rlabel metal3 s 159200 57536 160000 57656 6 localMemory_wb_data_o[1]
port 368 nsew signal output
rlabel metal3 s 159200 87184 160000 87304 6 localMemory_wb_data_o[20]
port 369 nsew signal output
rlabel metal3 s 159200 88680 160000 88800 6 localMemory_wb_data_o[21]
port 370 nsew signal output
rlabel metal3 s 159200 90176 160000 90296 6 localMemory_wb_data_o[22]
port 371 nsew signal output
rlabel metal3 s 159200 91672 160000 91792 6 localMemory_wb_data_o[23]
port 372 nsew signal output
rlabel metal3 s 159200 92624 160000 92744 6 localMemory_wb_data_o[24]
port 373 nsew signal output
rlabel metal3 s 159200 93576 160000 93696 6 localMemory_wb_data_o[25]
port 374 nsew signal output
rlabel metal3 s 159200 94528 160000 94648 6 localMemory_wb_data_o[26]
port 375 nsew signal output
rlabel metal3 s 159200 95616 160000 95736 6 localMemory_wb_data_o[27]
port 376 nsew signal output
rlabel metal3 s 159200 96568 160000 96688 6 localMemory_wb_data_o[28]
port 377 nsew signal output
rlabel metal3 s 159200 97520 160000 97640 6 localMemory_wb_data_o[29]
port 378 nsew signal output
rlabel metal3 s 159200 59440 160000 59560 6 localMemory_wb_data_o[2]
port 379 nsew signal output
rlabel metal3 s 159200 98608 160000 98728 6 localMemory_wb_data_o[30]
port 380 nsew signal output
rlabel metal3 s 159200 99560 160000 99680 6 localMemory_wb_data_o[31]
port 381 nsew signal output
rlabel metal3 s 159200 61480 160000 61600 6 localMemory_wb_data_o[3]
port 382 nsew signal output
rlabel metal3 s 159200 63384 160000 63504 6 localMemory_wb_data_o[4]
port 383 nsew signal output
rlabel metal3 s 159200 64880 160000 65000 6 localMemory_wb_data_o[5]
port 384 nsew signal output
rlabel metal3 s 159200 66376 160000 66496 6 localMemory_wb_data_o[6]
port 385 nsew signal output
rlabel metal3 s 159200 67872 160000 67992 6 localMemory_wb_data_o[7]
port 386 nsew signal output
rlabel metal3 s 159200 69368 160000 69488 6 localMemory_wb_data_o[8]
port 387 nsew signal output
rlabel metal3 s 159200 70864 160000 70984 6 localMemory_wb_data_o[9]
port 388 nsew signal output
rlabel metal3 s 159200 52504 160000 52624 6 localMemory_wb_error_o
port 389 nsew signal output
rlabel metal3 s 159200 56040 160000 56160 6 localMemory_wb_sel_i[0]
port 390 nsew signal input
rlabel metal3 s 159200 57944 160000 58064 6 localMemory_wb_sel_i[1]
port 391 nsew signal input
rlabel metal3 s 159200 59984 160000 60104 6 localMemory_wb_sel_i[2]
port 392 nsew signal input
rlabel metal3 s 159200 61888 160000 62008 6 localMemory_wb_sel_i[3]
port 393 nsew signal input
rlabel metal3 s 159200 53048 160000 53168 6 localMemory_wb_stall_o
port 394 nsew signal output
rlabel metal3 s 159200 53456 160000 53576 6 localMemory_wb_stb_i
port 395 nsew signal input
rlabel metal3 s 159200 54000 160000 54120 6 localMemory_wb_we_i
port 396 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 manufacturerID[0]
port 397 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 manufacturerID[10]
port 398 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 manufacturerID[1]
port 399 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 manufacturerID[2]
port 400 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 manufacturerID[3]
port 401 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 manufacturerID[4]
port 402 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 manufacturerID[5]
port 403 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 manufacturerID[6]
port 404 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 manufacturerID[7]
port 405 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 manufacturerID[8]
port 406 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 manufacturerID[9]
port 407 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 partID[0]
port 408 nsew signal input
rlabel metal2 s 120998 0 121054 800 6 partID[10]
port 409 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 partID[11]
port 410 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 partID[12]
port 411 nsew signal input
rlabel metal2 s 133234 0 133290 800 6 partID[13]
port 412 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 partID[14]
port 413 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 partID[15]
port 414 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 partID[1]
port 415 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 partID[2]
port 416 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 partID[3]
port 417 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 partID[4]
port 418 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 partID[5]
port 419 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 partID[6]
port 420 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 partID[7]
port 421 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 partID[8]
port 422 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 partID[9]
port 423 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 probe_errorCode[0]
port 424 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 probe_errorCode[1]
port 425 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 probe_errorCode[2]
port 426 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 probe_errorCode[3]
port 427 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 probe_isBranch
port 428 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 probe_isCompressed
port 429 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 probe_isLoad
port 430 nsew signal output
rlabel metal3 s 0 12656 800 12776 6 probe_isStore
port 431 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 probe_jtagInstruction[0]
port 432 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 probe_jtagInstruction[1]
port 433 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 probe_jtagInstruction[2]
port 434 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 probe_jtagInstruction[3]
port 435 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 probe_jtagInstruction[4]
port 436 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 probe_opcode[0]
port 437 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 probe_opcode[1]
port 438 nsew signal output
rlabel metal3 s 0 36320 800 36440 6 probe_opcode[2]
port 439 nsew signal output
rlabel metal3 s 0 43120 800 43240 6 probe_opcode[3]
port 440 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 probe_opcode[4]
port 441 nsew signal output
rlabel metal3 s 0 51552 800 51672 6 probe_opcode[5]
port 442 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 probe_opcode[6]
port 443 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 probe_programCounter[0]
port 444 nsew signal output
rlabel metal3 s 0 63384 800 63504 6 probe_programCounter[10]
port 445 nsew signal output
rlabel metal3 s 0 65152 800 65272 6 probe_programCounter[11]
port 446 nsew signal output
rlabel metal3 s 0 66784 800 66904 6 probe_programCounter[12]
port 447 nsew signal output
rlabel metal3 s 0 68552 800 68672 6 probe_programCounter[13]
port 448 nsew signal output
rlabel metal3 s 0 70184 800 70304 6 probe_programCounter[14]
port 449 nsew signal output
rlabel metal3 s 0 71952 800 72072 6 probe_programCounter[15]
port 450 nsew signal output
rlabel metal3 s 0 73584 800 73704 6 probe_programCounter[16]
port 451 nsew signal output
rlabel metal3 s 0 75352 800 75472 6 probe_programCounter[17]
port 452 nsew signal output
rlabel metal3 s 0 76984 800 77104 6 probe_programCounter[18]
port 453 nsew signal output
rlabel metal3 s 0 78752 800 78872 6 probe_programCounter[19]
port 454 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 probe_programCounter[1]
port 455 nsew signal output
rlabel metal3 s 0 80384 800 80504 6 probe_programCounter[20]
port 456 nsew signal output
rlabel metal3 s 0 82016 800 82136 6 probe_programCounter[21]
port 457 nsew signal output
rlabel metal3 s 0 83784 800 83904 6 probe_programCounter[22]
port 458 nsew signal output
rlabel metal3 s 0 85416 800 85536 6 probe_programCounter[23]
port 459 nsew signal output
rlabel metal3 s 0 87184 800 87304 6 probe_programCounter[24]
port 460 nsew signal output
rlabel metal3 s 0 88816 800 88936 6 probe_programCounter[25]
port 461 nsew signal output
rlabel metal3 s 0 90584 800 90704 6 probe_programCounter[26]
port 462 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 probe_programCounter[27]
port 463 nsew signal output
rlabel metal3 s 0 93984 800 94104 6 probe_programCounter[28]
port 464 nsew signal output
rlabel metal3 s 0 95616 800 95736 6 probe_programCounter[29]
port 465 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 probe_programCounter[2]
port 466 nsew signal output
rlabel metal3 s 0 97384 800 97504 6 probe_programCounter[30]
port 467 nsew signal output
rlabel metal3 s 0 99016 800 99136 6 probe_programCounter[31]
port 468 nsew signal output
rlabel metal3 s 0 44752 800 44872 6 probe_programCounter[3]
port 469 nsew signal output
rlabel metal3 s 0 49920 800 50040 6 probe_programCounter[4]
port 470 nsew signal output
rlabel metal3 s 0 53320 800 53440 6 probe_programCounter[5]
port 471 nsew signal output
rlabel metal3 s 0 56720 800 56840 6 probe_programCounter[6]
port 472 nsew signal output
rlabel metal3 s 0 58352 800 58472 6 probe_programCounter[7]
port 473 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 probe_programCounter[8]
port 474 nsew signal output
rlabel metal3 s 0 61752 800 61872 6 probe_programCounter[9]
port 475 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 probe_state[0]
port 476 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 probe_state[1]
port 477 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 probe_takeBranch
port 478 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal2 s 145562 0 145618 800 6 versionID[0]
port 480 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 versionID[1]
port 481 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 versionID[2]
port 482 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 versionID[3]
port 483 nsew signal input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal3 s 159200 144 160000 264 6 wb_clk_i
port 485 nsew signal input
rlabel metal3 s 159200 552 160000 672 6 wb_rst_i
port 486 nsew signal input
rlabel metal2 s 2870 99200 2926 100000 6 web0
port 487 nsew signal output
rlabel metal2 s 3698 99200 3754 100000 6 wmask0[0]
port 488 nsew signal output
rlabel metal2 s 4618 99200 4674 100000 6 wmask0[1]
port 489 nsew signal output
rlabel metal2 s 5446 99200 5502 100000 6 wmask0[2]
port 490 nsew signal output
rlabel metal2 s 6274 99200 6330 100000 6 wmask0[3]
port 491 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 160000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6976924
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/ExperiarCore/runs/ExperiarCore/results/signoff/ExperiarCore.magic.gds
string GDS_START 514332
<< end >>

