* NGSPICE file created from CaravelHost.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

.subckt CaravelHost caravel_uart_rx caravel_uart_tx caravel_wb_ack_i caravel_wb_adr_o[0]
+ caravel_wb_adr_o[10] caravel_wb_adr_o[11] caravel_wb_adr_o[12] caravel_wb_adr_o[13]
+ caravel_wb_adr_o[14] caravel_wb_adr_o[15] caravel_wb_adr_o[16] caravel_wb_adr_o[17]
+ caravel_wb_adr_o[18] caravel_wb_adr_o[19] caravel_wb_adr_o[1] caravel_wb_adr_o[20]
+ caravel_wb_adr_o[21] caravel_wb_adr_o[22] caravel_wb_adr_o[23] caravel_wb_adr_o[24]
+ caravel_wb_adr_o[25] caravel_wb_adr_o[26] caravel_wb_adr_o[27] caravel_wb_adr_o[2]
+ caravel_wb_adr_o[3] caravel_wb_adr_o[4] caravel_wb_adr_o[5] caravel_wb_adr_o[6]
+ caravel_wb_adr_o[7] caravel_wb_adr_o[8] caravel_wb_adr_o[9] caravel_wb_cyc_o caravel_wb_data_i[0]
+ caravel_wb_data_i[10] caravel_wb_data_i[11] caravel_wb_data_i[12] caravel_wb_data_i[13]
+ caravel_wb_data_i[14] caravel_wb_data_i[15] caravel_wb_data_i[16] caravel_wb_data_i[17]
+ caravel_wb_data_i[18] caravel_wb_data_i[19] caravel_wb_data_i[1] caravel_wb_data_i[20]
+ caravel_wb_data_i[21] caravel_wb_data_i[22] caravel_wb_data_i[23] caravel_wb_data_i[24]
+ caravel_wb_data_i[25] caravel_wb_data_i[26] caravel_wb_data_i[27] caravel_wb_data_i[28]
+ caravel_wb_data_i[29] caravel_wb_data_i[2] caravel_wb_data_i[30] caravel_wb_data_i[31]
+ caravel_wb_data_i[3] caravel_wb_data_i[4] caravel_wb_data_i[5] caravel_wb_data_i[6]
+ caravel_wb_data_i[7] caravel_wb_data_i[8] caravel_wb_data_i[9] caravel_wb_data_o[0]
+ caravel_wb_data_o[10] caravel_wb_data_o[11] caravel_wb_data_o[12] caravel_wb_data_o[13]
+ caravel_wb_data_o[14] caravel_wb_data_o[15] caravel_wb_data_o[16] caravel_wb_data_o[17]
+ caravel_wb_data_o[18] caravel_wb_data_o[19] caravel_wb_data_o[1] caravel_wb_data_o[20]
+ caravel_wb_data_o[21] caravel_wb_data_o[22] caravel_wb_data_o[23] caravel_wb_data_o[24]
+ caravel_wb_data_o[25] caravel_wb_data_o[26] caravel_wb_data_o[27] caravel_wb_data_o[28]
+ caravel_wb_data_o[29] caravel_wb_data_o[2] caravel_wb_data_o[30] caravel_wb_data_o[31]
+ caravel_wb_data_o[3] caravel_wb_data_o[4] caravel_wb_data_o[5] caravel_wb_data_o[6]
+ caravel_wb_data_o[7] caravel_wb_data_o[8] caravel_wb_data_o[9] caravel_wb_error_i
+ caravel_wb_sel_o[0] caravel_wb_sel_o[1] caravel_wb_sel_o[2] caravel_wb_sel_o[3]
+ caravel_wb_stall_i caravel_wb_stb_o caravel_wb_we_o core0Index[0] core0Index[1]
+ core0Index[2] core0Index[3] core0Index[4] core0Index[5] core0Index[6] core0Index[7]
+ core1Index[0] core1Index[1] core1Index[2] core1Index[3] core1Index[4] core1Index[5]
+ core1Index[6] core1Index[7] manufacturerID[0] manufacturerID[10] manufacturerID[1]
+ manufacturerID[2] manufacturerID[3] manufacturerID[4] manufacturerID[5] manufacturerID[6]
+ manufacturerID[7] manufacturerID[8] manufacturerID[9] partID[0] partID[10] partID[11]
+ partID[12] partID[13] partID[14] partID[15] partID[1] partID[2] partID[3] partID[4]
+ partID[5] partID[6] partID[7] partID[8] partID[9] vccd1 versionID[0] versionID[1]
+ versionID[2] versionID[3] vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_data_i[0] wbs_data_i[10] wbs_data_i[11] wbs_data_i[12] wbs_data_i[13] wbs_data_i[14]
+ wbs_data_i[15] wbs_data_i[16] wbs_data_i[17] wbs_data_i[18] wbs_data_i[19] wbs_data_i[1]
+ wbs_data_i[20] wbs_data_i[21] wbs_data_i[22] wbs_data_i[23] wbs_data_i[24] wbs_data_i[25]
+ wbs_data_i[26] wbs_data_i[27] wbs_data_i[28] wbs_data_i[29] wbs_data_i[2] wbs_data_i[30]
+ wbs_data_i[31] wbs_data_i[3] wbs_data_i[4] wbs_data_i[5] wbs_data_i[6] wbs_data_i[7]
+ wbs_data_i[8] wbs_data_i[9] wbs_data_o[0] wbs_data_o[10] wbs_data_o[11] wbs_data_o[12]
+ wbs_data_o[13] wbs_data_o[14] wbs_data_o[15] wbs_data_o[16] wbs_data_o[17] wbs_data_o[18]
+ wbs_data_o[19] wbs_data_o[1] wbs_data_o[20] wbs_data_o[21] wbs_data_o[22] wbs_data_o[23]
+ wbs_data_o[24] wbs_data_o[25] wbs_data_o[26] wbs_data_o[27] wbs_data_o[28] wbs_data_o[29]
+ wbs_data_o[2] wbs_data_o[30] wbs_data_o[31] wbs_data_o[3] wbs_data_o[4] wbs_data_o[5]
+ wbs_data_o[6] wbs_data_o[7] wbs_data_o[8] wbs_data_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
X_6465__521 _6465__521/A vssd1 vssd1 vccd1 vccd1 _7586_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6914_ _6911_/Y _6912_/X _6939_/A _6954_/A vssd1 vssd1 vccd1 vccd1 _6914_/X sky130_fd_sc_hd__a31o_1
XFILLER_23_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6845_ _6845_/A vssd1 vssd1 vccd1 vccd1 _6845_/X sky130_fd_sc_hd__buf_1
XFILLER_62_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3988_ _3988_/A vssd1 vssd1 vccd1 vccd1 _7636_/D sky130_fd_sc_hd__clkbuf_1
X_5727_ _5727_/A vssd1 vssd1 vccd1 vccd1 _6148_/S sky130_fd_sc_hd__buf_4
X_6754__141 _6757__144/A vssd1 vssd1 vccd1 vccd1 _7708_/CLK sky130_fd_sc_hd__inv_2
X_5658_ _6189_/A _5649_/X _5638_/X _7197_/Q _5639_/X vssd1 vssd1 vccd1 vccd1 _5659_/B
+ sky130_fd_sc_hd__a32o_1
X_4609_ _4609_/A vssd1 vssd1 vccd1 vccd1 _7391_/D sky130_fd_sc_hd__clkbuf_1
X_5589_ _7299_/Q _7291_/Q _7267_/Q _7115_/Q _5486_/X _5472_/X vssd1 vssd1 vccd1 vccd1
+ _5590_/B sky130_fd_sc_hd__mux4_2
X_7328_ _7329_/CLK _7328_/D vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_1
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7259_ _7259_/CLK _7259_/D vssd1 vssd1 vccd1 vccd1 _7259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3138_ clkbuf_0__3138_/X vssd1 vssd1 vccd1 vccd1 _6504__72/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6334__418 _6335__419/A vssd1 vssd1 vccd1 vccd1 _7481_/CLK sky130_fd_sc_hd__inv_2
X_6838__34 _6838__34/A vssd1 vssd1 vccd1 vccd1 _7776_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6547__106 _6548__107/A vssd1 vssd1 vccd1 vccd1 _7651_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6267__383 _6268__384/A vssd1 vssd1 vccd1 vccd1 _7436_/CLK sky130_fd_sc_hd__inv_2
X_4960_ _4960_/A vssd1 vssd1 vccd1 vccd1 _7166_/D sky130_fd_sc_hd__clkbuf_1
X_4891_ _4814_/X _7241_/Q _4893_/S vssd1 vssd1 vccd1 vccd1 _4892_/A sky130_fd_sc_hd__mux2_1
X_3911_ _3911_/A vssd1 vssd1 vccd1 vccd1 _7668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6630_ _6630_/A _6630_/B _6652_/B _6652_/C vssd1 vssd1 vccd1 vccd1 _6630_/X sky130_fd_sc_hd__or4bb_2
X_3842_ _3842_/A vssd1 vssd1 vccd1 vccd1 _7713_/D sky130_fd_sc_hd__clkbuf_1
X_6561_ _6569_/A vssd1 vssd1 vccd1 vccd1 _6621_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3773_ _3709_/X _7725_/Q _3775_/S vssd1 vssd1 vccd1 vccd1 _3774_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5512_ _5520_/A vssd1 vssd1 vccd1 vccd1 _5512_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_118_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3310_ _6820_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3310_/X sky130_fd_sc_hd__clkbuf_16
X_5443_ _5662_/A vssd1 vssd1 vccd1 vccd1 _7092_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_105_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7113_ _7113_/CLK _7113_/D vssd1 vssd1 vccd1 vccd1 _7113_/Q sky130_fd_sc_hd__dfxtp_1
X_4325_ _4155_/X _7516_/Q _4331_/S vssd1 vssd1 vccd1 vccd1 _4326_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4256_ _7825_/Q vssd1 vssd1 vccd1 vccd1 _4256_/X sky130_fd_sc_hd__buf_4
XFILLER_86_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7044_ _7044_/A vssd1 vssd1 vccd1 vccd1 _7838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4187_ _4187_/A vssd1 vssd1 vccd1 vccd1 _7558_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__2988_ clkbuf_0__2988_/X vssd1 vssd1 vccd1 vccd1 _6135__349/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5780__247 _5782__249/A vssd1 vssd1 vccd1 vccd1 _7264_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6108__327 _6108__327/A vssd1 vssd1 vccd1 vccd1 _7376_/CLK sky130_fd_sc_hd__inv_2
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5090_ _5090_/A _5098_/B vssd1 vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__and2_1
XFILLER_110_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4110_ _4150_/B _4194_/B _4865_/A vssd1 vssd1 vccd1 vccd1 _4883_/A sky130_fd_sc_hd__and3_4
XFILLER_96_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4041_ _4041_/A vssd1 vssd1 vccd1 vccd1 _7613_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5992_ _5987_/X _5991_/X _4452_/A vssd1 vssd1 vccd1 vccd1 _5992_/X sky130_fd_sc_hd__o21a_1
X_7800_ _7802_/CLK _7800_/D vssd1 vssd1 vccd1 vccd1 _7800_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__2773_ clkbuf_0__2773_/X vssd1 vssd1 vccd1 vccd1 _5813__274/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7731_ _7731_/CLK _7731_/D vssd1 vssd1 vccd1 vccd1 _7731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4943_ _4224_/X _7173_/Q _4947_/S vssd1 vssd1 vccd1 vccd1 _4944_/A sky130_fd_sc_hd__mux2_1
X_7662_ _7662_/CLK _7662_/D vssd1 vssd1 vccd1 vccd1 _7662_/Q sky130_fd_sc_hd__dfxtp_1
X_5356__188 _5357__189/A vssd1 vssd1 vccd1 vccd1 _7160_/CLK sky130_fd_sc_hd__inv_2
X_6613_ _6613_/A _6613_/B _6617_/D vssd1 vssd1 vccd1 vccd1 _6615_/A sky130_fd_sc_hd__nand3_1
X_4874_ _4874_/A vssd1 vssd1 vccd1 vccd1 _7249_/D sky130_fd_sc_hd__clkbuf_1
X_7593_ _7593_/CLK _7593_/D vssd1 vssd1 vccd1 vccd1 _7593_/Q sky130_fd_sc_hd__dfxtp_1
X_3825_ _3824_/X _7717_/Q _3829_/S vssd1 vssd1 vccd1 vccd1 _3826_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3756_ _3712_/X _7732_/Q _3756_/S vssd1 vssd1 vccd1 vccd1 _3757_/A sky130_fd_sc_hd__mux2_1
X_6544_ _6739_/A vssd1 vssd1 vccd1 vccd1 _6544_/X sky130_fd_sc_hd__buf_1
X_6475_ _6475_/A vssd1 vssd1 vccd1 vccd1 _6475_/X sky130_fd_sc_hd__buf_1
X_3687_ _3687_/A vssd1 vssd1 vccd1 vccd1 _7758_/D sky130_fd_sc_hd__clkbuf_1
X_5426_ _5426_/A vssd1 vssd1 vccd1 vccd1 _5426_/X sky130_fd_sc_hd__buf_4
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5288_ _5287_/X _7329_/Q _5283_/X _5284_/X _7129_/Q vssd1 vssd1 vccd1 vccd1 _7129_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_87_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_4 _4411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4308_ _5434_/A _4310_/B _6396_/A vssd1 vssd1 vccd1 vccd1 _4308_/Y sky130_fd_sc_hd__a21oi_1
X_7027_ _7027_/A vssd1 vssd1 vccd1 vccd1 _7827_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4239_ _7468_/Q vssd1 vssd1 vccd1 vccd1 _4239_/X sky130_fd_sc_hd__buf_2
Xclkbuf_0__3086_ _6282_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3086_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_74_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7895__222 vssd1 vssd1 vccd1 vccd1 _7895__222/HI partID[7] sky130_fd_sc_hd__conb_1
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6411__478 _6412__479/A vssd1 vssd1 vccd1 vccd1 _7543_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6735__128 _6736__129/A vssd1 vssd1 vccd1 vccd1 _7694_/CLK sky130_fd_sc_hd__inv_2
X_4590_ _7399_/Q _3944_/A _4594_/S vssd1 vssd1 vccd1 vccd1 _4591_/A sky130_fd_sc_hd__mux2_1
X_3610_ _3630_/C vssd1 vssd1 vccd1 vccd1 _4578_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3541_ _7465_/Q _7460_/Q vssd1 vssd1 vccd1 vccd1 _3541_/X sky130_fd_sc_hd__xor2_1
Xclkbuf_1_1_0__3110_ clkbuf_0__3110_/X vssd1 vssd1 vccd1 vccd1 _6363__441/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6260_ _6260_/A _6978_/A _6897_/B vssd1 vssd1 vccd1 vccd1 _6983_/A sky130_fd_sc_hd__and3_2
X_5211_ _5206_/X _5211_/B vssd1 vssd1 vccd1 vccd1 _5211_/X sky130_fd_sc_hd__and2b_1
X_6191_ _6191_/A _6866_/A _6191_/C vssd1 vssd1 vccd1 vccd1 _6253_/A sky130_fd_sc_hd__and3_1
X_5142_ _7344_/Q _5142_/B vssd1 vssd1 vccd1 vccd1 _5143_/A sky130_fd_sc_hd__and2_1
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5073_ _5073_/A _5077_/B vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__or2_1
XFILLER_57_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4024_ _3947_/X _7620_/Q _4026_/S vssd1 vssd1 vccd1 vccd1 _4025_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5975_ _7620_/Q _7612_/Q _7604_/Q _7596_/Q _5939_/X _5974_/X vssd1 vssd1 vccd1 vccd1
+ _5975_/X sky130_fd_sc_hd__mux4_2
XFILLER_40_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4926_ _4926_/A vssd1 vssd1 vccd1 vccd1 _7181_/D sky130_fd_sc_hd__clkbuf_1
X_7714_ _7714_/CLK _7714_/D vssd1 vssd1 vccd1 vccd1 _7714_/Q sky130_fd_sc_hd__dfxtp_1
X_7645_ _7645_/CLK _7645_/D vssd1 vssd1 vccd1 vccd1 _7645_/Q sky130_fd_sc_hd__dfxtp_1
X_4857_ _4817_/X _7256_/Q _4857_/S vssd1 vssd1 vccd1 vccd1 _4858_/A sky130_fd_sc_hd__mux2_1
X_7879__206 vssd1 vssd1 vccd1 vccd1 _7879__206/HI core1Index[6] sky130_fd_sc_hd__conb_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7576_ _7576_/CLK _7576_/D vssd1 vssd1 vccd1 vccd1 _7576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3808_ _7525_/Q vssd1 vssd1 vccd1 vccd1 _4111_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3308_ clkbuf_0__3308_/X vssd1 vssd1 vccd1 vccd1 _6813__14/A sky130_fd_sc_hd__clkbuf_4
X_4788_ _4788_/A vssd1 vssd1 vccd1 vccd1 _7284_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3739_ _3718_/X _7738_/Q _3741_/S vssd1 vssd1 vccd1 vccd1 _3740_/A sky130_fd_sc_hd__mux2_1
X_6499__68 _6500__69/A vssd1 vssd1 vccd1 vccd1 _7613_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5409_ _5572_/S vssd1 vssd1 vccd1 vccd1 _5432_/S sky130_fd_sc_hd__buf_4
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3138_ _6501_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3138_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _5691_/A vssd1 vssd1 vccd1 vccd1 _7207_/D sky130_fd_sc_hd__clkbuf_1
X_4711_ _4710_/X _7315_/Q _4720_/S vssd1 vssd1 vccd1 vccd1 _4712_/A sky130_fd_sc_hd__mux2_1
X_4642_ _3666_/X _7376_/Q _4642_/S vssd1 vssd1 vccd1 vccd1 _4643_/A sky130_fd_sc_hd__mux2_1
X_7430_ _7430_/CLK _7430_/D vssd1 vssd1 vccd1 vccd1 _7430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4573_ _4573_/A vssd1 vssd1 vccd1 vccd1 _7410_/D sky130_fd_sc_hd__clkbuf_1
X_7361_ _7361_/CLK _7361_/D vssd1 vssd1 vccd1 vccd1 _7361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3524_ _5462_/B _3522_/X _7405_/Q _5662_/A vssd1 vssd1 vccd1 vccd1 _3588_/A sky130_fd_sc_hd__and4bb_2
X_7292_ _7292_/CLK _7292_/D vssd1 vssd1 vccd1 vccd1 _7292_/Q sky130_fd_sc_hd__dfxtp_1
X_6312_ _6312_/A vssd1 vssd1 vccd1 vccd1 _7469_/D sky130_fd_sc_hd__clkbuf_1
X_6243_ _7846_/Q vssd1 vssd1 vccd1 vccd1 _6576_/A sky130_fd_sc_hd__inv_2
XFILLER_6_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5125_ _7336_/Q _5131_/B vssd1 vssd1 vccd1 vccd1 _5126_/A sky130_fd_sc_hd__and2_1
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5056_ _5056_/A vssd1 vssd1 vccd1 vccd1 _5056_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4007_ _3950_/X _7627_/Q _4007_/S vssd1 vssd1 vccd1 vccd1 _4008_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5958_ _6051_/A _5958_/B vssd1 vssd1 vccd1 vccd1 _5958_/X sky130_fd_sc_hd__or2_1
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4909_ _4814_/X _7233_/Q _4911_/S vssd1 vssd1 vccd1 vccd1 _4910_/A sky130_fd_sc_hd__mux2_1
X_5889_ _5889_/A vssd1 vssd1 vccd1 vccd1 _7339_/D sky130_fd_sc_hd__clkbuf_1
X_7628_ _7628_/CLK _7628_/D vssd1 vssd1 vccd1 vccd1 _7628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7559_ _7559_/CLK _7559_/D vssd1 vssd1 vccd1 vccd1 _7559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7339_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5801__264 _5801__264/A vssd1 vssd1 vccd1 vccd1 _7281_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6930_ _6930_/A _6933_/B vssd1 vssd1 vccd1 vccd1 _6930_/Y sky130_fd_sc_hd__nand2_1
X_6383__458 _6384__459/A vssd1 vssd1 vccd1 vccd1 _7521_/CLK sky130_fd_sc_hd__inv_2
X_6861_ _7841_/Q _6869_/A _6869_/B vssd1 vssd1 vccd1 vccd1 _6861_/X sky130_fd_sc_hd__and3_1
XFILLER_62_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6424__488 _6425__489/A vssd1 vssd1 vccd1 vccd1 _7553_/CLK sky130_fd_sc_hd__inv_2
X_5674_ _7202_/Q _5453_/A _5645_/A vssd1 vssd1 vccd1 vccd1 _7202_/D sky130_fd_sc_hd__a21o_1
XFILLER_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7413_ _7413_/CLK _7413_/D vssd1 vssd1 vccd1 vccd1 _7413_/Q sky130_fd_sc_hd__dfxtp_1
X_4625_ _4625_/A vssd1 vssd1 vccd1 vccd1 _7384_/D sky130_fd_sc_hd__clkbuf_1
X_7344_ _7344_/CLK _7344_/D vssd1 vssd1 vccd1 vccd1 _7344_/Q sky130_fd_sc_hd__dfxtp_1
X_4556_ _4262_/X _7417_/Q _4558_/S vssd1 vssd1 vccd1 vccd1 _4557_/A sky130_fd_sc_hd__mux2_1
X_3507_ _7464_/Q vssd1 vssd1 vccd1 vccd1 _3745_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7275_ _7275_/CLK _7275_/D vssd1 vssd1 vccd1 vccd1 _7275_/Q sky130_fd_sc_hd__dfxtp_1
X_4487_ _4937_/A _4505_/C vssd1 vssd1 vccd1 vccd1 _4503_/S sky130_fd_sc_hd__nand2_2
XFILLER_106_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6226_ _7798_/Q _6879_/A vssd1 vssd1 vccd1 vccd1 _6881_/B sky130_fd_sc_hd__xor2_2
XFILLER_106_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _5108_/A vssd1 vssd1 vccd1 vccd1 _5108_/X sky130_fd_sc_hd__clkbuf_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088_ _7728_/Q _7712_/Q _7431_/Q _7493_/Q _6024_/X _5940_/X vssd1 vssd1 vccd1 vccd1
+ _6088_/X sky130_fd_sc_hd__mux4_1
X_5039_ _5039_/A vssd1 vssd1 vccd1 vccd1 _5039_/X sky130_fd_sc_hd__clkbuf_1
X_6540__101 _6543__104/A vssd1 vssd1 vccd1 vccd1 _7646_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3085_ clkbuf_0__3085_/X vssd1 vssd1 vccd1 vccd1 _6281__394/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5744__218 _5745__219/A vssd1 vssd1 vccd1 vccd1 _7235_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput97 _5113_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[13] sky130_fd_sc_hd__buf_2
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4410_ _4410_/A vssd1 vssd1 vccd1 vccd1 _7481_/D sky130_fd_sc_hd__clkbuf_1
X_5390_ _5390_/A vssd1 vssd1 vccd1 vccd1 _5493_/B sky130_fd_sc_hd__clkbuf_1
X_4341_ _4149_/X _7509_/Q _4349_/S vssd1 vssd1 vccd1 vccd1 _4342_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7060_ _7060_/A vssd1 vssd1 vccd1 vccd1 _7106_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4272_ _4394_/A _4394_/B _4901_/C vssd1 vssd1 vccd1 vccd1 _4829_/B sky130_fd_sc_hd__and3b_2
X_6011_ _6011_/A vssd1 vssd1 vccd1 vccd1 _6011_/X sky130_fd_sc_hd__buf_2
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6913_ _7016_/A _3588_/X _5269_/A vssd1 vssd1 vccd1 vccd1 _6954_/A sky130_fd_sc_hd__a21o_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3987_ _7636_/Q _3672_/X _3989_/S vssd1 vssd1 vccd1 vccd1 _3988_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5726_ _5726_/A vssd1 vssd1 vccd1 vccd1 _7223_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5657_ _7842_/Q vssd1 vssd1 vccd1 vccd1 _6189_/A sky130_fd_sc_hd__clkbuf_4
X_4608_ _4259_/X _7391_/Q _4612_/S vssd1 vssd1 vccd1 vccd1 _4609_/A sky130_fd_sc_hd__mux2_1
X_5588_ _5466_/X _5587_/X _5403_/A vssd1 vssd1 vccd1 vccd1 _5588_/X sky130_fd_sc_hd__a21o_1
XFILLER_117_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7327_ _7329_/CLK _7327_/D vssd1 vssd1 vccd1 vccd1 _7327_/Q sky130_fd_sc_hd__dfxtp_1
X_4539_ _4265_/X _7424_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4540_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7258_ _7258_/CLK _7258_/D vssd1 vssd1 vccd1 vccd1 _7258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6209_ _7800_/Q vssd1 vssd1 vccd1 vccd1 _6933_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7189_ _7329_/CLK _7189_/D vssd1 vssd1 vccd1 vccd1 _7189_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3137_ clkbuf_0__3137_/X vssd1 vssd1 vccd1 vccd1 _6500__69/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4890_ _4890_/A vssd1 vssd1 vccd1 vccd1 _7242_/D sky130_fd_sc_hd__clkbuf_1
X_3910_ _3784_/X _7668_/Q _3918_/S vssd1 vssd1 vccd1 vccd1 _3911_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3841_ _3840_/X _7713_/Q _3841_/S vssd1 vssd1 vccd1 vccd1 _3842_/A sky130_fd_sc_hd__mux2_1
X_6560_ _7676_/Q _7675_/Q _7674_/Q _7673_/Q vssd1 vssd1 vccd1 vccd1 _6569_/A sky130_fd_sc_hd__and4_1
X_3772_ _3772_/A vssd1 vssd1 vccd1 vccd1 _7726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5511_ _5507_/X _5509_/X _5575_/S vssd1 vssd1 vccd1 vccd1 _5511_/X sky130_fd_sc_hd__mux2_1
X_5442_ _5492_/A _5672_/D _5442_/C vssd1 vssd1 vccd1 vccd1 _5442_/Y sky130_fd_sc_hd__nor3_1
XFILLER_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7112_ _7112_/CLK _7112_/D vssd1 vssd1 vccd1 vccd1 _7112_/Q sky130_fd_sc_hd__dfxtp_1
X_4324_ _4324_/A vssd1 vssd1 vccd1 vccd1 _7517_/D sky130_fd_sc_hd__clkbuf_1
X_6274__388 _6275__389/A vssd1 vssd1 vccd1 vccd1 _7441_/CLK sky130_fd_sc_hd__inv_2
X_7043_ _5680_/A _7043_/B vssd1 vssd1 vccd1 vccd1 _7044_/A sky130_fd_sc_hd__and2b_1
X_4255_ _4255_/A vssd1 vssd1 vccd1 vccd1 _7535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4186_ _4060_/X _7558_/Q _4186_/S vssd1 vssd1 vccd1 vccd1 _4187_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__2987_ clkbuf_0__2987_/X vssd1 vssd1 vccd1 vccd1 _6129__344/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6758_ _6764_/A vssd1 vssd1 vccd1 vccd1 _6758_/X sky130_fd_sc_hd__buf_1
X_5709_ _5709_/A vssd1 vssd1 vccd1 vccd1 _7215_/D sky130_fd_sc_hd__clkbuf_1
X_6689_ _6708_/A _6689_/B _6702_/C vssd1 vssd1 vccd1 vccd1 _6689_/X sky130_fd_sc_hd__or3_1
XFILLER_117_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6340__423 _6341__424/A vssd1 vssd1 vccd1 vccd1 _7486_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6553__111 _6555__113/A vssd1 vssd1 vccd1 vccd1 _7656_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4040_ _3944_/X _7613_/Q _4044_/S vssd1 vssd1 vccd1 vccd1 _4041_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5991_ _5953_/X _5988_/X _5990_/X _5959_/X vssd1 vssd1 vccd1 vccd1 _5991_/X sky130_fd_sc_hd__o211a_1
Xclkbuf_1_1_0__2772_ clkbuf_0__2772_/X vssd1 vssd1 vccd1 vccd1 _5807__269/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7730_ _7730_/CLK _7730_/D vssd1 vssd1 vccd1 vccd1 _7730_/Q sky130_fd_sc_hd__dfxtp_1
X_4942_ _4942_/A vssd1 vssd1 vccd1 vccd1 _7174_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7661_ _7661_/CLK _7661_/D vssd1 vssd1 vccd1 vccd1 _7661_/Q sky130_fd_sc_hd__dfxtp_1
X_6612_ _6612_/A _6689_/B vssd1 vssd1 vccd1 vccd1 _6612_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_60_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4873_ _7249_/Q _4405_/A _4875_/S vssd1 vssd1 vccd1 vccd1 _4874_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7592_ _7592_/CLK _7592_/D vssd1 vssd1 vccd1 vccd1 _7592_/Q sky130_fd_sc_hd__dfxtp_1
X_3824_ _4405_/A vssd1 vssd1 vccd1 vccd1 _3824_/X sky130_fd_sc_hd__buf_2
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3755_ _3755_/A vssd1 vssd1 vccd1 vccd1 _7733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3686_ _3558_/X _7758_/Q _3690_/S vssd1 vssd1 vccd1 vccd1 _3687_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5425_ _5479_/A vssd1 vssd1 vccd1 vccd1 _5426_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5287_ _5303_/A vssd1 vssd1 vccd1 vccd1 _5287_/X sky130_fd_sc_hd__buf_2
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4307_ _5433_/S _4314_/A vssd1 vssd1 vccd1 vccd1 _4310_/B sky130_fd_sc_hd__and2_1
XINSDIODE2_5 _4051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7026_ _7026_/A _7030_/B vssd1 vssd1 vccd1 vccd1 _7027_/A sky130_fd_sc_hd__and2_1
Xclkbuf_0__3085_ _6276_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3085_/X sky130_fd_sc_hd__clkbuf_16
X_4238_ _4238_/A vssd1 vssd1 vccd1 vccd1 _7540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4169_ _4169_/A vssd1 vssd1 vccd1 vccd1 _7565_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6478__532 _6478__532/A vssd1 vssd1 vccd1 vccd1 _7597_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6767__152 _6768__153/A vssd1 vssd1 vccd1 vccd1 _7719_/CLK sky130_fd_sc_hd__inv_2
X_6114__332 _6116__334/A vssd1 vssd1 vccd1 vccd1 _7381_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_39_wb_clk_i _7826_/CLK vssd1 vssd1 vccd1 vccd1 _7477_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_93_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3540_ _7464_/Q _7459_/Q vssd1 vssd1 vccd1 vccd1 _4447_/A sky130_fd_sc_hd__xor2_1
XFILLER_10_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5210_ _7137_/Q _5199_/X _5204_/X _5209_/X vssd1 vssd1 vccd1 vccd1 _5210_/X sky130_fd_sc_hd__o22a_4
X_6190_ _6869_/A _6869_/B _7841_/Q vssd1 vssd1 vccd1 vccd1 _6191_/C sky130_fd_sc_hd__a21bo_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5141_ _5141_/A vssd1 vssd1 vccd1 vccd1 _5141_/X sky130_fd_sc_hd__clkbuf_1
X_5072_ _5072_/A vssd1 vssd1 vccd1 vccd1 _5072_/X sky130_fd_sc_hd__clkbuf_1
X_5362__193 _5362__193/A vssd1 vssd1 vccd1 vccd1 _7165_/CLK sky130_fd_sc_hd__inv_2
X_4023_ _4023_/A vssd1 vssd1 vccd1 vccd1 _7621_/D sky130_fd_sc_hd__clkbuf_1
X_6347__429 _6347__429/A vssd1 vssd1 vccd1 vccd1 _7492_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5974_ _5998_/A vssd1 vssd1 vccd1 vccd1 _5974_/X sky130_fd_sc_hd__clkbuf_4
X_7713_ _7713_/CLK _7713_/D vssd1 vssd1 vccd1 vccd1 _7713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4925_ _4224_/X _7181_/Q _4929_/S vssd1 vssd1 vccd1 vccd1 _4926_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7644_ _7644_/CLK _7644_/D vssd1 vssd1 vccd1 vccd1 _7644_/Q sky130_fd_sc_hd__dfxtp_1
X_4856_ _4856_/A vssd1 vssd1 vccd1 vccd1 _7257_/D sky130_fd_sc_hd__clkbuf_1
X_5926__320 _5929__323/A vssd1 vssd1 vccd1 vccd1 _7361_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3807_ _4194_/A _4194_/B _4686_/A vssd1 vssd1 vccd1 vccd1 _4901_/D sky130_fd_sc_hd__nand3_2
X_7575_ _7575_/CLK _7575_/D vssd1 vssd1 vccd1 vccd1 _7575_/Q sky130_fd_sc_hd__dfxtp_1
X_6526_ _6538_/A vssd1 vssd1 vccd1 vccd1 _6526_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3307_ clkbuf_0__3307_/X vssd1 vssd1 vccd1 vccd1 _6803__5/A sky130_fd_sc_hd__clkbuf_4
X_4787_ _4705_/X _7284_/Q _4795_/S vssd1 vssd1 vccd1 vccd1 _4788_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3738_ _3738_/A vssd1 vssd1 vccd1 vccd1 _7739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3669_ _7824_/Q vssd1 vssd1 vccd1 vccd1 _3669_/X sky130_fd_sc_hd__buf_4
X_6457_ _6475_/A vssd1 vssd1 vccd1 vccd1 _6457_/X sky130_fd_sc_hd__buf_1
X_5408_ _5516_/A vssd1 vssd1 vccd1 vccd1 _5572_/S sky130_fd_sc_hd__clkbuf_4
X_5339_ _5307_/A _5317_/B _7060_/A vssd1 vssd1 vccd1 vccd1 _7228_/D sky130_fd_sc_hd__a21oi_1
XFILLER_48_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3137_ _6495_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3137_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_102_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7009_ _6996_/A _6997_/A _7819_/Q vssd1 vssd1 vccd1 vccd1 _7009_/X sky130_fd_sc_hd__a21o_1
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5793__258 _5794__259/A vssd1 vssd1 vccd1 vccd1 _7275_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _7207_/Q _5094_/A _5692_/S vssd1 vssd1 vccd1 vccd1 _5691_/A sky130_fd_sc_hd__mux2_1
X_4710_ _7474_/Q vssd1 vssd1 vccd1 vccd1 _4710_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4641_ _4641_/A vssd1 vssd1 vccd1 vccd1 _7377_/D sky130_fd_sc_hd__clkbuf_1
X_4572_ _4259_/X _7410_/Q _4576_/S vssd1 vssd1 vccd1 vccd1 _4573_/A sky130_fd_sc_hd__mux2_1
X_7360_ _7360_/CLK _7360_/D vssd1 vssd1 vccd1 vccd1 _7360_/Q sky130_fd_sc_hd__dfxtp_1
X_3523_ _7227_/Q _5679_/B vssd1 vssd1 vccd1 vccd1 _5662_/A sky130_fd_sc_hd__and2b_1
X_7291_ _7291_/CLK _7291_/D vssd1 vssd1 vccd1 vccd1 _7291_/Q sky130_fd_sc_hd__dfxtp_1
X_6311_ _7815_/Q _6319_/B vssd1 vssd1 vccd1 vccd1 _6312_/A sky130_fd_sc_hd__and2_1
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6242_ _6242_/A _6889_/B vssd1 vssd1 vccd1 vccd1 _6866_/B sky130_fd_sc_hd__xor2_1
XFILLER_103_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6173_ _6263_/A vssd1 vssd1 vccd1 vccd1 _6173_/X sky130_fd_sc_hd__buf_1
X_5124_ _5124_/A vssd1 vssd1 vccd1 vccd1 _5124_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5055_ _5055_/A _5055_/B vssd1 vssd1 vccd1 vccd1 _5056_/A sky130_fd_sc_hd__or2_1
XFILLER_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4006_ _4006_/A vssd1 vssd1 vccd1 vccd1 _7628_/D sky130_fd_sc_hd__clkbuf_1
X_6810__11 _6812__13/A vssd1 vssd1 vccd1 vccd1 _7753_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5957_ _7587_/Q _7555_/Q _7830_/Q _7531_/Q _6002_/A _5956_/X vssd1 vssd1 vccd1 vccd1
+ _5958_/B sky130_fd_sc_hd__mux4_1
XFILLER_52_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4908_ _4908_/A vssd1 vssd1 vccd1 vccd1 _7234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5888_ _5062_/A _7339_/Q _5890_/S vssd1 vssd1 vccd1 vccd1 _5889_/A sky130_fd_sc_hd__mux2_1
X_7627_ _7627_/CLK _7627_/D vssd1 vssd1 vccd1 vccd1 _7627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4839_ _4817_/X _7264_/Q _4839_/S vssd1 vssd1 vccd1 vccd1 _4840_/A sky130_fd_sc_hd__mux2_1
X_7558_ _7558_/CLK _7558_/D vssd1 vssd1 vccd1 vccd1 _7558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7489_ _7489_/CLK _7489_/D vssd1 vssd1 vccd1 vccd1 _7489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5369__199 _5369__199/A vssd1 vssd1 vccd1 vccd1 _7171_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3299_ clkbuf_0__3299_/X vssd1 vssd1 vccd1 vccd1 _6768__153/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6860_ _6869_/A _6869_/B _5661_/X vssd1 vssd1 vccd1 vccd1 _6860_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6127__342 _6127__342/A vssd1 vssd1 vccd1 vccd1 _7391_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5673_ _7201_/Q _5453_/A _5645_/A _5672_/X vssd1 vssd1 vccd1 vccd1 _7201_/D sky130_fd_sc_hd__a211o_1
XFILLER_30_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7412_ _7412_/CLK _7412_/D vssd1 vssd1 vccd1 vccd1 _7412_/Q sky130_fd_sc_hd__dfxtp_1
X_4624_ _3666_/X _7384_/Q _4624_/S vssd1 vssd1 vccd1 vccd1 _4625_/A sky130_fd_sc_hd__mux2_1
X_7343_ _7344_/CLK _7343_/D vssd1 vssd1 vccd1 vccd1 _7343_/Q sky130_fd_sc_hd__dfxtp_1
X_4555_ _4555_/A vssd1 vssd1 vccd1 vccd1 _7418_/D sky130_fd_sc_hd__clkbuf_1
X_3506_ _7466_/Q vssd1 vssd1 vccd1 vccd1 _4009_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7274_ _7274_/CLK _7274_/D vssd1 vssd1 vccd1 vccd1 _7274_/Q sky130_fd_sc_hd__dfxtp_1
X_4486_ _4486_/A vssd1 vssd1 vccd1 vccd1 _7449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6225_ _6218_/X _6219_/Y _6222_/Y _6223_/Y _6224_/X vssd1 vssd1 vccd1 vccd1 _6225_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_97_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5107_/A _5109_/B vssd1 vssd1 vccd1 vccd1 _5108_/A sky130_fd_sc_hd__and2_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6644__115 _6645__116/A vssd1 vssd1 vccd1 vccd1 _7662_/CLK sky130_fd_sc_hd__inv_2
X_6087_ _7371_/Q _6631_/B _6086_/X _5996_/A vssd1 vssd1 vccd1 vccd1 _7371_/D sky130_fd_sc_hd__o211a_1
X_5038_ _5038_/A _5044_/B vssd1 vssd1 vccd1 vccd1 _5039_/A sky130_fd_sc_hd__or2_1
XFILLER_38_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6989_ _6195_/A _6195_/B _6873_/B _6872_/A vssd1 vssd1 vccd1 vccd1 _6989_/X sky130_fd_sc_hd__o22a_1
XFILLER_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3084_ clkbuf_0__3084_/X vssd1 vssd1 vccd1 vccd1 _6273__387/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput98 _5115_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[14] sky130_fd_sc_hd__buf_2
XFILLER_110_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4340_ _4355_/S vssd1 vssd1 vccd1 vccd1 _4349_/S sky130_fd_sc_hd__buf_2
XFILLER_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4271_ _4271_/A _4285_/B vssd1 vssd1 vccd1 vccd1 _4278_/B sky130_fd_sc_hd__nand2_1
XFILLER_113_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6010_ _6005_/X _6006_/X _6009_/X _5959_/A vssd1 vssd1 vccd1 vccd1 _6010_/X sky130_fd_sc_hd__o211a_1
XFILLER_79_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6430__493 _6431__494/A vssd1 vssd1 vccd1 vccd1 _7558_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6912_ _6943_/A vssd1 vssd1 vccd1 vccd1 _6912_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3986_ _3986_/A vssd1 vssd1 vccd1 vccd1 _7637_/D sky130_fd_sc_hd__clkbuf_1
X_5725_ _7223_/Q _7338_/Q _5725_/S vssd1 vssd1 vccd1 vccd1 _5726_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5656_ _5656_/A vssd1 vssd1 vccd1 vccd1 _7196_/D sky130_fd_sc_hd__clkbuf_1
X_4607_ _4607_/A vssd1 vssd1 vccd1 vccd1 _7392_/D sky130_fd_sc_hd__clkbuf_1
X_6472__527 _6474__529/A vssd1 vssd1 vccd1 vccd1 _7592_/CLK sky130_fd_sc_hd__inv_2
X_5587_ _7307_/Q _7235_/Q _7703_/Q _7323_/Q _4296_/A _4302_/B vssd1 vssd1 vccd1 vccd1
+ _5587_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7326_ _7329_/CLK _7326_/D vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dfxtp_1
X_4538_ _4538_/A vssd1 vssd1 vccd1 vccd1 _7425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7257_ _7257_/CLK _7257_/D vssd1 vssd1 vccd1 vccd1 _7257_/Q sky130_fd_sc_hd__dfxtp_1
X_4469_ _4901_/D _4706_/A vssd1 vssd1 vccd1 vccd1 _4485_/S sky130_fd_sc_hd__or2_2
XFILLER_104_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6208_ _6991_/A _6208_/B _6991_/B vssd1 vssd1 vccd1 vccd1 _6238_/B sky130_fd_sc_hd__and3_1
X_7188_ _7839_/CLK _7188_/D vssd1 vssd1 vccd1 vccd1 _7188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6761__147 _6763__149/A vssd1 vssd1 vccd1 vccd1 _7714_/CLK sky130_fd_sc_hd__inv_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5750__223 _5751__224/A vssd1 vssd1 vccd1 vccd1 _7240_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3136_ clkbuf_0__3136_/X vssd1 vssd1 vccd1 vccd1 _6492__62/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3840_ _4417_/A vssd1 vssd1 vccd1 vccd1 _3840_/X sky130_fd_sc_hd__buf_2
X_3771_ _3706_/X _7726_/Q _3775_/S vssd1 vssd1 vccd1 vccd1 _3772_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5510_ _5516_/A vssd1 vssd1 vccd1 vccd1 _5575_/S sky130_fd_sc_hd__buf_4
XFILLER_118_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5920__315 _5920__315/A vssd1 vssd1 vccd1 vccd1 _7356_/CLK sky130_fd_sc_hd__inv_2
X_5441_ _5423_/Y _5434_/Y _6396_/B _5440_/X vssd1 vssd1 vccd1 vccd1 _5442_/C sky130_fd_sc_hd__o31a_1
XFILLER_113_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4323_ _4149_/X _7517_/Q _4331_/S vssd1 vssd1 vccd1 vccd1 _4324_/A sky130_fd_sc_hd__mux2_1
X_7111_ _7111_/CLK _7111_/D vssd1 vssd1 vccd1 vccd1 _7111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7042_ _5051_/A _6394_/A _7045_/S vssd1 vssd1 vccd1 vccd1 _7043_/B sky130_fd_sc_hd__mux2_1
X_6844__39 _6844__39/A vssd1 vssd1 vccd1 vccd1 _7781_/CLK sky130_fd_sc_hd__inv_2
X_4254_ _4253_/X _7535_/Q _4257_/S vssd1 vssd1 vccd1 vccd1 _4255_/A sky130_fd_sc_hd__mux2_1
X_4185_ _4185_/A vssd1 vssd1 vccd1 vccd1 _7559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__2986_ clkbuf_0__2986_/X vssd1 vssd1 vccd1 vccd1 _6123__339/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6826_ _6826_/A vssd1 vssd1 vccd1 vccd1 _6826_/X sky130_fd_sc_hd__buf_1
XFILLER_50_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5708_ _7215_/Q _5112_/A _5714_/S vssd1 vssd1 vccd1 vccd1 _5709_/A sky130_fd_sc_hd__mux2_1
X_3969_ _3969_/A vssd1 vssd1 vccd1 vccd1 _7644_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6688_ _6640_/C _6661_/X _6610_/Y vssd1 vssd1 vccd1 vccd1 _6688_/X sky130_fd_sc_hd__a21o_1
X_5639_ _5662_/A vssd1 vssd1 vccd1 vccd1 _5639_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6437__499 _6437__499/A vssd1 vssd1 vccd1 vccd1 _7564_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7309_ _7309_/CLK _7309_/D vssd1 vssd1 vccd1 vccd1 _7309_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3299_ _6764_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3299_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_86_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3119_ clkbuf_0__3119_/X vssd1 vssd1 vccd1 vccd1 _6412__479/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5757__229 _5757__229/A vssd1 vssd1 vccd1 vccd1 _7246_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5990_ _6051_/A _5990_/B vssd1 vssd1 vccd1 vccd1 _5990_/X sky130_fd_sc_hd__or2_1
XFILLER_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__2771_ clkbuf_0__2771_/X vssd1 vssd1 vccd1 vccd1 _5799__262/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4941_ _4221_/X _7174_/Q _4947_/S vssd1 vssd1 vccd1 vccd1 _4942_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7660_ _7684_/CLK _7660_/D vssd1 vssd1 vccd1 vccd1 _7660_/Q sky130_fd_sc_hd__dfxtp_1
X_4872_ _4872_/A vssd1 vssd1 vccd1 vccd1 _7250_/D sky130_fd_sc_hd__clkbuf_1
X_6611_ _6602_/B _6613_/B _6593_/A _6610_/Y vssd1 vssd1 vccd1 vccd1 _6689_/B sky130_fd_sc_hd__a22o_1
X_3823_ _7472_/Q vssd1 vssd1 vccd1 vccd1 _4405_/A sky130_fd_sc_hd__clkbuf_2
X_7591_ _7591_/CLK _7591_/D vssd1 vssd1 vccd1 vccd1 _7591_/Q sky130_fd_sc_hd__dfxtp_1
X_6280__393 _6281__394/A vssd1 vssd1 vccd1 vccd1 _7446_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_9_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7407_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3754_ _3709_/X _7733_/Q _3756_/S vssd1 vssd1 vccd1 vccd1 _3755_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3685_ _3685_/A vssd1 vssd1 vccd1 vccd1 _7759_/D sky130_fd_sc_hd__clkbuf_1
X_5424_ _7661_/Q _7494_/Q _7449_/Q _7309_/Q _5413_/X _5416_/X vssd1 vssd1 vccd1 vccd1
+ _5424_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5355_ _6725_/B _5350_/X _6677_/A _6690_/A vssd1 vssd1 vccd1 vccd1 _7159_/D sky130_fd_sc_hd__a211o_1
XFILLER_114_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6817__17 _6818__18/A vssd1 vssd1 vccd1 vccd1 _7759_/CLK sky130_fd_sc_hd__inv_2
X_5286_ _5278_/X hold4/X _5283_/X _5284_/X _7128_/Q vssd1 vssd1 vccd1 vccd1 _7128_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4306_ _5613_/A _4312_/A _4312_/B vssd1 vssd1 vccd1 vccd1 _4314_/A sky130_fd_sc_hd__and3_1
XINSDIODE2_6 _4057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7025_ _7025_/A vssd1 vssd1 vccd1 vccd1 _7826_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3084_ _6270_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3084_/X sky130_fd_sc_hd__clkbuf_16
X_4237_ _7540_/Q _4236_/X _4240_/S vssd1 vssd1 vccd1 vccd1 _4238_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4168_ _4167_/X _7565_/Q _4174_/S vssd1 vssd1 vccd1 vccd1 _4169_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4099_ _4099_/A vssd1 vssd1 vccd1 vccd1 _7591_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7789_ _7789_/CLK _7789_/D vssd1 vssd1 vccd1 vccd1 _7789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6774__157 _6776__159/A vssd1 vssd1 vccd1 vccd1 _7724_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6160__364 _6160__364/A vssd1 vssd1 vccd1 vccd1 _7416_/CLK sky130_fd_sc_hd__inv_2
X_6121__337 _6123__339/A vssd1 vssd1 vccd1 vccd1 _7386_/CLK sky130_fd_sc_hd__inv_2
X_5140_ _7343_/Q _5142_/B vssd1 vssd1 vccd1 vccd1 _5141_/A sky130_fd_sc_hd__and2_1
XFILLER_111_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5071_ _5071_/A _5077_/B vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__or2_1
X_4022_ _3944_/X _7621_/Q _4026_/S vssd1 vssd1 vccd1 vccd1 _4023_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5973_ _7754_/Q _7746_/Q _7738_/Q _7652_/Q _4465_/A _5937_/X vssd1 vssd1 vccd1 vccd1
+ _5973_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7712_ _7712_/CLK _7712_/D vssd1 vssd1 vccd1 vccd1 _7712_/Q sky130_fd_sc_hd__dfxtp_1
X_4924_ _4924_/A vssd1 vssd1 vccd1 vccd1 _7182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7643_ _7643_/CLK _7643_/D vssd1 vssd1 vccd1 vccd1 _7643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4855_ _4814_/X _7257_/Q _4857_/S vssd1 vssd1 vccd1 vccd1 _4856_/A sky130_fd_sc_hd__mux2_1
X_3806_ _7096_/A _3588_/A _5239_/A vssd1 vssd1 vccd1 vccd1 _4686_/A sky130_fd_sc_hd__a21oi_2
X_7574_ _7574_/CLK _7574_/D vssd1 vssd1 vccd1 vccd1 _7574_/Q sky130_fd_sc_hd__dfxtp_1
X_4786_ _4801_/S vssd1 vssd1 vccd1 vccd1 _4795_/S sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__3306_ clkbuf_0__3306_/X vssd1 vssd1 vccd1 vccd1 _6826_/A sky130_fd_sc_hd__clkbuf_4
X_3737_ _3715_/X _7739_/Q _3741_/S vssd1 vssd1 vccd1 vccd1 _3738_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3668_ _3668_/A vssd1 vssd1 vccd1 vccd1 _7764_/D sky130_fd_sc_hd__clkbuf_1
X_3599_ _3599_/A vssd1 vssd1 vccd1 vccd1 _7790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5407_ _7520_/Q vssd1 vssd1 vccd1 vccd1 _5516_/A sky130_fd_sc_hd__inv_2
XFILLER_102_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5338_ _5338_/A vssd1 vssd1 vccd1 vccd1 _7060_/A sky130_fd_sc_hd__buf_2
XFILLER_87_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3136_ _6489_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3136_/X sky130_fd_sc_hd__clkbuf_16
X_5269_ _5269_/A vssd1 vssd1 vccd1 vccd1 _5303_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7008_ _7819_/Q _6995_/X _7007_/X _7003_/X vssd1 vssd1 vccd1 vccd1 _7818_/D sky130_fd_sc_hd__o211a_1
XFILLER_75_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6287__399 _6287__399/A vssd1 vssd1 vccd1 vccd1 _7452_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6307__414 _6307__414/A vssd1 vssd1 vccd1 vccd1 _7467_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4640_ _3663_/X _7377_/Q _4642_/S vssd1 vssd1 vccd1 vccd1 _4641_/A sky130_fd_sc_hd__mux2_1
X_4571_ _4571_/A vssd1 vssd1 vccd1 vccd1 _7411_/D sky130_fd_sc_hd__clkbuf_1
X_6310_ _6310_/A vssd1 vssd1 vccd1 vccd1 _6319_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3522_ _7205_/Q _5390_/A _7204_/Q vssd1 vssd1 vccd1 vccd1 _3522_/X sky130_fd_sc_hd__or3b_1
X_7290_ _7290_/CLK _7290_/D vssd1 vssd1 vccd1 vccd1 _7290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6241_ _6193_/B _6241_/B vssd1 vssd1 vccd1 vccd1 _6889_/B sky130_fd_sc_hd__nand2b_2
X_6353__434 _6353__434/A vssd1 vssd1 vccd1 vccd1 _7497_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5123_ _7335_/Q _5131_/B vssd1 vssd1 vccd1 vccd1 _5124_/A sky130_fd_sc_hd__and2_1
XFILLER_111_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _5054_/A vssd1 vssd1 vccd1 vccd1 _5054_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7885__212 vssd1 vssd1 vccd1 vccd1 _7885__212/HI manufacturerID[4] sky130_fd_sc_hd__conb_1
X_4005_ _3947_/X _7628_/Q _4007_/S vssd1 vssd1 vccd1 vccd1 _4006_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5956_ _6024_/A vssd1 vssd1 vccd1 vccd1 _5956_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_53_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5887_ _5887_/A vssd1 vssd1 vccd1 vccd1 _7338_/D sky130_fd_sc_hd__clkbuf_1
X_4907_ _4811_/X _7234_/Q _4911_/S vssd1 vssd1 vccd1 vccd1 _4908_/A sky130_fd_sc_hd__mux2_1
X_4838_ _4838_/A vssd1 vssd1 vccd1 vccd1 _7265_/D sky130_fd_sc_hd__clkbuf_1
X_7626_ _7626_/CLK _7626_/D vssd1 vssd1 vccd1 vccd1 _7626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7557_ _7557_/CLK _7557_/D vssd1 vssd1 vccd1 vccd1 _7557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4769_ _4705_/X _7292_/Q _4777_/S vssd1 vssd1 vccd1 vccd1 _4770_/A sky130_fd_sc_hd__mux2_1
X_7488_ _7488_/CLK _7488_/D vssd1 vssd1 vccd1 vccd1 _7488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__3119_ _6407_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3119_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_29_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3298_ clkbuf_0__3298_/X vssd1 vssd1 vccd1 vccd1 _6763__149/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_23_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7845_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_82_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7411_ _7411_/CLK _7411_/D vssd1 vssd1 vccd1 vccd1 _7411_/Q sky130_fd_sc_hd__dfxtp_1
X_5672_ _6394_/A _5679_/A _7407_/Q _5672_/D vssd1 vssd1 vccd1 vccd1 _5672_/X sky130_fd_sc_hd__and4_1
X_4623_ _4623_/A vssd1 vssd1 vccd1 vccd1 _7385_/D sky130_fd_sc_hd__clkbuf_1
X_7342_ _7344_/CLK _7342_/D vssd1 vssd1 vccd1 vccd1 _7342_/Q sky130_fd_sc_hd__dfxtp_1
X_4554_ _4259_/X _7418_/Q _4558_/S vssd1 vssd1 vccd1 vccd1 _4555_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3505_ _3926_/A vssd1 vssd1 vccd1 vccd1 _3505_/X sky130_fd_sc_hd__clkbuf_2
X_7273_ _7273_/CLK _7273_/D vssd1 vssd1 vccd1 vccd1 _7273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6224_ _7855_/Q _6911_/A vssd1 vssd1 vccd1 vccd1 _6224_/X sky130_fd_sc_hd__or2_1
X_4485_ _4417_/X _7449_/Q _4485_/S vssd1 vssd1 vccd1 vccd1 _4486_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6155_ _6167_/A vssd1 vssd1 vccd1 vccd1 _6155_/X sky130_fd_sc_hd__buf_1
XFILLER_58_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5106_/A vssd1 vssd1 vccd1 vccd1 _5106_/X sky130_fd_sc_hd__clkbuf_1
X_6086_ _5932_/A _6076_/X _6085_/X _5993_/A vssd1 vssd1 vccd1 vccd1 _6086_/X sky130_fd_sc_hd__a211o_2
XFILLER_85_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5037_ _5037_/A vssd1 vssd1 vccd1 vccd1 _5037_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6988_ _6235_/Y _6236_/X _6987_/Y _6229_/X _6225_/X vssd1 vssd1 vccd1 vccd1 _6993_/B
+ sky130_fd_sc_hd__o2111a_1
Xclkbuf_1_0_0__3083_ clkbuf_0__3083_/X vssd1 vssd1 vccd1 vccd1 _6282_/A sky130_fd_sc_hd__clkbuf_4
X_5939_ _6024_/A vssd1 vssd1 vccd1 vccd1 _5939_/X sky130_fd_sc_hd__buf_4
XFILLER_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7609_ _7609_/CLK _7609_/D vssd1 vssd1 vccd1 vccd1 _7609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput99 _5117_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[15] sky130_fd_sc_hd__buf_2
XFILLER_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__3296_ clkbuf_0__3296_/X vssd1 vssd1 vccd1 vccd1 _6749__137/A sky130_fd_sc_hd__clkbuf_16
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4270_ _4285_/B _4270_/B vssd1 vssd1 vccd1 vccd1 _7528_/D sky130_fd_sc_hd__nor2_1
XFILLER_4_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6911_ _6911_/A vssd1 vssd1 vccd1 vccd1 _6911_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3985_ _7637_/Q _3669_/X _3989_/S vssd1 vssd1 vccd1 vccd1 _3986_/A sky130_fd_sc_hd__mux2_1
X_5724_ _5724_/A vssd1 vssd1 vccd1 vccd1 _7222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5655_ _5667_/A _5655_/B vssd1 vssd1 vccd1 vccd1 _5656_/A sky130_fd_sc_hd__or2_1
X_4606_ _4256_/X _7392_/Q _4606_/S vssd1 vssd1 vccd1 vccd1 _4607_/A sky130_fd_sc_hd__mux2_1
X_7325_ _7331_/CLK _7325_/D vssd1 vssd1 vccd1 vccd1 _7325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5586_ _5590_/A _5586_/B vssd1 vssd1 vccd1 vccd1 _5586_/X sky130_fd_sc_hd__and2_1
X_6650__120 _6651__121/A vssd1 vssd1 vccd1 vccd1 _7667_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4537_ _4262_/X _7425_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4538_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4468_ _4468_/A vssd1 vssd1 vccd1 vccd1 _7457_/D sky130_fd_sc_hd__clkbuf_1
X_7256_ _7256_/CLK _7256_/D vssd1 vssd1 vccd1 vccd1 _7256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7187_ _7407_/CLK _7187_/D vssd1 vssd1 vccd1 vccd1 _7187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6207_ _6605_/A _6883_/A _6883_/B vssd1 vssd1 vccd1 vccd1 _6991_/B sky130_fd_sc_hd__nand3_1
XFILLER_112_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4399_ _4399_/A vssd1 vssd1 vccd1 vccd1 _4399_/X sky130_fd_sc_hd__buf_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _6064_/X _6068_/X _6036_/X vssd1 vssd1 vccd1 vccd1 _6069_/X sky130_fd_sc_hd__o21a_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6366__444 _6366__444/A vssd1 vssd1 vccd1 vccd1 _7507_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3135_ clkbuf_0__3135_/X vssd1 vssd1 vccd1 vccd1 _6486__57/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3770_ _3770_/A vssd1 vssd1 vccd1 vccd1 _7727_/D sky130_fd_sc_hd__clkbuf_1
X_5440_ _5462_/A _7040_/B _5493_/B _5462_/D vssd1 vssd1 vccd1 vccd1 _5440_/X sky130_fd_sc_hd__or4_1
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4322_ _4337_/S vssd1 vssd1 vccd1 vccd1 _4331_/S sky130_fd_sc_hd__buf_2
X_7110_ _7110_/CLK _7110_/D vssd1 vssd1 vccd1 vccd1 _7110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4253_ _7826_/Q vssd1 vssd1 vccd1 vccd1 _4253_/X sky130_fd_sc_hd__buf_4
X_7041_ _7407_/Q _7077_/B vssd1 vssd1 vccd1 vccd1 _7045_/S sky130_fd_sc_hd__nand2_1
XFILLER_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4184_ _4057_/X _7559_/Q _4186_/S vssd1 vssd1 vccd1 vccd1 _4185_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__2985_ clkbuf_0__2985_/X vssd1 vssd1 vccd1 vccd1 _6142_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3968_ _3947_/X _7644_/Q _3970_/S vssd1 vssd1 vccd1 vccd1 _3969_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5707_ _5707_/A vssd1 vssd1 vccd1 vccd1 _7214_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6687_ _6685_/X _6686_/X _6665_/X vssd1 vssd1 vccd1 vccd1 _7675_/D sky130_fd_sc_hd__a21oi_1
X_3899_ _3828_/X _7691_/Q _3899_/S vssd1 vssd1 vccd1 vccd1 _3900_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5638_ _5638_/A vssd1 vssd1 vccd1 vccd1 _5638_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5569_ _5567_/X _5568_/X _5569_/S vssd1 vssd1 vccd1 vccd1 _5569_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7308_ _7308_/CLK _7308_/D vssd1 vssd1 vccd1 vccd1 _7308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7239_ _7239_/CLK _7239_/D vssd1 vssd1 vccd1 vccd1 _7239_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3298_ _6758_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3298_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3118_ clkbuf_0__3118_/X vssd1 vssd1 vccd1 vccd1 _6406__474/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6531__94 _6531__94/A vssd1 vssd1 vccd1 vccd1 _7639_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__2770_ clkbuf_0__2770_/X vssd1 vssd1 vccd1 vccd1 _5820_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4940_ _4940_/A vssd1 vssd1 vccd1 vccd1 _7175_/D sky130_fd_sc_hd__clkbuf_1
X_4871_ _7250_/Q _4402_/A _4875_/S vssd1 vssd1 vccd1 vccd1 _4872_/A sky130_fd_sc_hd__mux2_1
X_6610_ _7676_/Q vssd1 vssd1 vccd1 vccd1 _6610_/Y sky130_fd_sc_hd__inv_2
X_7590_ _7590_/CLK _7590_/D vssd1 vssd1 vccd1 vccd1 _7590_/Q sky130_fd_sc_hd__dfxtp_1
X_3822_ _3822_/A vssd1 vssd1 vccd1 vccd1 _7718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3753_ _3753_/A vssd1 vssd1 vccd1 vccd1 _7734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3684_ _3554_/X _7759_/Q _3690_/S vssd1 vssd1 vccd1 vccd1 _3685_/A sky130_fd_sc_hd__mux2_1
X_5423_ _5404_/X _5410_/X _5422_/X vssd1 vssd1 vccd1 vccd1 _5423_/Y sky130_fd_sc_hd__a21oi_1
X_5354_ _7100_/A _3588_/X _7060_/A vssd1 vssd1 vccd1 vccd1 _6690_/A sky130_fd_sc_hd__a21o_2
X_4305_ _4305_/A _7530_/Q _5396_/A vssd1 vssd1 vccd1 vccd1 _4312_/B sky130_fd_sc_hd__and3_1
X_5285_ _5278_/X _7327_/Q _5283_/X _5284_/X _7127_/Q vssd1 vssd1 vccd1 vccd1 _7127_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_59_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_7 _4224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7024_ _7024_/A _7024_/B vssd1 vssd1 vccd1 vccd1 _7025_/A sky130_fd_sc_hd__and2_1
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4236_ _7469_/Q vssd1 vssd1 vccd1 vccd1 _4236_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3083_ _6269_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3083_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_101_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4167_ _4411_/A vssd1 vssd1 vccd1 vccd1 _4167_/X sky130_fd_sc_hd__buf_2
XFILLER_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4098_ _4057_/X _7591_/Q _4100_/S vssd1 vssd1 vccd1 vccd1 _4099_/A sky130_fd_sc_hd__mux2_1
X_5374__203 _5374__203/A vssd1 vssd1 vccd1 vccd1 _7175_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6808_ _6814_/A vssd1 vssd1 vccd1 vccd1 _6808_/X sky130_fd_sc_hd__buf_1
X_7788_ _7788_/CLK _7788_/D vssd1 vssd1 vccd1 vccd1 _7788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6739_ _6739_/A vssd1 vssd1 vccd1 vccd1 _6739_/X sky130_fd_sc_hd__buf_1
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5763__234 _5763__234/A vssd1 vssd1 vccd1 vccd1 _7251_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6504__72 _6504__72/A vssd1 vssd1 vccd1 vccd1 _7617_/CLK sky130_fd_sc_hd__inv_2
X_5070_ _5070_/A vssd1 vssd1 vccd1 vccd1 _5070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4021_ _4021_/A vssd1 vssd1 vccd1 vccd1 _7622_/D sky130_fd_sc_hd__clkbuf_1
X_6822__21 _6822__21/A vssd1 vssd1 vccd1 vccd1 _7763_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5972_ _7722_/Q _7706_/Q _7425_/Q _7487_/Q _5933_/X _4457_/A vssd1 vssd1 vccd1 vccd1
+ _5972_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7711_ _7711_/CLK _7711_/D vssd1 vssd1 vccd1 vccd1 _7711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4923_ _4221_/X _7182_/Q _4929_/S vssd1 vssd1 vccd1 vccd1 _4924_/A sky130_fd_sc_hd__mux2_1
X_7642_ _7642_/CLK _7642_/D vssd1 vssd1 vccd1 vccd1 _7642_/Q sky130_fd_sc_hd__dfxtp_1
X_4854_ _4854_/A vssd1 vssd1 vccd1 vccd1 _7258_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3805_ _3805_/A vssd1 vssd1 vccd1 vccd1 _7096_/A sky130_fd_sc_hd__buf_6
X_4785_ _4901_/D _4955_/B vssd1 vssd1 vccd1 vccd1 _4801_/S sky130_fd_sc_hd__or2_4
X_7573_ _7573_/CLK _7573_/D vssd1 vssd1 vccd1 vccd1 _7573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3736_ _3736_/A vssd1 vssd1 vccd1 vccd1 _7740_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3305_ clkbuf_0__3305_/X vssd1 vssd1 vccd1 vccd1 _6800__179/A sky130_fd_sc_hd__clkbuf_4
XFILLER_119_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3667_ _7764_/Q _3666_/X _3667_/S vssd1 vssd1 vccd1 vccd1 _3668_/A sky130_fd_sc_hd__mux2_1
X_3598_ _3558_/X _7790_/Q _3602_/S vssd1 vssd1 vccd1 vccd1 _3599_/A sky130_fd_sc_hd__mux2_1
X_6386_ _6392_/A vssd1 vssd1 vccd1 vccd1 _6386_/X sky130_fd_sc_hd__buf_1
X_5406_ _7176_/Q _7357_/Q _7713_/Q _7253_/Q _4305_/A _4312_/A vssd1 vssd1 vccd1 vccd1
+ _5406_/X sky130_fd_sc_hd__mux4_1
X_5337_ _5239_/A _5337_/B _5337_/C vssd1 vssd1 vccd1 vccd1 _5682_/C sky130_fd_sc_hd__and3b_2
X_5268_ _5245_/B _7150_/Q _5262_/X _5266_/X _7118_/Q vssd1 vssd1 vccd1 vccd1 _7118_/D
+ sky130_fd_sc_hd__o32a_1
Xclkbuf_0__3135_ _6483_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3135_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4219_ _7546_/Q _4213_/X _4231_/S vssd1 vssd1 vccd1 vccd1 _4220_/A sky130_fd_sc_hd__mux2_1
X_7007_ _6996_/X _6997_/X _7818_/Q vssd1 vssd1 vccd1 vccd1 _7007_/X sky130_fd_sc_hd__a21o_1
X_5199_ _5199_/A vssd1 vssd1 vccd1 vccd1 _5199_/X sky130_fd_sc_hd__buf_2
XFILLER_18_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6780__162 _6782__164/A vssd1 vssd1 vccd1 vccd1 _7729_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4570_ _4256_/X _7411_/Q _4570_/S vssd1 vssd1 vccd1 vccd1 _4571_/A sky130_fd_sc_hd__mux2_1
X_3521_ _5458_/C _5458_/D vssd1 vssd1 vccd1 vccd1 _5390_/A sky130_fd_sc_hd__or2_1
XFILLER_116_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6240_ _7805_/Q _6245_/A _6245_/B _6245_/C _7806_/Q vssd1 vssd1 vccd1 vccd1 _6241_/B
+ sky130_fd_sc_hd__a41o_1
X_5122_ _5122_/A vssd1 vssd1 vccd1 vccd1 _5131_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5053_ _5053_/A _5055_/B vssd1 vssd1 vccd1 vccd1 _5054_/A sky130_fd_sc_hd__or2_1
XFILLER_38_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4004_ _4004_/A vssd1 vssd1 vccd1 vccd1 _7629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5955_ _7785_/Q _7777_/Q _7769_/Q _7761_/Q _4446_/A _5954_/X vssd1 vssd1 vccd1 vccd1
+ _5955_/X sky130_fd_sc_hd__mux4_1
X_6360__439 _6360__439/A vssd1 vssd1 vccd1 vccd1 _7502_/CLK sky130_fd_sc_hd__inv_2
X_5886_ _5060_/A _7338_/Q _5890_/S vssd1 vssd1 vccd1 vccd1 _5887_/A sky130_fd_sc_hd__mux2_1
X_4906_ _4906_/A vssd1 vssd1 vccd1 vccd1 _7235_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4837_ _4814_/X _7265_/Q _4839_/S vssd1 vssd1 vccd1 vccd1 _4838_/A sky130_fd_sc_hd__mux2_1
X_7625_ _7625_/CLK _7625_/D vssd1 vssd1 vccd1 vccd1 _7625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7556_ _7556_/CLK _7556_/D vssd1 vssd1 vccd1 vccd1 _7556_/Q sky130_fd_sc_hd__dfxtp_1
X_4768_ _4783_/S vssd1 vssd1 vccd1 vccd1 _4777_/S sky130_fd_sc_hd__buf_2
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3719_ _3718_/X _7746_/Q _3722_/S vssd1 vssd1 vccd1 vccd1 _3720_/A sky130_fd_sc_hd__mux2_1
X_7487_ _7487_/CLK _7487_/D vssd1 vssd1 vccd1 vccd1 _7487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4699_ _4411_/X _7319_/Q _4703_/S vssd1 vssd1 vccd1 vccd1 _4700_/A sky130_fd_sc_hd__mux2_1
X_6507_ _6507_/A vssd1 vssd1 vccd1 vccd1 _6507_/X sky130_fd_sc_hd__buf_1
X_6438_ _6444_/A vssd1 vssd1 vccd1 vccd1 _6438_/X sky130_fd_sc_hd__buf_1
XFILLER_20_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3118_ _6401_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3118_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3297_ clkbuf_0__3297_/X vssd1 vssd1 vccd1 vccd1 _6757__144/A sky130_fd_sc_hd__clkbuf_4
XFILLER_12_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5740_ _5740_/A vssd1 vssd1 vccd1 vccd1 _5740_/X sky130_fd_sc_hd__buf_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7410_ _7410_/CLK _7410_/D vssd1 vssd1 vccd1 vccd1 _7410_/Q sky130_fd_sc_hd__dfxtp_1
X_5671_ _7838_/Q vssd1 vssd1 vccd1 vccd1 _6394_/A sky130_fd_sc_hd__clkbuf_4
X_4622_ _3663_/X _7385_/Q _4624_/S vssd1 vssd1 vccd1 vccd1 _4623_/A sky130_fd_sc_hd__mux2_1
X_7341_ _7344_/CLK _7341_/D vssd1 vssd1 vccd1 vccd1 _7341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4553_ _4553_/A vssd1 vssd1 vccd1 vccd1 _7419_/D sky130_fd_sc_hd__clkbuf_1
X_3504_ _7829_/Q vssd1 vssd1 vccd1 vccd1 _3926_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7272_ _7272_/CLK _7272_/D vssd1 vssd1 vccd1 vccd1 _7272_/Q sky130_fd_sc_hd__dfxtp_1
X_4484_ _4484_/A vssd1 vssd1 vccd1 vccd1 _7450_/D sky130_fd_sc_hd__clkbuf_1
X_6787__168 _6787__168/A vssd1 vssd1 vccd1 vccd1 _7735_/CLK sky130_fd_sc_hd__inv_2
X_6223_ _7855_/Q _6911_/A vssd1 vssd1 vccd1 vccd1 _6223_/Y sky130_fd_sc_hd__nand2_1
X_6134__348 _6135__349/A vssd1 vssd1 vccd1 vccd1 _7397_/CLK sky130_fd_sc_hd__inv_2
X_6154_ _6269_/A vssd1 vssd1 vccd1 vccd1 _6154_/X sky130_fd_sc_hd__buf_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5105_/A _5109_/B vssd1 vssd1 vccd1 vccd1 _5106_/A sky130_fd_sc_hd__and2_1
X_6085_ _6080_/X _6084_/X _6036_/X vssd1 vssd1 vccd1 vccd1 _6085_/X sky130_fd_sc_hd__o21a_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5776__244 _5776__244/A vssd1 vssd1 vccd1 vccd1 _7261_/CLK sky130_fd_sc_hd__inv_2
X_5036_ _5036_/A _5044_/B vssd1 vssd1 vccd1 vccd1 _5037_/A sky130_fd_sc_hd__or2_1
XFILLER_57_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6442__503 _6442__503/A vssd1 vssd1 vccd1 vccd1 _7568_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6987_ _6195_/A _6195_/B _6208_/B vssd1 vssd1 vccd1 vccd1 _6987_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5938_ _7753_/Q _7745_/Q _7737_/Q _7651_/Q _5935_/X _5937_/X vssd1 vssd1 vccd1 vccd1
+ _5938_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3082_ clkbuf_0__3082_/X vssd1 vssd1 vccd1 vccd1 _6268__384/A sky130_fd_sc_hd__clkbuf_4
X_5869_ _5869_/A vssd1 vssd1 vccd1 vccd1 _7330_/D sky130_fd_sc_hd__clkbuf_1
X_6399__468 _6400__469/A vssd1 vssd1 vccd1 vccd1 _7533_/CLK sky130_fd_sc_hd__inv_2
X_7608_ _7608_/CLK _7608_/D vssd1 vssd1 vccd1 vccd1 _7608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7539_ _7539_/CLK _7539_/D vssd1 vssd1 vccd1 vccd1 _7539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6856__49 _6856__49/A vssd1 vssd1 vccd1 vccd1 _7791_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6910_ _6902_/S _6900_/Y _6908_/X _6909_/X vssd1 vssd1 vccd1 vccd1 _7794_/D sky130_fd_sc_hd__o211a_1
XFILLER_50_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3984_ _3984_/A vssd1 vssd1 vccd1 vccd1 _7638_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5723_ _7222_/Q _7337_/Q _5725_/S vssd1 vssd1 vccd1 vccd1 _5724_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5654_ _6195_/A _5649_/X _5638_/X _7196_/Q _5639_/X vssd1 vssd1 vccd1 vccd1 _5655_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4605_ _4605_/A vssd1 vssd1 vccd1 vccd1 _7393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5585_ _7667_/Q _7500_/Q _7455_/Q _7315_/Q _5427_/A _5472_/X vssd1 vssd1 vccd1 vccd1
+ _5586_/B sky130_fd_sc_hd__mux4_1
X_7324_ _7324_/CLK _7324_/D vssd1 vssd1 vccd1 vccd1 _7324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4536_ _4536_/A vssd1 vssd1 vccd1 vccd1 _7426_/D sky130_fd_sc_hd__clkbuf_1
X_4467_ _4457_/B _4467_/B _6328_/B vssd1 vssd1 vccd1 vccd1 _4468_/A sky130_fd_sc_hd__and3b_1
X_7255_ _7255_/CLK _7255_/D vssd1 vssd1 vccd1 vccd1 _7255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7186_ _7839_/CLK _7186_/D vssd1 vssd1 vccd1 vccd1 _7186_/Q sky130_fd_sc_hd__dfxtp_1
X_6206_ _6231_/A _6231_/B _6612_/A vssd1 vssd1 vccd1 vccd1 _6208_/B sky130_fd_sc_hd__a21o_1
X_4398_ _4398_/A vssd1 vssd1 vccd1 vccd1 _7485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6068_ _6005_/X _6065_/X _6067_/X _5959_/X vssd1 vssd1 vccd1 vccd1 _6068_/X sky130_fd_sc_hd__o211a_1
XFILLER_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5019_ _5019_/A vssd1 vssd1 vccd1 vccd1 _5019_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3134_ clkbuf_0__3134_/X vssd1 vssd1 vccd1 vccd1 _6507_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6449__509 _6449__509/A vssd1 vssd1 vccd1 vccd1 _7574_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7870__197 vssd1 vssd1 vccd1 vccd1 _7870__197/HI core0Index[4] sky130_fd_sc_hd__conb_1
XFILLER_91_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5370_ _5376_/A vssd1 vssd1 vccd1 vccd1 _5370_/X sky130_fd_sc_hd__buf_1
X_6829__27 _6831__29/A vssd1 vssd1 vccd1 vccd1 _7769_/CLK sky130_fd_sc_hd__inv_2
X_4321_ _4883_/A _4505_/C vssd1 vssd1 vccd1 vccd1 _4337_/S sky130_fd_sc_hd__nand2_4
XFILLER_99_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4252_ _4252_/A vssd1 vssd1 vccd1 vccd1 _7536_/D sky130_fd_sc_hd__clkbuf_1
X_7040_ _7040_/A _7040_/B _7040_/C vssd1 vssd1 vccd1 vccd1 _7077_/B sky130_fd_sc_hd__nor3_2
XFILLER_86_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4183_ _4183_/A vssd1 vssd1 vccd1 vccd1 _7560_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__2984_ clkbuf_0__2984_/X vssd1 vssd1 vccd1 vccd1 _6113__331/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3967_ _3967_/A vssd1 vssd1 vccd1 vccd1 _7645_/D sky130_fd_sc_hd__clkbuf_1
X_5706_ _7214_/Q _5109_/A _5714_/S vssd1 vssd1 vccd1 vccd1 _5707_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6686_ _6708_/A _6686_/B _6702_/C vssd1 vssd1 vccd1 vccd1 _6686_/X sky130_fd_sc_hd__or3_1
X_3898_ _3898_/A vssd1 vssd1 vccd1 vccd1 _7692_/D sky130_fd_sc_hd__clkbuf_1
X_5637_ _5679_/A _7406_/Q vssd1 vssd1 vccd1 vccd1 _5638_/A sky130_fd_sc_hd__and2_1
X_6292__403 _6292__403/A vssd1 vssd1 vccd1 vccd1 _7456_/CLK sky130_fd_sc_hd__inv_2
X_5568_ _7306_/Q _7234_/Q _7702_/Q _7322_/Q _5426_/A _5518_/X vssd1 vssd1 vccd1 vccd1
+ _5568_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7307_ _7307_/CLK _7307_/D vssd1 vssd1 vccd1 vccd1 _7307_/Q sky130_fd_sc_hd__dfxtp_1
X_4519_ _7434_/Q _4236_/X _4521_/S vssd1 vssd1 vccd1 vccd1 _4520_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5499_ _7185_/Q _5453_/X _5498_/X vssd1 vssd1 vccd1 vccd1 _7185_/D sky130_fd_sc_hd__a21o_1
X_7238_ _7238_/CLK _7238_/D vssd1 vssd1 vccd1 vccd1 _7238_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3297_ _6752_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3297_/X sky130_fd_sc_hd__clkbuf_16
X_7169_ _7169_/CLK _7169_/D vssd1 vssd1 vccd1 vccd1 _7169_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6455__513 _6455__513/A vssd1 vssd1 vccd1 vccd1 _7578_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6516__81 _6516__81/A vssd1 vssd1 vccd1 vccd1 _7626_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6834__30 _6836__32/A vssd1 vssd1 vccd1 vccd1 _7772_/CLK sky130_fd_sc_hd__inv_2
X_6744__133 _6745__134/A vssd1 vssd1 vccd1 vccd1 _7700_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4870_ _4870_/A vssd1 vssd1 vccd1 vccd1 _7251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3821_ _3820_/X _7718_/Q _3829_/S vssd1 vssd1 vccd1 vccd1 _3822_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3752_ _3706_/X _7734_/Q _3756_/S vssd1 vssd1 vccd1 vccd1 _3753_/A sky130_fd_sc_hd__mux2_1
X_3683_ _3683_/A vssd1 vssd1 vccd1 vccd1 _7760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5422_ _5433_/S _5420_/X _5421_/Y vssd1 vssd1 vccd1 vccd1 _5422_/X sky130_fd_sc_hd__a21o_1
X_5353_ _6714_/A vssd1 vssd1 vccd1 vccd1 _6677_/A sky130_fd_sc_hd__buf_2
X_4304_ _4302_/X _4304_/B _4304_/C vssd1 vssd1 vccd1 vccd1 _5396_/A sky130_fd_sc_hd__nand3b_2
X_5284_ _5284_/A vssd1 vssd1 vccd1 vccd1 _5284_/X sky130_fd_sc_hd__clkbuf_2
X_7023_ _7023_/A vssd1 vssd1 vccd1 vccd1 _7825_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_8 _4224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0__3082_ _6263_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3082_/X sky130_fd_sc_hd__clkbuf_16
X_4235_ _4235_/A vssd1 vssd1 vccd1 vccd1 _7541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4166_ _4166_/A vssd1 vssd1 vccd1 vccd1 _7566_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4097_ _4097_/A vssd1 vssd1 vccd1 vccd1 _7592_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4999_ _4999_/A vssd1 vssd1 vccd1 vccd1 _4999_/X sky130_fd_sc_hd__clkbuf_1
X_7787_ _7787_/CLK _7787_/D vssd1 vssd1 vccd1 vccd1 _7787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6738_ _6738_/A vssd1 vssd1 vccd1 vccd1 _7696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6669_ _6705_/A vssd1 vssd1 vccd1 vccd1 _6711_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6299__409 _6299__409/A vssd1 vssd1 vccd1 vccd1 _7462_/CLK sky130_fd_sc_hd__inv_2
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7344_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4020_ _3941_/X _7622_/Q _4020_/S vssd1 vssd1 vccd1 vccd1 _4021_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5770__239 _5770__239/A vssd1 vssd1 vccd1 vccd1 _7256_/CLK sky130_fd_sc_hd__inv_2
X_5971_ _7365_/Q _5931_/X _5967_/X _5970_/X vssd1 vssd1 vccd1 vccd1 _7365_/D sky130_fd_sc_hd__o211a_1
XFILLER_80_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7710_ _7710_/CLK _7710_/D vssd1 vssd1 vccd1 vccd1 _7710_/Q sky130_fd_sc_hd__dfxtp_1
X_4922_ _4922_/A vssd1 vssd1 vccd1 vccd1 _7183_/D sky130_fd_sc_hd__clkbuf_1
X_7641_ _7641_/CLK _7641_/D vssd1 vssd1 vccd1 vccd1 _7641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4853_ _4811_/X _7258_/Q _4857_/S vssd1 vssd1 vccd1 vccd1 _4854_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3804_ _4285_/A _3865_/A vssd1 vssd1 vccd1 vccd1 _4194_/B sky130_fd_sc_hd__and2b_1
X_7572_ _7572_/CLK _7572_/D vssd1 vssd1 vccd1 vccd1 _7572_/Q sky130_fd_sc_hd__dfxtp_1
X_4784_ _4784_/A vssd1 vssd1 vccd1 vccd1 _7285_/D sky130_fd_sc_hd__clkbuf_1
X_3735_ _3712_/X _7740_/Q _3735_/S vssd1 vssd1 vccd1 vccd1 _3736_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3304_ clkbuf_0__3304_/X vssd1 vssd1 vccd1 vccd1 _6792__172/A sky130_fd_sc_hd__clkbuf_4
XFILLER_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3666_ _7825_/Q vssd1 vssd1 vccd1 vccd1 _3666_/X sky130_fd_sc_hd__clkbuf_4
X_5405_ _7579_/Q _7563_/Q _7547_/Q _7539_/Q _4305_/A _4312_/A vssd1 vssd1 vccd1 vccd1
+ _5405_/X sky130_fd_sc_hd__mux4_1
X_3597_ _3597_/A vssd1 vssd1 vccd1 vccd1 _7791_/D sky130_fd_sc_hd__clkbuf_1
X_6385_ _6385_/A vssd1 vssd1 vccd1 vccd1 _6385_/X sky130_fd_sc_hd__buf_1
X_5336_ _7158_/Q _4998_/A _7157_/Q vssd1 vssd1 vccd1 vccd1 _5336_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5267_ _5245_/B _7149_/Q _5262_/X _5266_/X _7117_/Q vssd1 vssd1 vccd1 vccd1 _7117_/D
+ sky130_fd_sc_hd__o32a_1
Xclkbuf_0__3134_ _6482_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3134_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_102_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4218_ _4240_/S vssd1 vssd1 vccd1 vccd1 _4231_/S sky130_fd_sc_hd__clkbuf_2
X_7006_ _7818_/Q _6995_/X _7005_/X _7003_/X vssd1 vssd1 vccd1 vccd1 _7817_/D sky130_fd_sc_hd__o211a_1
X_5198_ _5198_/A vssd1 vssd1 vccd1 vccd1 _5199_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4149_ _4393_/A vssd1 vssd1 vccd1 vccd1 _4149_/X sky130_fd_sc_hd__buf_2
XFILLER_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7862__236 vssd1 vssd1 vccd1 vccd1 partID[10] _7862__236/LO sky130_fd_sc_hd__conb_1
X_7839_ _7839_/CLK _7839_/D vssd1 vssd1 vccd1 vccd1 _7839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3520_ _5399_/C _3520_/B vssd1 vssd1 vccd1 vccd1 _5458_/D sky130_fd_sc_hd__or2_2
XFILLER_115_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5121_ _5121_/A vssd1 vssd1 vccd1 vccd1 _5121_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5052_ _5052_/A vssd1 vssd1 vccd1 vccd1 _5052_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4003_ _3944_/X _7629_/Q _4007_/S vssd1 vssd1 vccd1 vccd1 _4004_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5954_ _6011_/A vssd1 vssd1 vccd1 vccd1 _5954_/X sky130_fd_sc_hd__clkbuf_4
X_5885_ _5885_/A vssd1 vssd1 vccd1 vccd1 _7337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4905_ _4808_/X _7235_/Q _4911_/S vssd1 vssd1 vccd1 vccd1 _4906_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4836_ _4836_/A vssd1 vssd1 vccd1 vccd1 _7266_/D sky130_fd_sc_hd__clkbuf_1
X_7624_ _7624_/CLK _7624_/D vssd1 vssd1 vccd1 vccd1 _7624_/Q sky130_fd_sc_hd__dfxtp_1
X_7555_ _7555_/CLK _7555_/D vssd1 vssd1 vccd1 vccd1 _7555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4767_ _4767_/A _4829_/B vssd1 vssd1 vccd1 vccd1 _4783_/S sky130_fd_sc_hd__nand2_4
X_3718_ _3947_/A vssd1 vssd1 vccd1 vccd1 _3718_/X sky130_fd_sc_hd__clkbuf_2
X_7486_ _7486_/CLK _7486_/D vssd1 vssd1 vccd1 vccd1 _7486_/Q sky130_fd_sc_hd__dfxtp_1
X_4698_ _4698_/A vssd1 vssd1 vccd1 vccd1 _7320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3649_ _7829_/Q vssd1 vssd1 vccd1 vccd1 _3649_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_114_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5319_ _5334_/S vssd1 vssd1 vccd1 vccd1 _5328_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5670_ _7200_/Q _5453_/A _5645_/A _5669_/X vssd1 vssd1 vccd1 vccd1 _7200_/D sky130_fd_sc_hd__a211o_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_32_wb_clk_i _7474_/CLK vssd1 vssd1 vccd1 vccd1 _7808_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1_0__2451_ clkbuf_0__2451_/X vssd1 vssd1 vccd1 vccd1 _5740_/A sky130_fd_sc_hd__clkbuf_4
X_4621_ _4621_/A vssd1 vssd1 vccd1 vccd1 _7386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7340_ _7344_/CLK _7340_/D vssd1 vssd1 vccd1 vccd1 _7340_/Q sky130_fd_sc_hd__dfxtp_2
X_4552_ _4256_/X _7419_/Q _4552_/S vssd1 vssd1 vccd1 vccd1 _4553_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7271_ _7271_/CLK _7271_/D vssd1 vssd1 vccd1 vccd1 _7271_/Q sky130_fd_sc_hd__dfxtp_1
X_4483_ _4414_/X _7450_/Q _4485_/S vssd1 vssd1 vccd1 vccd1 _4484_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6222_ _6918_/A _6222_/B vssd1 vssd1 vccd1 vccd1 _6222_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_112_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _5104_/A vssd1 vssd1 vccd1 vccd1 _5104_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6084_ _6005_/X _6081_/X _6083_/X _5959_/X vssd1 vssd1 vccd1 vccd1 _6084_/X sky130_fd_sc_hd__o211a_1
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5081_/B vssd1 vssd1 vccd1 vccd1 _5044_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6986_ _6986_/A vssd1 vssd1 vccd1 vccd1 _7813_/D sky130_fd_sc_hd__clkbuf_1
X_5937_ _6011_/A vssd1 vssd1 vccd1 vccd1 _5937_/X sky130_fd_sc_hd__buf_4
XFILLER_53_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5868_ _5042_/A _7330_/Q _5872_/S vssd1 vssd1 vccd1 vccd1 _5869_/A sky130_fd_sc_hd__mux2_1
X_7607_ _7607_/CLK _7607_/D vssd1 vssd1 vccd1 vccd1 _7607_/Q sky130_fd_sc_hd__dfxtp_1
X_4819_ _4819_/A vssd1 vssd1 vccd1 vccd1 _7272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7538_ _7538_/CLK _7538_/D vssd1 vssd1 vccd1 vccd1 _7538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7469_ _7818_/CLK _7469_/D vssd1 vssd1 vccd1 vccd1 _7469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7875__202 vssd1 vssd1 vccd1 vccd1 _7875__202/HI core1Index[2] sky130_fd_sc_hd__conb_1
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6771_ _6783_/A vssd1 vssd1 vccd1 vccd1 _6771_/X sky130_fd_sc_hd__buf_1
XFILLER_62_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5722_ _5722_/A vssd1 vssd1 vccd1 vccd1 _7221_/D sky130_fd_sc_hd__clkbuf_1
X_3983_ _7638_/Q _3666_/X _3983_/S vssd1 vssd1 vccd1 vccd1 _3984_/A sky130_fd_sc_hd__mux2_1
X_6793__173 _6794__174/A vssd1 vssd1 vccd1 vccd1 _7740_/CLK sky130_fd_sc_hd__inv_2
X_5653_ _7843_/Q vssd1 vssd1 vccd1 vccd1 _6195_/A sky130_fd_sc_hd__buf_2
X_6140__353 _6141__354/A vssd1 vssd1 vccd1 vccd1 _7402_/CLK sky130_fd_sc_hd__inv_2
X_4604_ _4253_/X _7393_/Q _4606_/S vssd1 vssd1 vccd1 vccd1 _4605_/A sky130_fd_sc_hd__mux2_1
X_5584_ _7849_/Q vssd1 vssd1 vccd1 vccd1 _5584_/X sky130_fd_sc_hd__clkbuf_4
X_4535_ _4259_/X _7426_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4536_/A sky130_fd_sc_hd__mux2_1
X_7323_ _7323_/CLK _7323_/D vssd1 vssd1 vccd1 vccd1 _7323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4466_ _7477_/Q _6328_/C _4465_/X vssd1 vssd1 vccd1 vccd1 _4467_/B sky130_fd_sc_hd__a21o_1
X_7254_ _7254_/CLK _7254_/D vssd1 vssd1 vccd1 vccd1 _7254_/Q sky130_fd_sc_hd__dfxtp_1
X_7185_ _7839_/CLK _7185_/D vssd1 vssd1 vccd1 vccd1 _7185_/Q sky130_fd_sc_hd__dfxtp_1
X_6205_ _7848_/Q vssd1 vssd1 vccd1 vccd1 _6612_/A sky130_fd_sc_hd__inv_2
X_4397_ _4393_/X _7485_/Q _4409_/S vssd1 vssd1 vccd1 vccd1 _4398_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6136_ _6142_/A vssd1 vssd1 vccd1 vccd1 _6136_/X sky130_fd_sc_hd__buf_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6067_ _6099_/A _6067_/B vssd1 vssd1 vccd1 vccd1 _6067_/X sky130_fd_sc_hd__or2_1
X_5018_ _7096_/A _5022_/B vssd1 vssd1 vccd1 vccd1 _5019_/A sky130_fd_sc_hd__or2_1
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3133_ clkbuf_0__3133_/X vssd1 vssd1 vccd1 vccd1 _6739_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6969_ _7810_/Q _6969_/B vssd1 vssd1 vccd1 vccd1 _6969_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6156__360 _6158__362/A vssd1 vssd1 vccd1 vccd1 _7412_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2779_ clkbuf_0__2779_/X vssd1 vssd1 vccd1 vccd1 _5839__294/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4320_ _4901_/C _4394_/B _4394_/A vssd1 vssd1 vccd1 vccd1 _4505_/C sky130_fd_sc_hd__and3b_4
X_4251_ _4250_/X _7536_/Q _4257_/S vssd1 vssd1 vccd1 vccd1 _4252_/A sky130_fd_sc_hd__mux2_1
X_4182_ _4054_/X _7560_/Q _4186_/S vssd1 vssd1 vccd1 vccd1 _4183_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__2983_ clkbuf_0__2983_/X vssd1 vssd1 vccd1 vccd1 _6110__329/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3966_ _3944_/X _7645_/Q _3970_/S vssd1 vssd1 vccd1 vccd1 _3967_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5705_ _5727_/A vssd1 vssd1 vccd1 vccd1 _5714_/S sky130_fd_sc_hd__clkbuf_2
X_6685_ _6679_/X _6684_/X _7675_/Q vssd1 vssd1 vccd1 vccd1 _6685_/X sky130_fd_sc_hd__a21bo_1
XFILLER_10_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5636_ _5647_/A vssd1 vssd1 vccd1 vccd1 _5645_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3897_ _3824_/X _7692_/Q _3899_/S vssd1 vssd1 vccd1 vccd1 _3898_/A sky130_fd_sc_hd__mux2_1
X_5567_ _7666_/Q _7499_/Q _7454_/Q _7314_/Q _5502_/X _5416_/A vssd1 vssd1 vccd1 vccd1
+ _5567_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5498_ _5455_/X _5460_/X _5496_/X _5497_/X vssd1 vssd1 vccd1 vccd1 _5498_/X sky130_fd_sc_hd__a31o_1
XFILLER_2_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7306_ _7306_/CLK _7306_/D vssd1 vssd1 vccd1 vccd1 _7306_/Q sky130_fd_sc_hd__dfxtp_1
X_4518_ _4518_/A vssd1 vssd1 vccd1 vccd1 _7435_/D sky130_fd_sc_hd__clkbuf_1
X_4449_ _4449_/A vssd1 vssd1 vccd1 vccd1 _6328_/C sky130_fd_sc_hd__buf_2
X_7237_ _7237_/CLK _7237_/D vssd1 vssd1 vccd1 vccd1 _7237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3296_ _6746_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3296_/X sky130_fd_sc_hd__clkbuf_16
X_7168_ _7168_/CLK _7168_/D vssd1 vssd1 vccd1 vccd1 _7168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7099_ _7104_/B _7854_/Q vssd1 vssd1 vccd1 vccd1 _7101_/B sky130_fd_sc_hd__and2b_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3116_ clkbuf_0__3116_/X vssd1 vssd1 vccd1 vccd1 _6400__469/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6349__430 _6349__430/A vssd1 vssd1 vccd1 vccd1 _7493_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__2777_ clkbuf_0__2777_/X vssd1 vssd1 vccd1 vccd1 _5840_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_94_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3820_ _4402_/A vssd1 vssd1 vccd1 vccd1 _3820_/X sky130_fd_sc_hd__buf_2
X_3751_ _3751_/A vssd1 vssd1 vccd1 vccd1 _7735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3682_ _3505_/X _7760_/Q _3690_/S vssd1 vssd1 vccd1 vccd1 _3683_/A sky130_fd_sc_hd__mux2_1
X_5421_ _7522_/Q vssd1 vssd1 vccd1 vccd1 _5421_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5352_ _5949_/B vssd1 vssd1 vccd1 vccd1 _6714_/A sky130_fd_sc_hd__buf_2
X_4303_ _3796_/X _4303_/B _4303_/C _4303_/D vssd1 vssd1 vccd1 vccd1 _4304_/C sky130_fd_sc_hd__and4b_1
XFILLER_114_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5283_ _5307_/A vssd1 vssd1 vccd1 vccd1 _5283_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7022_ _7092_/A _7024_/B vssd1 vssd1 vccd1 vccd1 _7023_/A sky130_fd_sc_hd__and2_1
XINSDIODE2_9 _4230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4234_ _7541_/Q _4233_/X _4240_/S vssd1 vssd1 vccd1 vccd1 _4235_/A sky130_fd_sc_hd__mux2_1
X_4165_ _4164_/X _7566_/Q _4165_/S vssd1 vssd1 vccd1 vccd1 _4166_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4096_ _4054_/X _7592_/Q _4100_/S vssd1 vssd1 vccd1 vccd1 _4097_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7855_ _7855_/CLK _7855_/D vssd1 vssd1 vccd1 vccd1 _7855_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4998_ _4998_/A _5002_/B vssd1 vssd1 vccd1 vccd1 _4999_/A sky130_fd_sc_hd__and2_1
X_7786_ _7786_/CLK _7786_/D vssd1 vssd1 vccd1 vccd1 _7786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3949_ _3949_/A vssd1 vssd1 vccd1 vccd1 _7652_/D sky130_fd_sc_hd__clkbuf_1
X_6737_ _7696_/Q _5950_/A _6737_/S vssd1 vssd1 vccd1 vccd1 _6738_/A sky130_fd_sc_hd__mux2_1
X_6668_ _6725_/B _6668_/B vssd1 vssd1 vccd1 vccd1 _6705_/A sky130_fd_sc_hd__or2_1
X_6599_ _6598_/Y _6670_/B _6602_/B vssd1 vssd1 vccd1 vccd1 _6600_/B sky130_fd_sc_hd__a21oi_1
X_5619_ _5466_/X _5618_/X _5403_/A vssd1 vssd1 vccd1 vccd1 _5619_/X sky130_fd_sc_hd__a21o_1
X_5381__209 _5381__209/A vssd1 vssd1 vccd1 vccd1 _7181_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5804__266 _5805__267/A vssd1 vssd1 vccd1 vccd1 _7283_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5970_ _6723_/A vssd1 vssd1 vccd1 vccd1 _5970_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4921_ _4213_/X _7183_/Q _4929_/S vssd1 vssd1 vccd1 vccd1 _4922_/A sky130_fd_sc_hd__mux2_1
X_7640_ _7640_/CLK _7640_/D vssd1 vssd1 vccd1 vccd1 _7640_/Q sky130_fd_sc_hd__dfxtp_1
X_4852_ _4852_/A vssd1 vssd1 vccd1 vccd1 _7259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3803_ _7529_/Q _5461_/A vssd1 vssd1 vccd1 vccd1 _3865_/A sky130_fd_sc_hd__and2_1
XFILLER_21_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3303_ clkbuf_0__3303_/X vssd1 vssd1 vccd1 vccd1 _6788__169/A sky130_fd_sc_hd__clkbuf_4
X_7571_ _7571_/CLK _7571_/D vssd1 vssd1 vccd1 vccd1 _7571_/Q sky130_fd_sc_hd__dfxtp_1
X_4783_ _4728_/X _7285_/Q _4783_/S vssd1 vssd1 vccd1 vccd1 _4784_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3734_ _3734_/A vssd1 vssd1 vccd1 vccd1 _7741_/D sky130_fd_sc_hd__clkbuf_1
X_3665_ _3665_/A vssd1 vssd1 vccd1 vccd1 _7765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3234_ clkbuf_0__3234_/X vssd1 vssd1 vccd1 vccd1 _6730__124/A sky130_fd_sc_hd__clkbuf_4
X_5404_ _5404_/A vssd1 vssd1 vccd1 vccd1 _5404_/X sky130_fd_sc_hd__buf_2
X_3596_ _3554_/X _7791_/Q _3602_/S vssd1 vssd1 vccd1 vccd1 _3597_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5335_ _5335_/A vssd1 vssd1 vccd1 vccd1 _7156_/D sky130_fd_sc_hd__clkbuf_1
X_5266_ _5284_/A vssd1 vssd1 vccd1 vccd1 _5266_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_0__3133_ _6481_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3133_/X sky130_fd_sc_hd__clkbuf_16
X_6510__77 _6510__77/A vssd1 vssd1 vccd1 vccd1 _7622_/CLK sky130_fd_sc_hd__inv_2
X_7005_ _6996_/X _6997_/X _7817_/Q vssd1 vssd1 vccd1 vccd1 _7005_/X sky130_fd_sc_hd__a21o_1
X_4217_ _6310_/A _4217_/B _4284_/A vssd1 vssd1 vccd1 vccd1 _4240_/S sky130_fd_sc_hd__and3_4
X_5197_ _7134_/Q _5187_/X input11/X _5138_/D _5196_/X vssd1 vssd1 vccd1 vccd1 _5197_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4148_ _4148_/A vssd1 vssd1 vccd1 vccd1 _7571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4079_ _4079_/A vssd1 vssd1 vccd1 vccd1 _7600_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7838_ _7838_/CLK _7838_/D vssd1 vssd1 vccd1 vccd1 _7838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7769_ _7769_/CLK _7769_/D vssd1 vssd1 vccd1 vccd1 _7769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__2779_ _5834_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2779_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_50_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5120_ _7334_/Q _5120_/B vssd1 vssd1 vccd1 vccd1 _5121_/A sky130_fd_sc_hd__and2_1
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5051_ _5051_/A _5055_/B vssd1 vssd1 vccd1 vccd1 _5052_/A sky130_fd_sc_hd__or2_1
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6468__524 _6468__524/A vssd1 vssd1 vccd1 vccd1 _7589_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4002_ _4002_/A vssd1 vssd1 vccd1 vccd1 _7630_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5953_ _6016_/A vssd1 vssd1 vccd1 vccd1 _5953_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_52_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5884_ _5058_/A _7337_/Q _5884_/S vssd1 vssd1 vccd1 vccd1 _5885_/A sky130_fd_sc_hd__mux2_1
X_6757__144 _6757__144/A vssd1 vssd1 vccd1 vccd1 _7711_/CLK sky130_fd_sc_hd__inv_2
X_5258__186 _5259__187/A vssd1 vssd1 vccd1 vccd1 _7115_/CLK sky130_fd_sc_hd__inv_2
X_4904_ _4904_/A vssd1 vssd1 vccd1 vccd1 _7236_/D sky130_fd_sc_hd__clkbuf_1
X_4835_ _4811_/X _7266_/Q _4839_/S vssd1 vssd1 vccd1 vccd1 _4836_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7623_ _7623_/CLK _7623_/D vssd1 vssd1 vccd1 vccd1 _7623_/Q sky130_fd_sc_hd__dfxtp_1
X_6104__324 _6104__324/A vssd1 vssd1 vccd1 vccd1 _7373_/CLK sky130_fd_sc_hd__inv_2
X_7554_ _7554_/CLK _7554_/D vssd1 vssd1 vccd1 vccd1 _7554_/Q sky130_fd_sc_hd__dfxtp_1
X_4766_ _4766_/A vssd1 vssd1 vccd1 vccd1 _7293_/D sky130_fd_sc_hd__clkbuf_1
X_3717_ _3717_/A vssd1 vssd1 vccd1 vccd1 _7747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7892__219 vssd1 vssd1 vccd1 vccd1 _7892__219/HI partID[1] sky130_fd_sc_hd__conb_1
X_4697_ _4408_/X _7320_/Q _4697_/S vssd1 vssd1 vccd1 vccd1 _4698_/A sky130_fd_sc_hd__mux2_1
X_7485_ _7485_/CLK _7485_/D vssd1 vssd1 vccd1 vccd1 _7485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3648_ _3648_/A vssd1 vssd1 vccd1 vccd1 _7769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3579_ _3578_/X _7830_/Q _3579_/S vssd1 vssd1 vccd1 vccd1 _3580_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3148_ clkbuf_0__3148_/X vssd1 vssd1 vccd1 vccd1 _6642__114/A sky130_fd_sc_hd__clkbuf_4
X_6367_ _6373_/A vssd1 vssd1 vccd1 vccd1 _6367_/X sky130_fd_sc_hd__buf_1
X_5318_ _5318_/A _5892_/B vssd1 vssd1 vccd1 vccd1 _5334_/S sky130_fd_sc_hd__nand2_2
XFILLER_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3116_ _6392_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3116_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_48_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_2_wb_clk_i _7826_/CLK vssd1 vssd1 vccd1 vccd1 _7825_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5249_ _5249_/A vssd1 vssd1 vccd1 vccd1 _5249_/X sky130_fd_sc_hd__buf_1
XFILLER_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3295_ clkbuf_0__3295_/X vssd1 vssd1 vccd1 vccd1 _6745__134/A sky130_fd_sc_hd__clkbuf_4
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5916__312 _5916__312/A vssd1 vssd1 vccd1 vccd1 _7353_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1_0__2450_ clkbuf_0__2450_/X vssd1 vssd1 vccd1 vccd1 _5378__206/A sky130_fd_sc_hd__clkbuf_4
X_4620_ _3660_/X _7386_/Q _4624_/S vssd1 vssd1 vccd1 vccd1 _4621_/A sky130_fd_sc_hd__mux2_1
X_4551_ _4551_/A vssd1 vssd1 vccd1 vccd1 _7420_/D sky130_fd_sc_hd__clkbuf_1
X_4482_ _4482_/A vssd1 vssd1 vccd1 vccd1 _7451_/D sky130_fd_sc_hd__clkbuf_1
X_7270_ _7270_/CLK _7270_/D vssd1 vssd1 vccd1 vccd1 _7270_/Q sky130_fd_sc_hd__dfxtp_1
X_6221_ _7854_/Q _6911_/A vssd1 vssd1 vccd1 vccd1 _6222_/B sky130_fd_sc_hd__xor2_1
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5103_/A _5109_/B vssd1 vssd1 vccd1 vccd1 _5104_/A sky130_fd_sc_hd__and2_1
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6083_ _6099_/A _6083_/B vssd1 vssd1 vccd1 vccd1 _6083_/X sky130_fd_sc_hd__or2_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5034_/A vssd1 vssd1 vccd1 vccd1 _5034_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6985_ _7003_/A _6985_/B _6985_/C vssd1 vssd1 vccd1 vccd1 _6986_/A sky130_fd_sc_hd__and3_1
X_5936_ _5936_/A vssd1 vssd1 vccd1 vccd1 _6011_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5867_ _5867_/A vssd1 vssd1 vccd1 vccd1 _7329_/D sky130_fd_sc_hd__clkbuf_1
X_7606_ _7606_/CLK _7606_/D vssd1 vssd1 vccd1 vccd1 _7606_/Q sky130_fd_sc_hd__dfxtp_1
X_4818_ _4817_/X _7272_/Q _4818_/S vssd1 vssd1 vccd1 vccd1 _4819_/A sky130_fd_sc_hd__mux2_1
X_7537_ _7537_/CLK _7537_/D vssd1 vssd1 vccd1 vccd1 _7537_/Q sky130_fd_sc_hd__dfxtp_1
X_4749_ _4883_/A _4829_/B vssd1 vssd1 vccd1 vccd1 _4765_/S sky130_fd_sc_hd__nand2_4
XFILLER_119_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7468_ _7799_/CLK _7468_/D vssd1 vssd1 vccd1 vccd1 _7468_/Q sky130_fd_sc_hd__dfxtp_1
X_6419_ _6450_/A vssd1 vssd1 vccd1 vccd1 _6419_/X sky130_fd_sc_hd__buf_1
X_7399_ _7399_/CLK _7399_/D vssd1 vssd1 vccd1 vccd1 _7399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6343__425 _6343__425/A vssd1 vssd1 vccd1 vccd1 _7488_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3982_ _3982_/A vssd1 vssd1 vccd1 vccd1 _7639_/D sky130_fd_sc_hd__clkbuf_1
X_6770_ _6770_/A vssd1 vssd1 vccd1 vccd1 _6770_/X sky130_fd_sc_hd__buf_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5721_ _7221_/Q _7336_/Q _5725_/S vssd1 vssd1 vccd1 vccd1 _5722_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5652_ _5652_/A vssd1 vssd1 vccd1 vccd1 _7195_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4603_ _4603_/A vssd1 vssd1 vccd1 vccd1 _7394_/D sky130_fd_sc_hd__clkbuf_1
X_5583_ _7189_/Q _5453_/X _5582_/X vssd1 vssd1 vccd1 vccd1 _7189_/D sky130_fd_sc_hd__a21o_1
X_4534_ _4534_/A vssd1 vssd1 vccd1 vccd1 _7427_/D sky130_fd_sc_hd__clkbuf_1
X_7322_ _7322_/CLK _7322_/D vssd1 vssd1 vccd1 vccd1 _7322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4465_ _4465_/A vssd1 vssd1 vccd1 vccd1 _4465_/X sky130_fd_sc_hd__buf_2
X_7253_ _7253_/CLK _7253_/D vssd1 vssd1 vccd1 vccd1 _7253_/Q sky130_fd_sc_hd__dfxtp_1
X_7184_ _7855_/CLK _7184_/D vssd1 vssd1 vccd1 vccd1 _7184_/Q sky130_fd_sc_hd__dfxtp_1
X_6204_ _7801_/Q _7800_/Q _7799_/Q _6245_/A _7802_/Q vssd1 vssd1 vccd1 vccd1 _6231_/B
+ sky130_fd_sc_hd__a41o_1
X_4396_ _4418_/S vssd1 vssd1 vccd1 vccd1 _4409_/S sky130_fd_sc_hd__buf_2
XFILLER_100_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6066_ _7592_/Q _7560_/Q _7835_/Q _7536_/Q _6013_/X _6014_/X vssd1 vssd1 vccd1 vccd1
+ _6067_/B sky130_fd_sc_hd__mux4_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _5017_/A vssd1 vssd1 vccd1 vccd1 _5017_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3132_ clkbuf_0__3132_/X vssd1 vssd1 vccd1 vccd1 _6480__534/A sky130_fd_sc_hd__clkbuf_4
X_7032__51 _7035__54/A vssd1 vssd1 vccd1 vccd1 _7830_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6968_ _6966_/Y _6967_/X _6954_/X vssd1 vssd1 vccd1 vccd1 _7809_/D sky130_fd_sc_hd__a21oi_1
XFILLER_41_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5919_ _5925_/A vssd1 vssd1 vccd1 vccd1 _5919_/X sky130_fd_sc_hd__buf_1
X_6899_ _6916_/A _6900_/B vssd1 vssd1 vccd1 vccd1 _6899_/X sky130_fd_sc_hd__or2_1
XFILLER_22_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7898__225 vssd1 vssd1 vccd1 vccd1 _7898__225/HI partID[13] sky130_fd_sc_hd__conb_1
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6528__91 _6529__92/A vssd1 vssd1 vccd1 vccd1 _7636_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6846__40 _6848__42/A vssd1 vssd1 vccd1 vccd1 _7782_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5759__230 _5763__234/A vssd1 vssd1 vccd1 vccd1 _7247_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__2778_ clkbuf_0__2778_/X vssd1 vssd1 vccd1 vccd1 _5833__289/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4250_ _7827_/Q vssd1 vssd1 vccd1 vccd1 _4250_/X sky130_fd_sc_hd__clkbuf_4
X_4181_ _4181_/A vssd1 vssd1 vccd1 vccd1 _7561_/D sky130_fd_sc_hd__clkbuf_1
X_5365__195 _5369__199/A vssd1 vssd1 vccd1 vccd1 _7167_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3965_ _3965_/A vssd1 vssd1 vccd1 vccd1 _7646_/D sky130_fd_sc_hd__clkbuf_1
X_5704_ _5704_/A vssd1 vssd1 vccd1 vccd1 _7213_/D sky130_fd_sc_hd__clkbuf_1
X_6684_ _6684_/A vssd1 vssd1 vccd1 vccd1 _6684_/X sky130_fd_sc_hd__clkbuf_2
X_3896_ _3896_/A vssd1 vssd1 vccd1 vccd1 _7693_/D sky130_fd_sc_hd__clkbuf_1
X_5635_ _5633_/X _5634_/X _5245_/B vssd1 vssd1 vccd1 vccd1 _7192_/D sky130_fd_sc_hd__a21o_1
X_5566_ _5565_/X _7405_/Q _5457_/A _5459_/X vssd1 vssd1 vccd1 vccd1 _5566_/X sky130_fd_sc_hd__a31o_1
XFILLER_117_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5497_ _7060_/A vssd1 vssd1 vccd1 vccd1 _5497_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7305_ _7305_/CLK _7305_/D vssd1 vssd1 vccd1 vccd1 _7305_/Q sky130_fd_sc_hd__dfxtp_1
X_4517_ _7435_/Q _4233_/X _4521_/S vssd1 vssd1 vccd1 vccd1 _4518_/A sky130_fd_sc_hd__mux2_1
X_4448_ _3541_/X _4448_/B _4448_/C _4448_/D vssd1 vssd1 vccd1 vccd1 _4449_/A sky130_fd_sc_hd__nand4b_4
X_7236_ _7236_/CLK _7236_/D vssd1 vssd1 vccd1 vccd1 _7236_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3295_ _6740_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3295_/X sky130_fd_sc_hd__clkbuf_16
X_4379_ _7492_/Q _3932_/A _4385_/S vssd1 vssd1 vccd1 vccd1 _4380_/A sky130_fd_sc_hd__mux2_1
X_7167_ _7167_/CLK _7167_/D vssd1 vssd1 vccd1 vccd1 _7167_/Q sky130_fd_sc_hd__dfxtp_1
X_6118_ _6130_/A vssd1 vssd1 vccd1 vccd1 _6118_/X sky130_fd_sc_hd__buf_1
XFILLER_86_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7098_ _7098_/A vssd1 vssd1 vccd1 vccd1 _7853_/D sky130_fd_sc_hd__clkbuf_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _7789_/Q _7781_/Q _7773_/Q _7765_/Q _6031_/X _6011_/X vssd1 vssd1 vccd1 vccd1
+ _6049_/X sky130_fd_sc_hd__mux4_2
XFILLER_85_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3115_ clkbuf_0__3115_/X vssd1 vssd1 vccd1 vccd1 _6389__462/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f__3130_ clkbuf_0__3130_/X vssd1 vssd1 vccd1 vccd1 _6468__524/A sky130_fd_sc_hd__clkbuf_16
XFILLER_6_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2776_ clkbuf_0__2776_/X vssd1 vssd1 vccd1 vccd1 _6117_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6462__519 _6462__519/A vssd1 vssd1 vccd1 vccd1 _7584_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3750_ _3703_/X _7735_/Q _3756_/S vssd1 vssd1 vccd1 vccd1 _3751_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3681_ _3696_/S vssd1 vssd1 vccd1 vccd1 _3690_/S sky130_fd_sc_hd__buf_2
X_6751__139 _6751__139/A vssd1 vssd1 vccd1 vccd1 _7706_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6356__435 _6359__438/A vssd1 vssd1 vccd1 vccd1 _7498_/CLK sky130_fd_sc_hd__inv_2
X_5420_ _5417_/X _5418_/X _5590_/A vssd1 vssd1 vccd1 vccd1 _5420_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5351_ _7660_/Q _7659_/Q vssd1 vssd1 vccd1 vccd1 _5949_/B sky130_fd_sc_hd__nor2_1
X_5282_ _5282_/A vssd1 vssd1 vccd1 vccd1 _5307_/A sky130_fd_sc_hd__buf_2
X_4302_ _4285_/A _4302_/B vssd1 vssd1 vccd1 vccd1 _4302_/X sky130_fd_sc_hd__and2b_1
XFILLER_114_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6522__86 _6524__88/A vssd1 vssd1 vccd1 vccd1 _7631_/CLK sky130_fd_sc_hd__inv_2
X_7021_ _7021_/A vssd1 vssd1 vccd1 vccd1 _7824_/D sky130_fd_sc_hd__clkbuf_1
X_4233_ _7470_/Q vssd1 vssd1 vccd1 vccd1 _4233_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4164_ _4408_/A vssd1 vssd1 vccd1 vccd1 _4164_/X sky130_fd_sc_hd__clkbuf_4
X_4095_ _4095_/A vssd1 vssd1 vccd1 vccd1 _7593_/D sky130_fd_sc_hd__clkbuf_1
X_6840__35 _6842__37/A vssd1 vssd1 vccd1 vccd1 _7777_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7854_ _7854_/CLK _7854_/D vssd1 vssd1 vccd1 vccd1 _7854_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7785_ _7785_/CLK _7785_/D vssd1 vssd1 vccd1 vccd1 _7785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4997_ _4997_/A vssd1 vssd1 vccd1 vccd1 _4997_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3948_ _3947_/X _7652_/Q _3951_/S vssd1 vssd1 vccd1 vccd1 _3949_/A sky130_fd_sc_hd__mux2_1
X_6667_ _6656_/X _6658_/X _7671_/Q vssd1 vssd1 vccd1 vccd1 _6667_/Y sky130_fd_sc_hd__a21boi_1
X_3879_ _3879_/A vssd1 vssd1 vccd1 vccd1 _7700_/D sky130_fd_sc_hd__clkbuf_1
X_6598_ _7672_/Q vssd1 vssd1 vccd1 vccd1 _6598_/Y sky130_fd_sc_hd__inv_2
X_5618_ _7308_/Q _7236_/Q _7704_/Q _7324_/Q _5467_/X _4302_/B vssd1 vssd1 vccd1 vccd1
+ _5618_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5549_ _7692_/Q _7281_/Q _7164_/Q _7273_/Q _5426_/A _5518_/X vssd1 vssd1 vccd1 vccd1
+ _5549_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7219_ _7336_/CLK _7219_/D vssd1 vssd1 vccd1 vccd1 _7219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5251__181 _5252__182/A vssd1 vssd1 vccd1 vccd1 _7110_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_26_wb_clk_i _7474_/CLK vssd1 vssd1 vccd1 vccd1 _7854_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6169__371 _6169__371/A vssd1 vssd1 vccd1 vccd1 _7423_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4920_ _4935_/S vssd1 vssd1 vccd1 vccd1 _4929_/S sky130_fd_sc_hd__buf_2
X_4851_ _4808_/X _7259_/Q _4857_/S vssd1 vssd1 vccd1 vccd1 _4852_/A sky130_fd_sc_hd__mux2_1
X_3802_ _3802_/A _3802_/B _3802_/C vssd1 vssd1 vccd1 vccd1 _5461_/A sky130_fd_sc_hd__or3_2
Xclkbuf_1_1_0__3302_ clkbuf_0__3302_/X vssd1 vssd1 vccd1 vccd1 _6782__164/A sky130_fd_sc_hd__clkbuf_4
X_7570_ _7570_/CLK _7570_/D vssd1 vssd1 vccd1 vccd1 _7570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4782_ _4782_/A vssd1 vssd1 vccd1 vccd1 _7286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3733_ _3709_/X _7741_/Q _3735_/S vssd1 vssd1 vccd1 vccd1 _3734_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3664_ _7765_/Q _3663_/X _3667_/S vssd1 vssd1 vccd1 vccd1 _3665_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3233_ clkbuf_0__3233_/X vssd1 vssd1 vccd1 vccd1 _6645__116/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5403_ _5403_/A vssd1 vssd1 vccd1 vccd1 _5404_/A sky130_fd_sc_hd__clkinv_2
X_3595_ _3595_/A vssd1 vssd1 vccd1 vccd1 _7792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5334_ _7030_/A _7156_/Q _5334_/S vssd1 vssd1 vccd1 vccd1 _5335_/A sky130_fd_sc_hd__mux2_1
X_5265_ _5308_/A vssd1 vssd1 vccd1 vccd1 _5284_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3132_ _6475_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3132_/X sky130_fd_sc_hd__clkbuf_16
X_5196_ _7201_/Q _5217_/A _5198_/A vssd1 vssd1 vccd1 vccd1 _5196_/X sky130_fd_sc_hd__and3_1
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7004_ _7817_/Q _6995_/X _7002_/X _7003_/X vssd1 vssd1 vccd1 vccd1 _7816_/D sky130_fd_sc_hd__o211a_1
X_4216_ _4865_/B vssd1 vssd1 vccd1 vccd1 _4284_/A sky130_fd_sc_hd__clkbuf_2
X_4147_ _4069_/X _7571_/Q _4147_/S vssd1 vssd1 vccd1 vccd1 _4148_/A sky130_fd_sc_hd__mux2_1
X_6543__104 _6543__104/A vssd1 vssd1 vccd1 vccd1 _7649_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4078_ _4054_/X _7600_/Q _4082_/S vssd1 vssd1 vccd1 vccd1 _4079_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7837_ _7837_/CLK _7837_/D vssd1 vssd1 vccd1 vccd1 _7837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7768_ _7768_/CLK _7768_/D vssd1 vssd1 vccd1 vccd1 _7768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6719_ _6723_/A _6719_/B _6719_/C vssd1 vssd1 vccd1 vccd1 _6720_/A sky130_fd_sc_hd__and3_1
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2778_ _5828_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2778_/X sky130_fd_sc_hd__clkbuf_16
X_7699_ _7699_/CLK _7699_/D vssd1 vssd1 vccd1 vccd1 _7699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5810__271 _5812__273/A vssd1 vssd1 vccd1 vccd1 _7288_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5050_ _5050_/A vssd1 vssd1 vccd1 vccd1 _5050_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6433__495 _6435__497/A vssd1 vssd1 vccd1 vccd1 _7560_/CLK sky130_fd_sc_hd__inv_2
X_4001_ _3941_/X _7630_/Q _4001_/S vssd1 vssd1 vccd1 vccd1 _4002_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5952_ _6095_/A vssd1 vssd1 vccd1 vccd1 _6016_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4903_ _4803_/X _7236_/Q _4911_/S vssd1 vssd1 vccd1 vccd1 _4904_/A sky130_fd_sc_hd__mux2_1
X_5883_ _5883_/A vssd1 vssd1 vccd1 vccd1 _7336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4834_ _4834_/A vssd1 vssd1 vccd1 vccd1 _7267_/D sky130_fd_sc_hd__clkbuf_1
X_7622_ _7622_/CLK _7622_/D vssd1 vssd1 vccd1 vccd1 _7622_/Q sky130_fd_sc_hd__dfxtp_1
X_7553_ _7553_/CLK _7553_/D vssd1 vssd1 vccd1 vccd1 _7553_/Q sky130_fd_sc_hd__dfxtp_1
X_4765_ _4728_/X _7293_/Q _4765_/S vssd1 vssd1 vccd1 vccd1 _4766_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3716_ _3715_/X _7747_/Q _3722_/S vssd1 vssd1 vccd1 vccd1 _3717_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4696_ _4696_/A vssd1 vssd1 vccd1 vccd1 _7321_/D sky130_fd_sc_hd__clkbuf_1
X_7484_ _7484_/CLK _7484_/D vssd1 vssd1 vccd1 vccd1 _7484_/Q sky130_fd_sc_hd__dfxtp_1
X_3647_ _3578_/X _7769_/Q _3647_/S vssd1 vssd1 vccd1 vccd1 _3648_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3147_ clkbuf_0__3147_/X vssd1 vssd1 vccd1 vccd1 _6550__109/A sky130_fd_sc_hd__clkbuf_4
X_3578_ _3950_/A vssd1 vssd1 vccd1 vccd1 _3578_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5317_ _5338_/A _5317_/B vssd1 vssd1 vccd1 vccd1 _5892_/B sky130_fd_sc_hd__nor2_2
XFILLER_88_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__3115_ _6386_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3115_/X sky130_fd_sc_hd__clkbuf_16
X_5248_ _5795_/A vssd1 vssd1 vccd1 vccd1 _5248_/X sky130_fd_sc_hd__buf_1
X_6150__356 _6152__358/A vssd1 vssd1 vccd1 vccd1 _7408_/CLK sky130_fd_sc_hd__inv_2
X_5179_ _7194_/Q _5189_/B _5185_/C vssd1 vssd1 vccd1 vccd1 _5179_/X sky130_fd_sc_hd__and3_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5753__225 _5755__227/A vssd1 vssd1 vccd1 vccd1 _7242_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7866__193 vssd1 vssd1 vccd1 vccd1 _7866__193/HI core0Index[0] sky130_fd_sc_hd__conb_1
XFILLER_37_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3294_ clkbuf_0__3294_/X vssd1 vssd1 vccd1 vccd1 _6764_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4550_ _4253_/X _7420_/Q _4552_/S vssd1 vssd1 vccd1 vccd1 _4551_/A sky130_fd_sc_hd__mux2_1
X_4481_ _4411_/X _7451_/Q _4485_/S vssd1 vssd1 vccd1 vccd1 _4482_/A sky130_fd_sc_hd__mux2_1
X_6220_ _7795_/Q vssd1 vssd1 vccd1 vccd1 _6911_/A sky130_fd_sc_hd__clkbuf_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5102_/A vssd1 vssd1 vccd1 vccd1 _5102_/X sky130_fd_sc_hd__clkbuf_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6082_ _7593_/Q _7561_/Q _7836_/Q _7537_/Q _6013_/X _6014_/X vssd1 vssd1 vccd1 vccd1
+ _6083_/B sky130_fd_sc_hd__mux4_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5033_/A _5033_/B vssd1 vssd1 vccd1 vccd1 _5034_/A sky130_fd_sc_hd__or2_1
XFILLER_111_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5817__277 _5818__278/A vssd1 vssd1 vccd1 vccd1 _7294_/CLK sky130_fd_sc_hd__inv_2
X_6984_ _7813_/Q _6974_/B vssd1 vssd1 vccd1 vccd1 _6985_/C sky130_fd_sc_hd__or2b_1
X_5935_ _6024_/A vssd1 vssd1 vccd1 vccd1 _5935_/X sky130_fd_sc_hd__buf_4
X_5866_ _5040_/A _7329_/Q _5866_/S vssd1 vssd1 vccd1 vccd1 _5867_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4817_ _7471_/Q vssd1 vssd1 vccd1 vccd1 _4817_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7605_ _7605_/CLK _7605_/D vssd1 vssd1 vccd1 vccd1 _7605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7900__227 vssd1 vssd1 vccd1 vccd1 _7900__227/HI versionID[1] sky130_fd_sc_hd__conb_1
XFILLER_119_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7536_ _7536_/CLK _7536_/D vssd1 vssd1 vccd1 vccd1 _7536_/Q sky130_fd_sc_hd__dfxtp_1
X_4748_ _4748_/A vssd1 vssd1 vccd1 vccd1 _7301_/D sky130_fd_sc_hd__clkbuf_1
X_4679_ _4679_/A vssd1 vssd1 vccd1 vccd1 _7352_/D sky130_fd_sc_hd__clkbuf_1
X_7467_ _7467_/CLK _7467_/D vssd1 vssd1 vccd1 vccd1 _7467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7398_ _7398_/CLK _7398_/D vssd1 vssd1 vccd1 vccd1 _7398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3981_ _7639_/Q _3663_/X _3983_/S vssd1 vssd1 vccd1 vccd1 _3982_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5720_ _5720_/A vssd1 vssd1 vccd1 vccd1 _7220_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6283__395 _6286__398/A vssd1 vssd1 vccd1 vccd1 _7448_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5651_ _5667_/A _5651_/B vssd1 vssd1 vccd1 vccd1 _5652_/A sky130_fd_sc_hd__or2_1
X_4602_ _4250_/X _7394_/Q _4606_/S vssd1 vssd1 vccd1 vccd1 _4603_/A sky130_fd_sc_hd__mux2_1
X_5582_ _5634_/B _5566_/X _5581_/X _5497_/X vssd1 vssd1 vccd1 vccd1 _5582_/X sky130_fd_sc_hd__a31o_1
X_4533_ _4256_/X _7427_/Q _4533_/S vssd1 vssd1 vccd1 vccd1 _4534_/A sky130_fd_sc_hd__mux2_1
X_7321_ _7321_/CLK _7321_/D vssd1 vssd1 vccd1 vccd1 _7321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7252_ _7252_/CLK _7252_/D vssd1 vssd1 vccd1 vccd1 _7252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4464_ _5933_/A vssd1 vssd1 vccd1 vccd1 _4465_/A sky130_fd_sc_hd__clkbuf_4
X_6203_ _6233_/D _6245_/B vssd1 vssd1 vccd1 vccd1 _6231_/A sky130_fd_sc_hd__nand2_1
X_7183_ _7183_/CLK _7183_/D vssd1 vssd1 vccd1 vccd1 _7183_/Q sky130_fd_sc_hd__dfxtp_1
X_4395_ _4767_/A _4937_/B vssd1 vssd1 vccd1 vccd1 _4418_/S sky130_fd_sc_hd__nand2_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _7790_/Q _7782_/Q _7774_/Q _7766_/Q _6031_/X _6011_/X vssd1 vssd1 vccd1 vccd1
+ _6065_/X sky130_fd_sc_hd__mux4_2
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _7100_/A _5022_/B vssd1 vssd1 vccd1 vccd1 _5017_/A sky130_fd_sc_hd__or2_1
XFILLER_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3131_ clkbuf_0__3131_/X vssd1 vssd1 vccd1 vccd1 _6471__526/A sky130_fd_sc_hd__clkbuf_4
X_6967_ _6912_/X _6919_/X _6870_/B vssd1 vssd1 vccd1 vccd1 _6967_/X sky130_fd_sc_hd__a21o_1
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6303__410 _6306__413/A vssd1 vssd1 vccd1 vccd1 _7463_/CLK sky130_fd_sc_hd__inv_2
X_6898_ _7794_/Q vssd1 vssd1 vccd1 vccd1 _6916_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7519_ _7519_/CLK _7519_/D vssd1 vssd1 vccd1 vccd1 _7519_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_5_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6163__366 _6163__366/A vssd1 vssd1 vccd1 vccd1 _7418_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5766__235 _5770__239/A vssd1 vssd1 vccd1 vccd1 _7252_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4180_ _4051_/X _7561_/Q _4186_/S vssd1 vssd1 vccd1 vccd1 _4181_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3964_ _3941_/X _7646_/Q _3964_/S vssd1 vssd1 vccd1 vccd1 _3965_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5929__323 _5929__323/A vssd1 vssd1 vccd1 vccd1 _7364_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6752_ _6764_/A vssd1 vssd1 vccd1 vccd1 _6752_/X sky130_fd_sc_hd__buf_1
X_5703_ _7213_/Q _5107_/A _5703_/S vssd1 vssd1 vccd1 vccd1 _5704_/A sky130_fd_sc_hd__mux2_1
X_6683_ _6680_/X _6682_/X _6665_/X vssd1 vssd1 vccd1 vccd1 _7674_/D sky130_fd_sc_hd__a21oi_1
X_3895_ _3820_/X _7693_/Q _3899_/S vssd1 vssd1 vccd1 vccd1 _3896_/A sky130_fd_sc_hd__mux2_1
X_5634_ _7192_/Q _5634_/B vssd1 vssd1 vccd1 vccd1 _5634_/X sky130_fd_sc_hd__or2_1
XFILLER_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7858__232 vssd1 vssd1 vccd1 vccd1 partID[2] _7858__232/LO sky130_fd_sc_hd__conb_1
X_5565_ _7850_/Q vssd1 vssd1 vccd1 vccd1 _5565_/X sky130_fd_sc_hd__clkbuf_4
X_7304_ _7304_/CLK _7304_/D vssd1 vssd1 vccd1 vccd1 _7304_/Q sky130_fd_sc_hd__dfxtp_1
X_5496_ _5461_/Y _5463_/Y _5494_/X _5495_/X vssd1 vssd1 vccd1 vccd1 _5496_/X sky130_fd_sc_hd__a22o_1
X_4516_ _4516_/A vssd1 vssd1 vccd1 vccd1 _7436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4447_ _4447_/A _4447_/B _4447_/C vssd1 vssd1 vccd1 vccd1 _4448_/D sky130_fd_sc_hd__nor3_1
X_7235_ _7235_/CLK _7235_/D vssd1 vssd1 vccd1 vccd1 _7235_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3294_ _6739_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3294_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7166_ _7166_/CLK _7166_/D vssd1 vssd1 vccd1 vccd1 _7166_/Q sky130_fd_sc_hd__dfxtp_1
X_6117_ _6117_/A vssd1 vssd1 vccd1 vccd1 _6117_/X sky130_fd_sc_hd__buf_1
XFILLER_98_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4378_ _4378_/A vssd1 vssd1 vccd1 vccd1 _7493_/D sky130_fd_sc_hd__clkbuf_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _7106_/A _7097_/B _7097_/C vssd1 vssd1 vccd1 vccd1 _7098_/A sky130_fd_sc_hd__or3_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _5978_/X _6045_/X _6047_/X _5964_/X vssd1 vssd1 vccd1 vccd1 _6048_/X sky130_fd_sc_hd__o211a_1
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3114_ clkbuf_0__3114_/X vssd1 vssd1 vccd1 vccd1 _6413_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3680_ _4131_/D _3928_/B vssd1 vssd1 vccd1 vccd1 _3696_/S sky130_fd_sc_hd__or2_2
XFILLER_9_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5350_ _7687_/Q _5346_/X _5348_/X _6668_/B vssd1 vssd1 vccd1 vccd1 _5350_/X sky130_fd_sc_hd__a211o_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5281_ _5278_/X hold2/X _5274_/X _5275_/X _7126_/Q vssd1 vssd1 vccd1 vccd1 _7126_/D
+ sky130_fd_sc_hd__o32a_1
X_4301_ _4301_/A vssd1 vssd1 vccd1 vccd1 _4302_/B sky130_fd_sc_hd__buf_4
X_7020_ _7096_/A _7024_/B vssd1 vssd1 vccd1 vccd1 _7021_/A sky130_fd_sc_hd__and2_1
X_4232_ _4232_/A vssd1 vssd1 vccd1 vccd1 _7542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4163_ _4163_/A vssd1 vssd1 vccd1 vccd1 _7567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4094_ _4051_/X _7593_/Q _4100_/S vssd1 vssd1 vccd1 vccd1 _4095_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7853_ _7853_/CLK _7853_/D vssd1 vssd1 vccd1 vccd1 _7853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4996_ _5337_/B _5002_/B vssd1 vssd1 vccd1 vccd1 _4997_/A sky130_fd_sc_hd__and2_1
X_7784_ _7784_/CLK _7784_/D vssd1 vssd1 vccd1 vccd1 _7784_/Q sky130_fd_sc_hd__dfxtp_1
X_3947_ _3947_/A vssd1 vssd1 vccd1 vccd1 _3947_/X sky130_fd_sc_hd__clkbuf_4
X_6666_ _6662_/X _6664_/X _6665_/X vssd1 vssd1 vccd1 vccd1 _7670_/D sky130_fd_sc_hd__a21oi_1
X_3878_ _3828_/X _7700_/Q _3878_/S vssd1 vssd1 vccd1 vccd1 _3879_/A sky130_fd_sc_hd__mux2_1
X_6597_ _6606_/B _6606_/C vssd1 vssd1 vccd1 vccd1 _6682_/B sky130_fd_sc_hd__nand2_1
X_5617_ _7668_/Q _7501_/Q _7456_/Q _7316_/Q _5427_/X _5416_/X vssd1 vssd1 vccd1 vccd1
+ _5617_/X sky130_fd_sc_hd__mux4_1
X_5548_ _7297_/Q _7289_/Q _7265_/Q _7113_/Q _5502_/X _5416_/A vssd1 vssd1 vccd1 vccd1
+ _5548_/X sky130_fd_sc_hd__mux4_1
X_7218_ _7336_/CLK _7218_/D vssd1 vssd1 vccd1 vccd1 _7218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5479_ _5479_/A vssd1 vssd1 vccd1 vccd1 _5479_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_59_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7149_ _7687_/CLK _7149_/D vssd1 vssd1 vccd1 vccd1 _7149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5910__308 _5911__309/A vssd1 vssd1 vccd1 vccd1 _7349_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5836__291 _5839__294/A vssd1 vssd1 vccd1 vccd1 _7308_/CLK sky130_fd_sc_hd__inv_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4850_ _4850_/A vssd1 vssd1 vccd1 vccd1 _7260_/D sky130_fd_sc_hd__clkbuf_1
X_6362__440 _6363__441/A vssd1 vssd1 vccd1 vccd1 _7503_/CLK sky130_fd_sc_hd__inv_2
X_3801_ _4271_/A _4303_/C _4303_/D _3791_/B vssd1 vssd1 vccd1 vccd1 _3802_/C sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_1_1_0__3301_ clkbuf_0__3301_/X vssd1 vssd1 vccd1 vccd1 _6773__156/A sky130_fd_sc_hd__clkbuf_4
X_6520_ _6520_/A vssd1 vssd1 vccd1 vccd1 _6520_/X sky130_fd_sc_hd__buf_1
X_4781_ _4725_/X _7286_/Q _4783_/S vssd1 vssd1 vccd1 vccd1 _4782_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3732_ _3732_/A vssd1 vssd1 vccd1 vccd1 _7742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3663_ _7826_/Q vssd1 vssd1 vccd1 vccd1 _3663_/X sky130_fd_sc_hd__clkbuf_4
X_6451_ _6469_/A vssd1 vssd1 vccd1 vccd1 _6451_/X sky130_fd_sc_hd__buf_1
X_5402_ _5649_/A vssd1 vssd1 vccd1 vccd1 _5672_/D sky130_fd_sc_hd__clkbuf_2
X_5333_ _5333_/A vssd1 vssd1 vccd1 vccd1 _7155_/D sky130_fd_sc_hd__clkbuf_1
X_3594_ _3505_/X _7792_/Q _3602_/S vssd1 vssd1 vccd1 vccd1 _3595_/A sky130_fd_sc_hd__mux2_1
X_5264_ _5338_/A _5317_/B vssd1 vssd1 vccd1 vccd1 _5308_/A sky130_fd_sc_hd__or2_2
Xclkbuf_0__3131_ _6469_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3131_/X sky130_fd_sc_hd__clkbuf_16
X_6647__118 _6648__119/A vssd1 vssd1 vccd1 vccd1 _7665_/CLK sky130_fd_sc_hd__inv_2
X_5195_ _7133_/Q _5187_/X input10/X _5138_/D _5194_/X vssd1 vssd1 vccd1 vccd1 _5195_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4215_ _7524_/Q _4285_/A _4285_/B vssd1 vssd1 vccd1 vccd1 _4865_/B sky130_fd_sc_hd__and3_1
X_7003_ _7003_/A vssd1 vssd1 vccd1 vccd1 _7003_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4146_ _4146_/A vssd1 vssd1 vccd1 vccd1 _7572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6813__14 _6813__14/A vssd1 vssd1 vccd1 vccd1 _7756_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6805__7 _6807__9/A vssd1 vssd1 vccd1 vccd1 _7749_/CLK sky130_fd_sc_hd__inv_2
X_4077_ _4077_/A vssd1 vssd1 vccd1 vccd1 _7601_/D sky130_fd_sc_hd__clkbuf_1
X_7836_ _7836_/CLK _7836_/D vssd1 vssd1 vccd1 vccd1 _7836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7767_ _7767_/CLK _7767_/D vssd1 vssd1 vccd1 vccd1 _7767_/Q sky130_fd_sc_hd__dfxtp_1
X_4979_ _7113_/Q _4405_/A _4979_/S vssd1 vssd1 vccd1 vccd1 _4980_/A sky130_fd_sc_hd__mux2_1
X_6718_ _6718_/A _6726_/B vssd1 vssd1 vccd1 vccd1 _6719_/C sky130_fd_sc_hd__nand2_1
X_7698_ _7698_/CLK _7698_/D vssd1 vssd1 vccd1 vccd1 _7698_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2777_ _5827_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2777_/X sky130_fd_sc_hd__clkbuf_16
X_6649_ _6731_/A vssd1 vssd1 vccd1 vccd1 _6649_/X sky130_fd_sc_hd__buf_1
X_6550__109 _6550__109/A vssd1 vssd1 vccd1 vccd1 _7654_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4000_ _4000_/A vssd1 vssd1 vccd1 vccd1 _7631_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5951_ _5951_/A vssd1 vssd1 vccd1 vccd1 _5993_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4902_ _4917_/S vssd1 vssd1 vccd1 vccd1 _4911_/S sky130_fd_sc_hd__clkbuf_2
X_5882_ _5055_/A _7336_/Q _5884_/S vssd1 vssd1 vccd1 vccd1 _5883_/A sky130_fd_sc_hd__mux2_1
X_4833_ _4808_/X _7267_/Q _4839_/S vssd1 vssd1 vccd1 vccd1 _4834_/A sky130_fd_sc_hd__mux2_1
X_7621_ _7621_/CLK _7621_/D vssd1 vssd1 vccd1 vccd1 _7621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7552_ _7552_/CLK _7552_/D vssd1 vssd1 vccd1 vccd1 _7552_/Q sky130_fd_sc_hd__dfxtp_1
X_4764_ _4764_/A vssd1 vssd1 vccd1 vccd1 _7294_/D sky130_fd_sc_hd__clkbuf_1
X_3715_ _3944_/A vssd1 vssd1 vccd1 vccd1 _3715_/X sky130_fd_sc_hd__buf_2
X_7483_ _7483_/CLK _7483_/D vssd1 vssd1 vccd1 vccd1 _7483_/Q sky130_fd_sc_hd__dfxtp_1
X_4695_ _4405_/X _7321_/Q _4697_/S vssd1 vssd1 vccd1 vccd1 _4696_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3646_ _3646_/A vssd1 vssd1 vccd1 vccd1 _7770_/D sky130_fd_sc_hd__clkbuf_1
X_3577_ _7822_/Q vssd1 vssd1 vccd1 vccd1 _3950_/A sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__3146_ clkbuf_0__3146_/X vssd1 vssd1 vccd1 vccd1 _6731_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5316_ _5311_/X _7348_/Q _5274_/A _5284_/A _7148_/Q vssd1 vssd1 vccd1 vccd1 _7148_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5247_ _6300_/A vssd1 vssd1 vccd1 vccd1 _5247_/X sky130_fd_sc_hd__buf_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3114_ _6385_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3114_/X sky130_fd_sc_hd__clkbuf_16
X_5178_ _5200_/A vssd1 vssd1 vccd1 vccd1 _5189_/B sky130_fd_sc_hd__clkbuf_1
X_6369__446 _6372__449/A vssd1 vssd1 vccd1 vccd1 _7509_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4129_ _3840_/X _7579_/Q _4129_/S vssd1 vssd1 vccd1 vccd1 _4130_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7819_ _7819_/CLK _7819_/D vssd1 vssd1 vccd1 vccd1 _7819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5923__318 _5924__319/A vssd1 vssd1 vccd1 vccd1 _7359_/CLK sky130_fd_sc_hd__inv_2
X_4480_ _4480_/A vssd1 vssd1 vccd1 vccd1 _7452_/D sky130_fd_sc_hd__clkbuf_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5101_/A _5109_/B vssd1 vssd1 vccd1 vccd1 _5102_/A sky130_fd_sc_hd__and2_1
XFILLER_111_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6081_ _7791_/Q _7783_/Q _7775_/Q _7767_/Q _6031_/X _6011_/X vssd1 vssd1 vccd1 vccd1
+ _6081_/X sky130_fd_sc_hd__mux4_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5032_/A vssd1 vssd1 vccd1 vccd1 _5032_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7329_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6983_ _6983_/A _6983_/B _6982_/X vssd1 vssd1 vccd1 vccd1 _6985_/B sky130_fd_sc_hd__or3b_1
X_5934_ _7721_/Q _7705_/Q _7424_/Q _7486_/Q _5933_/X _4457_/A vssd1 vssd1 vccd1 vccd1
+ _5934_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5865_ _5865_/A vssd1 vssd1 vccd1 vccd1 _7328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4816_ _4816_/A vssd1 vssd1 vccd1 vccd1 _7273_/D sky130_fd_sc_hd__clkbuf_1
X_7604_ _7604_/CLK _7604_/D vssd1 vssd1 vccd1 vccd1 _7604_/Q sky130_fd_sc_hd__dfxtp_1
X_5796_ _5820_/A vssd1 vssd1 vccd1 vccd1 _5796_/X sky130_fd_sc_hd__buf_1
XFILLER_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7535_ _7535_/CLK _7535_/D vssd1 vssd1 vccd1 vccd1 _7535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4747_ _4728_/X _7301_/Q _4747_/S vssd1 vssd1 vccd1 vccd1 _4748_/A sky130_fd_sc_hd__mux2_1
X_4678_ _3666_/X _7352_/Q _4678_/S vssd1 vssd1 vccd1 vccd1 _4679_/A sky130_fd_sc_hd__mux2_1
X_7466_ _7466_/CLK _7466_/D vssd1 vssd1 vccd1 vccd1 _7466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7397_ _7397_/CLK _7397_/D vssd1 vssd1 vccd1 vccd1 _7397_/Q sky130_fd_sc_hd__dfxtp_1
X_3629_ _3629_/A vssd1 vssd1 vccd1 vccd1 _7777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6858__50 _6858__50/A vssd1 vssd1 vccd1 vccd1 _7792_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3129_ clkbuf_0__3129_/X vssd1 vssd1 vccd1 vccd1 _6459__516/A sky130_fd_sc_hd__clkbuf_4
X_6348_ _6348_/A vssd1 vssd1 vccd1 vccd1 _6348_/X sky130_fd_sc_hd__buf_1
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7882__209 vssd1 vssd1 vccd1 vccd1 _7882__209/HI manufacturerID[1] sky130_fd_sc_hd__conb_1
X_3980_ _3980_/A vssd1 vssd1 vccd1 vccd1 _7640_/D sky130_fd_sc_hd__clkbuf_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5650_ _6242_/A _5649_/X _5638_/X _7195_/Q _5639_/X vssd1 vssd1 vccd1 vccd1 _5651_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_43_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4601_ _4601_/A vssd1 vssd1 vccd1 vccd1 _7395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5581_ _7467_/Q _5463_/Y _5580_/X _5495_/X vssd1 vssd1 vccd1 vccd1 _5581_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4532_ _4532_/A vssd1 vssd1 vccd1 vccd1 _7428_/D sky130_fd_sc_hd__clkbuf_1
X_7320_ _7320_/CLK _7320_/D vssd1 vssd1 vccd1 vccd1 _7320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4463_ _6031_/A vssd1 vssd1 vccd1 vccd1 _5933_/A sky130_fd_sc_hd__clkbuf_4
X_7251_ _7251_/CLK _7251_/D vssd1 vssd1 vccd1 vccd1 _7251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6202_ _6883_/A _6883_/B _6605_/A vssd1 vssd1 vccd1 vccd1 _6991_/A sky130_fd_sc_hd__a21o_1
X_5823__282 _5824__283/A vssd1 vssd1 vccd1 vccd1 _7299_/CLK sky130_fd_sc_hd__inv_2
X_7182_ _7182_/CLK _7182_/D vssd1 vssd1 vccd1 vccd1 _7182_/Q sky130_fd_sc_hd__dfxtp_1
X_4394_ _4394_/A _4394_/B _4901_/C vssd1 vssd1 vccd1 vccd1 _4937_/B sky130_fd_sc_hd__and3_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _5978_/X _6061_/X _6063_/X _5964_/A vssd1 vssd1 vccd1 vccd1 _6064_/X sky130_fd_sc_hd__o211a_1
XFILLER_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5015_ _5015_/A vssd1 vssd1 vccd1 vccd1 _7100_/A sky130_fd_sc_hd__buf_6
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5377__205 _5378__206/A vssd1 vssd1 vccd1 vccd1 _7177_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6966_ _7809_/Q _6969_/B vssd1 vssd1 vccd1 vccd1 _6966_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5830__286 _5830__286/A vssd1 vssd1 vccd1 vccd1 _7303_/CLK sky130_fd_sc_hd__inv_2
X_6897_ _6897_/A _6897_/B vssd1 vssd1 vccd1 vccd1 _6897_/X sky130_fd_sc_hd__or2_1
XFILLER_108_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7518_ _7518_/CLK _7518_/D vssd1 vssd1 vccd1 vccd1 _7518_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_107_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7449_ _7449_/CLK _7449_/D vssd1 vssd1 vccd1 vccd1 _7449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6534__96 _6535__97/A vssd1 vssd1 vccd1 vccd1 _7641_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6852__45 _6856__49/A vssd1 vssd1 vccd1 vccd1 _7787_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6820_ _6826_/A vssd1 vssd1 vccd1 vccd1 _6820_/X sky130_fd_sc_hd__buf_1
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3963_ _3963_/A vssd1 vssd1 vccd1 vccd1 _7647_/D sky130_fd_sc_hd__clkbuf_1
X_5702_ _5702_/A vssd1 vssd1 vccd1 vccd1 _7212_/D sky130_fd_sc_hd__clkbuf_1
X_6682_ _6708_/A _6682_/B _6702_/C vssd1 vssd1 vccd1 vccd1 _6682_/X sky130_fd_sc_hd__or3_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_3894_ _3894_/A vssd1 vssd1 vccd1 vccd1 _7694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5633_ _5448_/X _5631_/X _5632_/X _7092_/B vssd1 vssd1 vccd1 vccd1 _5633_/X sky130_fd_sc_hd__a211o_1
XFILLER_117_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5564_ _7188_/Q _5453_/X _5563_/X vssd1 vssd1 vccd1 vccd1 _7188_/D sky130_fd_sc_hd__a21o_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4515_ _7436_/Q _4230_/X _4515_/S vssd1 vssd1 vccd1 vccd1 _4516_/A sky130_fd_sc_hd__mux2_1
X_7303_ _7303_/CLK _7303_/D vssd1 vssd1 vccd1 vccd1 _7303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5495_ _5495_/A vssd1 vssd1 vccd1 vccd1 _5495_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4446_ _4446_/A vssd1 vssd1 vccd1 vccd1 _4450_/A sky130_fd_sc_hd__clkbuf_4
X_7234_ _7234_/CLK _7234_/D vssd1 vssd1 vccd1 vccd1 _7234_/Q sky130_fd_sc_hd__dfxtp_1
X_4377_ _7493_/Q _3926_/A _4385_/S vssd1 vssd1 vccd1 vccd1 _4378_/A sky130_fd_sc_hd__mux2_1
X_7165_ _7165_/CLK _7165_/D vssd1 vssd1 vccd1 vccd1 _7165_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7096_ _7096_/A _7105_/B _7100_/C vssd1 vssd1 vccd1 vccd1 _7097_/C sky130_fd_sc_hd__and3_1
XFILLER_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _6079_/A _6047_/B vssd1 vssd1 vccd1 vccd1 _6047_/X sky130_fd_sc_hd__or2_1
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3113_ clkbuf_0__3113_/X vssd1 vssd1 vccd1 vccd1 _6384__459/A sky130_fd_sc_hd__clkbuf_4
X_6949_ _7804_/Q _6952_/B vssd1 vssd1 vccd1 vccd1 _6949_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5772__240 _5775__243/A vssd1 vssd1 vccd1 vccd1 _7257_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5280_ _5278_/X _7325_/Q _5274_/X _5275_/X _7125_/Q vssd1 vssd1 vccd1 vccd1 _7125_/D
+ sky130_fd_sc_hd__o32a_1
X_4300_ _4300_/A vssd1 vssd1 vccd1 vccd1 _4305_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4231_ _7542_/Q _4230_/X _4231_/S vssd1 vssd1 vccd1 vccd1 _4232_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7888__215 vssd1 vssd1 vccd1 vccd1 _7888__215/HI manufacturerID[7] sky130_fd_sc_hd__conb_1
X_4162_ _4161_/X _7567_/Q _4165_/S vssd1 vssd1 vccd1 vccd1 _4163_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4093_ _4093_/A vssd1 vssd1 vccd1 vccd1 _7594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7852_ _7854_/CLK _7852_/D vssd1 vssd1 vccd1 vccd1 _7852_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4995_ _5122_/A vssd1 vssd1 vccd1 vccd1 _5002_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7783_ _7783_/CLK _7783_/D vssd1 vssd1 vccd1 vccd1 _7783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3946_ _3946_/A vssd1 vssd1 vccd1 vccd1 _7653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6665_ _6690_/A vssd1 vssd1 vccd1 vccd1 _6665_/X sky130_fd_sc_hd__clkbuf_2
X_3877_ _3877_/A vssd1 vssd1 vccd1 vccd1 _7701_/D sky130_fd_sc_hd__clkbuf_1
X_6596_ _6595_/B _6602_/B _6595_/A vssd1 vssd1 vccd1 vccd1 _6606_/C sky130_fd_sc_hd__a21o_1
X_5616_ _5433_/S _5611_/X _5613_/Y _5615_/Y vssd1 vssd1 vccd1 vccd1 _5616_/X sky130_fd_sc_hd__a2bb2o_1
X_5547_ _7851_/Q _7405_/Q _5457_/A _5459_/X vssd1 vssd1 vccd1 vccd1 _5547_/X sky130_fd_sc_hd__a31o_1
XFILLER_2_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5478_ _7518_/Q vssd1 vssd1 vccd1 vccd1 _5518_/A sky130_fd_sc_hd__buf_2
X_7217_ _7333_/CLK _7217_/D vssd1 vssd1 vccd1 vccd1 _7217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4429_ _3991_/C _4431_/B _6328_/B vssd1 vssd1 vccd1 vccd1 _4429_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_113_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7148_ _7685_/CLK _7148_/D vssd1 vssd1 vccd1 vccd1 _7148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7079_ _6872_/A _7030_/A _7100_/C vssd1 vssd1 vccd1 vccd1 _7080_/B sky130_fd_sc_hd__mux2_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3800_ _3800_/A _3800_/B vssd1 vssd1 vccd1 vccd1 _3802_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4780_ _4780_/A vssd1 vssd1 vccd1 vccd1 _7287_/D sky130_fd_sc_hd__clkbuf_1
X_3731_ _3706_/X _7742_/Q _3735_/S vssd1 vssd1 vccd1 vccd1 _3732_/A sky130_fd_sc_hd__mux2_1
X_6403__471 _6404__472/A vssd1 vssd1 vccd1 vccd1 _7536_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3300_ clkbuf_0__3300_/X vssd1 vssd1 vccd1 vccd1 _6795_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_35_wb_clk_i _7474_/CLK vssd1 vssd1 vccd1 vccd1 _7821_/CLK sky130_fd_sc_hd__clkbuf_16
X_3662_ _3662_/A vssd1 vssd1 vccd1 vccd1 _7766_/D sky130_fd_sc_hd__clkbuf_1
X_6450_ _6450_/A vssd1 vssd1 vccd1 vccd1 _6450_/X sky130_fd_sc_hd__buf_1
X_3593_ _3608_/S vssd1 vssd1 vccd1 vccd1 _3602_/S sky130_fd_sc_hd__buf_2
X_5401_ _5462_/A _7040_/B _5401_/C _5493_/C vssd1 vssd1 vccd1 vccd1 _5649_/A sky130_fd_sc_hd__nor4_1
X_5332_ _7028_/A hold1/A _5334_/S vssd1 vssd1 vccd1 vccd1 _5333_/A sky130_fd_sc_hd__mux2_1
X_6176__377 _6177__378/A vssd1 vssd1 vccd1 vccd1 _7429_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3130_ _6463_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3130_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_114_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5263_ _7158_/Q _7157_/Q vssd1 vssd1 vccd1 vccd1 _5317_/B sky130_fd_sc_hd__nand2b_2
XFILLER_88_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5779__246 _5779__246/A vssd1 vssd1 vccd1 vccd1 _7263_/CLK sky130_fd_sc_hd__inv_2
X_5194_ _7200_/Q _5217_/A _5198_/A vssd1 vssd1 vccd1 vccd1 _5194_/X sky130_fd_sc_hd__and3_1
X_7002_ _6996_/X _6997_/X _7816_/Q vssd1 vssd1 vccd1 vccd1 _7002_/X sky130_fd_sc_hd__a21o_1
X_4214_ _4686_/A vssd1 vssd1 vccd1 vccd1 _6310_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4145_ _4066_/X _7572_/Q _4147_/S vssd1 vssd1 vccd1 vccd1 _4146_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6445__505 _6449__509/A vssd1 vssd1 vccd1 vccd1 _7570_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4076_ _4051_/X _7601_/Q _4082_/S vssd1 vssd1 vccd1 vccd1 _4077_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7835_ _7835_/CLK _7835_/D vssd1 vssd1 vccd1 vccd1 _7835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7766_ _7766_/CLK _7766_/D vssd1 vssd1 vccd1 vccd1 _7766_/Q sky130_fd_sc_hd__dfxtp_1
X_4978_ _4978_/A vssd1 vssd1 vccd1 vccd1 _7114_/D sky130_fd_sc_hd__clkbuf_1
X_6717_ _6637_/A _6676_/A _6684_/A _6630_/A vssd1 vssd1 vccd1 vccd1 _6726_/B sky130_fd_sc_hd__o211a_1
X_3929_ _3951_/S vssd1 vssd1 vccd1 vccd1 _3942_/S sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__2776_ _5826_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2776_/X sky130_fd_sc_hd__clkbuf_16
X_7697_ _7697_/CLK _7697_/D vssd1 vssd1 vccd1 vccd1 _7697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6579_ _7670_/Q _7669_/Q _7671_/Q vssd1 vssd1 vccd1 vccd1 _6670_/C sky130_fd_sc_hd__a21o_1
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__2389_ clkbuf_0__2389_/X vssd1 vssd1 vccd1 vccd1 _6300_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5950_ _5950_/A _4449_/A vssd1 vssd1 vccd1 vccd1 _5951_/A sky130_fd_sc_hd__or2b_1
XFILLER_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4901_ _4901_/A _4901_/B _4901_/C _4901_/D vssd1 vssd1 vccd1 vccd1 _4917_/S sky130_fd_sc_hd__or4_4
X_5881_ _5881_/A vssd1 vssd1 vccd1 vccd1 _7335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7620_ _7620_/CLK _7620_/D vssd1 vssd1 vccd1 vccd1 _7620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4832_ _4832_/A vssd1 vssd1 vccd1 vccd1 _7268_/D sky130_fd_sc_hd__clkbuf_1
X_7551_ _7551_/CLK _7551_/D vssd1 vssd1 vccd1 vccd1 _7551_/Q sky130_fd_sc_hd__dfxtp_1
X_4763_ _4725_/X _7294_/Q _4765_/S vssd1 vssd1 vccd1 vccd1 _4764_/A sky130_fd_sc_hd__mux2_1
X_3714_ _3714_/A vssd1 vssd1 vccd1 vccd1 _7748_/D sky130_fd_sc_hd__clkbuf_1
X_7482_ _7482_/CLK _7482_/D vssd1 vssd1 vccd1 vccd1 _7482_/Q sky130_fd_sc_hd__dfxtp_1
X_4694_ _4694_/A vssd1 vssd1 vccd1 vccd1 _7322_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3145_ clkbuf_0__3145_/X vssd1 vssd1 vccd1 vccd1 _6539__100/A sky130_fd_sc_hd__clkbuf_4
X_3645_ _3574_/X _7770_/Q _3647_/S vssd1 vssd1 vccd1 vccd1 _3646_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3576_ _3576_/A vssd1 vssd1 vccd1 vccd1 _7831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5315_ _5311_/X _7347_/Q _5274_/A _5284_/A _7147_/Q vssd1 vssd1 vccd1 vccd1 _7147_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_88_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3113_ _6379_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3113_/X sky130_fd_sc_hd__clkbuf_16
X_5246_ _5246_/A vssd1 vssd1 vccd1 vccd1 _5246_/X sky130_fd_sc_hd__buf_1
XFILLER_102_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5177_ _5177_/A vssd1 vssd1 vccd1 vccd1 _5177_/X sky130_fd_sc_hd__buf_2
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4128_ _4128_/A vssd1 vssd1 vccd1 vccd1 _7580_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3292_ clkbuf_0__3292_/X vssd1 vssd1 vccd1 vccd1 _6733__126/A sky130_fd_sc_hd__clkbuf_4
X_4059_ _4059_/A vssd1 vssd1 vccd1 vccd1 _7607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7818_ _7818_/CLK _7818_/D vssd1 vssd1 vccd1 vccd1 _7818_/Q sky130_fd_sc_hd__dfxtp_1
X_7749_ _7749_/CLK _7749_/D vssd1 vssd1 vccd1 vccd1 _7749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6486__57 _6486__57/A vssd1 vssd1 vccd1 vccd1 _7602_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5100_ _5122_/A vssd1 vssd1 vccd1 vccd1 _5109_/B sky130_fd_sc_hd__clkbuf_1
X_6080_ _5978_/X _6077_/X _6079_/X _5964_/A vssd1 vssd1 vccd1 vccd1 _6080_/X sky130_fd_sc_hd__o211a_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5031_/A _5033_/B vssd1 vssd1 vccd1 vccd1 _5032_/A sky130_fd_sc_hd__or2_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6982_ _6259_/A _6259_/B _6897_/X vssd1 vssd1 vccd1 vccd1 _6982_/X sky130_fd_sc_hd__a21o_1
X_5933_ _5933_/A vssd1 vssd1 vccd1 vccd1 _5933_/X sky130_fd_sc_hd__buf_4
XFILLER_34_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5864_ _5038_/A hold4/A _5866_/S vssd1 vssd1 vccd1 vccd1 _5865_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4815_ _4814_/X _7273_/Q _4818_/S vssd1 vssd1 vccd1 vccd1 _4816_/A sky130_fd_sc_hd__mux2_1
X_7603_ _7603_/CLK _7603_/D vssd1 vssd1 vccd1 vccd1 _7603_/Q sky130_fd_sc_hd__dfxtp_1
X_7534_ _7534_/CLK _7534_/D vssd1 vssd1 vccd1 vccd1 _7534_/Q sky130_fd_sc_hd__dfxtp_1
X_5795_ _5795_/A vssd1 vssd1 vccd1 vccd1 _5795_/X sky130_fd_sc_hd__buf_1
X_6295__405 _6298__408/A vssd1 vssd1 vccd1 vccd1 _7458_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4746_ _4746_/A vssd1 vssd1 vccd1 vccd1 _7302_/D sky130_fd_sc_hd__clkbuf_1
X_4677_ _4677_/A vssd1 vssd1 vccd1 vccd1 _7353_/D sky130_fd_sc_hd__clkbuf_1
X_7465_ _7465_/CLK _7465_/D vssd1 vssd1 vccd1 vccd1 _7465_/Q sky130_fd_sc_hd__dfxtp_2
X_6375__451 _6376__452/A vssd1 vssd1 vccd1 vccd1 _7514_/CLK sky130_fd_sc_hd__inv_2
X_7396_ _7396_/CLK _7396_/D vssd1 vssd1 vccd1 vccd1 _7396_/Q sky130_fd_sc_hd__dfxtp_1
X_3628_ _3578_/X _7777_/Q _3628_/S vssd1 vssd1 vccd1 vccd1 _3629_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3128_ clkbuf_0__3128_/X vssd1 vssd1 vccd1 vccd1 _6456__514/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3559_ _3558_/X _7835_/Q _3567_/S vssd1 vssd1 vccd1 vccd1 _3560_/A sky130_fd_sc_hd__mux2_1
X_5229_ _7145_/Q _5199_/A _5204_/A _5228_/X vssd1 vssd1 vccd1 vccd1 _5229_/X sky130_fd_sc_hd__o22a_4
XFILLER_102_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6458__515 _6459__516/A vssd1 vssd1 vccd1 vccd1 _7580_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_79_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6747__135 _6749__137/A vssd1 vssd1 vccd1 vccd1 _7702_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4600_ _4247_/X _7395_/Q _4606_/S vssd1 vssd1 vccd1 vccd1 _4601_/A sky130_fd_sc_hd__mux2_1
X_5580_ _5492_/Y _5579_/X _5493_/X vssd1 vssd1 vccd1 vccd1 _5580_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4531_ _4253_/X _7428_/Q _4533_/S vssd1 vssd1 vccd1 vccd1 _4532_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4462_ _7457_/Q vssd1 vssd1 vccd1 vccd1 _6031_/A sky130_fd_sc_hd__buf_2
X_7250_ _7250_/CLK _7250_/D vssd1 vssd1 vccd1 vccd1 _7250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6201_ _7847_/Q vssd1 vssd1 vccd1 vccd1 _6605_/A sky130_fd_sc_hd__inv_2
X_7181_ _7181_/CLK _7181_/D vssd1 vssd1 vccd1 vccd1 _7181_/Q sky130_fd_sc_hd__dfxtp_1
X_4393_ _4393_/A vssd1 vssd1 vccd1 vccd1 _4393_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6063_ _6079_/A _6063_/B vssd1 vssd1 vccd1 vccd1 _6063_/X sky130_fd_sc_hd__or2_1
XFILLER_97_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _5014_/A vssd1 vssd1 vccd1 vccd1 _5014_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _6963_/Y _6964_/X _6954_/X vssd1 vssd1 vccd1 vccd1 _7808_/D sky130_fd_sc_hd__a21oi_1
X_6896_ _6919_/A vssd1 vssd1 vccd1 vccd1 _6939_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7517_ _7517_/CLK _7517_/D vssd1 vssd1 vccd1 vccd1 _7517_/Q sky130_fd_sc_hd__dfxtp_1
X_4729_ _4728_/X _7309_/Q _4729_/S vssd1 vssd1 vccd1 vccd1 _4730_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7448_ _7448_/CLK _7448_/D vssd1 vssd1 vccd1 vccd1 _7448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7379_ _7379_/CLK _7379_/D vssd1 vssd1 vccd1 vccd1 _7379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__2389_ _5246_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2389_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_67_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2775_ clkbuf_0__2775_/X vssd1 vssd1 vccd1 vccd1 _5824__283/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5701_ _7212_/Q _5105_/A _5703_/S vssd1 vssd1 vccd1 vccd1 _5702_/A sky130_fd_sc_hd__mux2_1
X_3962_ _3938_/X _7647_/Q _3964_/S vssd1 vssd1 vccd1 vccd1 _3963_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6539__100 _6539__100/A vssd1 vssd1 vccd1 vccd1 _7645_/CLK sky130_fd_sc_hd__inv_2
X_6681_ _6714_/A vssd1 vssd1 vccd1 vccd1 _6708_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3893_ _3816_/X _7694_/Q _3899_/S vssd1 vssd1 vccd1 vccd1 _3894_/A sky130_fd_sc_hd__mux2_1
X_5632_ _5682_/A _5394_/C _7847_/Q _7406_/Q vssd1 vssd1 vccd1 vccd1 _5632_/X sky130_fd_sc_hd__and4bb_1
X_5563_ _5634_/B _5547_/X _5562_/X _5497_/X vssd1 vssd1 vccd1 vccd1 _5563_/X sky130_fd_sc_hd__a31o_1
XFILLER_117_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4514_ _4514_/A vssd1 vssd1 vccd1 vccd1 _7437_/D sky130_fd_sc_hd__clkbuf_1
X_7302_ _7302_/CLK _7302_/D vssd1 vssd1 vccd1 vccd1 _7302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5494_ _5490_/X _5492_/Y _5493_/X vssd1 vssd1 vccd1 vccd1 _5494_/X sky130_fd_sc_hd__a21o_1
XFILLER_117_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4445_ _6024_/A vssd1 vssd1 vccd1 vccd1 _4446_/A sky130_fd_sc_hd__buf_4
X_7233_ _7233_/CLK _7233_/D vssd1 vssd1 vccd1 vccd1 _7233_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3292_ _6731_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3292_/X sky130_fd_sc_hd__clkbuf_16
X_4376_ _4391_/S vssd1 vssd1 vccd1 vccd1 _4385_/S sky130_fd_sc_hd__buf_2
X_7164_ _7164_/CLK _7164_/D vssd1 vssd1 vccd1 vccd1 _7164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7104_/B _7095_/B vssd1 vssd1 vccd1 vccd1 _7097_/B sky130_fd_sc_hd__and2b_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _7393_/Q _7377_/Q _7647_/Q _7639_/Q _5983_/X _5984_/X vssd1 vssd1 vccd1 vccd1
+ _6047_/B sky130_fd_sc_hd__mux4_1
XFILLER_85_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3112_ clkbuf_0__3112_/X vssd1 vssd1 vccd1 vccd1 _6376__452/A sky130_fd_sc_hd__clkbuf_4
X_6948_ _6946_/Y _6947_/X _6935_/X vssd1 vssd1 vccd1 vccd1 _7803_/D sky130_fd_sc_hd__a21oi_1
XFILLER_53_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6879_ _6879_/A _6879_/B vssd1 vssd1 vccd1 vccd1 _6880_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6388__461 _6389__462/A vssd1 vssd1 vccd1 vccd1 _7524_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5848__301 _5849__302/A vssd1 vssd1 vccd1 vccd1 _7318_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4230_ _7471_/Q vssd1 vssd1 vccd1 vccd1 _4230_/X sky130_fd_sc_hd__buf_4
XFILLER_101_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4161_ _4405_/A vssd1 vssd1 vccd1 vccd1 _4161_/X sky130_fd_sc_hd__clkbuf_4
X_6825__24 _6825__24/A vssd1 vssd1 vccd1 vccd1 _7766_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4092_ _4046_/X _7594_/Q _4100_/S vssd1 vssd1 vccd1 vccd1 _4093_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7851_ _7853_/CLK _7851_/D vssd1 vssd1 vccd1 vccd1 _7851_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6802_ _6814_/A vssd1 vssd1 vccd1 vccd1 _6802_/X sky130_fd_sc_hd__buf_1
XFILLER_36_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4994_ _5004_/A vssd1 vssd1 vccd1 vccd1 _5122_/A sky130_fd_sc_hd__clkbuf_4
X_7782_ _7782_/CLK _7782_/D vssd1 vssd1 vccd1 vccd1 _7782_/Q sky130_fd_sc_hd__dfxtp_1
X_3945_ _3944_/X _7653_/Q _3951_/S vssd1 vssd1 vccd1 vccd1 _3946_/A sky130_fd_sc_hd__mux2_1
X_6664_ _6677_/A _6714_/C _6584_/B vssd1 vssd1 vccd1 vccd1 _6664_/X sky130_fd_sc_hd__or3b_1
XFILLER_23_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3876_ _3824_/X _7701_/Q _3878_/S vssd1 vssd1 vccd1 vccd1 _3877_/A sky130_fd_sc_hd__mux2_1
X_5615_ _5432_/S _5614_/X _5404_/X vssd1 vssd1 vccd1 vccd1 _5615_/Y sky130_fd_sc_hd__a21oi_1
X_6595_ _6595_/A _6595_/B _6602_/B vssd1 vssd1 vccd1 vccd1 _6606_/B sky130_fd_sc_hd__nand3_1
XFILLER_117_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5546_ _7187_/Q _5453_/X _5545_/X vssd1 vssd1 vccd1 vccd1 _7187_/D sky130_fd_sc_hd__a21o_1
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5477_ _5590_/A _5473_/X _5476_/X vssd1 vssd1 vccd1 vccd1 _5477_/X sky130_fd_sc_hd__a21o_1
X_7216_ _7333_/CLK _7216_/D vssd1 vssd1 vccd1 vccd1 _7216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4428_ _4428_/A vssd1 vssd1 vccd1 vccd1 _7465_/D sky130_fd_sc_hd__clkbuf_1
X_7147_ _7348_/CLK _7147_/D vssd1 vssd1 vccd1 vccd1 _7147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4359_ _4149_/X _7501_/Q _4367_/S vssd1 vssd1 vccd1 vccd1 _4360_/A sky130_fd_sc_hd__mux2_1
X_7078_ _7105_/C vssd1 vssd1 vccd1 vccd1 _7100_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_59_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_5_wb_clk_i _7826_/CLK vssd1 vssd1 vccd1 vccd1 _7829_/CLK sky130_fd_sc_hd__clkbuf_16
X_6029_ _6099_/A _6029_/B vssd1 vssd1 vccd1 vccd1 _6029_/X sky130_fd_sc_hd__or2_1
XFILLER_104_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7037__2 _7039__4/A vssd1 vssd1 vccd1 vccd1 _7835_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5843__297 _5843__297/A vssd1 vssd1 vccd1 vccd1 _7314_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3730_ _3730_/A vssd1 vssd1 vccd1 vccd1 _7743_/D sky130_fd_sc_hd__clkbuf_1
X_3661_ _7766_/Q _3660_/X _3667_/S vssd1 vssd1 vccd1 vccd1 _3662_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3592_ _3653_/B _4596_/A vssd1 vssd1 vccd1 vccd1 _3608_/S sky130_fd_sc_hd__nand2_2
X_5400_ _5491_/A vssd1 vssd1 vccd1 vccd1 _5493_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5331_ _5331_/A vssd1 vssd1 vccd1 vccd1 _7154_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5262_ _5274_/A vssd1 vssd1 vccd1 vccd1 _5262_/X sky130_fd_sc_hd__clkbuf_2
X_7001_ _7816_/Q _6995_/X _7000_/X _6909_/X vssd1 vssd1 vccd1 vccd1 _7815_/D sky130_fd_sc_hd__o211a_1
X_5193_ _7132_/Q _5187_/X input9/X _5138_/D _5192_/X vssd1 vssd1 vccd1 vccd1 _5193_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4213_ _7475_/Q vssd1 vssd1 vccd1 vccd1 _4213_/X sky130_fd_sc_hd__clkbuf_4
X_4144_ _4144_/A vssd1 vssd1 vccd1 vccd1 _7573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4075_ _4075_/A vssd1 vssd1 vccd1 vccd1 _7602_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7834_ _7834_/CLK _7834_/D vssd1 vssd1 vccd1 vccd1 _7834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7765_ _7765_/CLK _7765_/D vssd1 vssd1 vccd1 vccd1 _7765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6716_ _6725_/B _6630_/A _6714_/C _6718_/A vssd1 vssd1 vccd1 vccd1 _6719_/B sky130_fd_sc_hd__a31o_1
X_4977_ _7114_/Q _4402_/A _4979_/S vssd1 vssd1 vccd1 vccd1 _4978_/A sky130_fd_sc_hd__mux2_1
X_7696_ _7845_/CLK _7696_/D vssd1 vssd1 vccd1 vccd1 _7696_/Q sky130_fd_sc_hd__dfxtp_1
X_3928_ _4243_/B _3928_/B vssd1 vssd1 vccd1 vccd1 _3951_/S sky130_fd_sc_hd__or2_4
Xclkbuf_0__2775_ _5820_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2775_/X sky130_fd_sc_hd__clkbuf_16
X_3859_ _3721_/X _7705_/Q _3859_/S vssd1 vssd1 vccd1 vccd1 _3860_/A sky130_fd_sc_hd__mux2_1
X_6339__422 _6339__422/A vssd1 vssd1 vccd1 vccd1 _7485_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6578_ _7671_/Q _7670_/Q _6583_/B vssd1 vssd1 vccd1 vccd1 _6670_/B sky130_fd_sc_hd__nand3_1
X_5529_ _7852_/Q _6326_/A _5457_/X _5459_/X vssd1 vssd1 vccd1 vccd1 _5529_/X sky130_fd_sc_hd__a31o_1
XFILLER_105_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5880_ _5053_/A _7335_/Q _5884_/S vssd1 vssd1 vccd1 vccd1 _5881_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4900_ _4900_/A vssd1 vssd1 vccd1 vccd1 _7237_/D sky130_fd_sc_hd__clkbuf_1
X_6796__175 _6798__177/A vssd1 vssd1 vccd1 vccd1 _7742_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4831_ _4803_/X _7268_/Q _4839_/S vssd1 vssd1 vccd1 vccd1 _4832_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6143__355 _6153__359/A vssd1 vssd1 vccd1 vccd1 _7404_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7550_ _7550_/CLK _7550_/D vssd1 vssd1 vccd1 vccd1 _7550_/Q sky130_fd_sc_hd__dfxtp_1
X_5785__251 _5785__251/A vssd1 vssd1 vccd1 vccd1 _7268_/CLK sky130_fd_sc_hd__inv_2
X_4762_ _4762_/A vssd1 vssd1 vccd1 vccd1 _7295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3713_ _3712_/X _7748_/Q _3713_/S vssd1 vssd1 vccd1 vccd1 _3714_/A sky130_fd_sc_hd__mux2_1
X_4693_ _4402_/X _7322_/Q _4697_/S vssd1 vssd1 vccd1 vccd1 _4694_/A sky130_fd_sc_hd__mux2_1
X_7481_ _7481_/CLK _7481_/D vssd1 vssd1 vccd1 vccd1 _7481_/Q sky130_fd_sc_hd__dfxtp_1
X_6501_ _6501_/A vssd1 vssd1 vccd1 vccd1 _6501_/X sky130_fd_sc_hd__buf_1
X_3644_ _3644_/A vssd1 vssd1 vccd1 vccd1 _7771_/D sky130_fd_sc_hd__clkbuf_1
X_6432_ _6432_/A vssd1 vssd1 vccd1 vccd1 _6432_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3144_ clkbuf_0__3144_/X vssd1 vssd1 vccd1 vccd1 _6535__97/A sky130_fd_sc_hd__clkbuf_4
X_3575_ _3574_/X _7831_/Q _3579_/S vssd1 vssd1 vccd1 vccd1 _3576_/A sky130_fd_sc_hd__mux2_1
X_5314_ _5311_/X _7346_/Q _5307_/X _5308_/X _7146_/Q vssd1 vssd1 vccd1 vccd1 _7146_/D
+ sky130_fd_sc_hd__o32a_1
X_6294_ _6294_/A vssd1 vssd1 vccd1 vccd1 _6294_/X sky130_fd_sc_hd__buf_1
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5245_ _7203_/Q _5245_/B _5245_/C vssd1 vssd1 vccd1 vccd1 _7108_/D sky130_fd_sc_hd__nor3_1
Xclkbuf_0__3112_ _6373_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3112_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_102_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5176_ _7126_/Q _5173_/X input34/X _5163_/X _5175_/X vssd1 vssd1 vccd1 vccd1 _5176_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_28_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4127_ _3836_/X _7580_/Q _4129_/S vssd1 vssd1 vccd1 vccd1 _4128_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4058_ _4057_/X _7607_/Q _4061_/S vssd1 vssd1 vccd1 vccd1 _4059_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7817_ _7818_/CLK _7817_/D vssd1 vssd1 vccd1 vccd1 _7817_/Q sky130_fd_sc_hd__dfxtp_1
X_7748_ _7748_/CLK _7748_/D vssd1 vssd1 vccd1 vccd1 _7748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7679_ _7679_/CLK _7679_/D vssd1 vssd1 vccd1 vccd1 _7679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5030_/A vssd1 vssd1 vccd1 vccd1 _5030_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6981_ _7812_/Q _6974_/Y _6980_/X _6909_/X vssd1 vssd1 vccd1 vccd1 _7812_/D sky130_fd_sc_hd__o211a_1
X_5932_ _5932_/A vssd1 vssd1 vccd1 vccd1 _5932_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5863_ _5863_/A vssd1 vssd1 vccd1 vccd1 _7327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4814_ _7472_/Q vssd1 vssd1 vccd1 vccd1 _4814_/X sky130_fd_sc_hd__buf_2
X_7602_ _7602_/CLK _7602_/D vssd1 vssd1 vccd1 vccd1 _7602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7533_ _7533_/CLK _7533_/D vssd1 vssd1 vccd1 vccd1 _7533_/Q sky130_fd_sc_hd__dfxtp_1
X_4745_ _4725_/X _7302_/Q _4747_/S vssd1 vssd1 vccd1 vccd1 _4746_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4676_ _3663_/X _7353_/Q _4678_/S vssd1 vssd1 vccd1 vccd1 _4677_/A sky130_fd_sc_hd__mux2_1
X_7464_ _7464_/CLK _7464_/D vssd1 vssd1 vccd1 vccd1 _7464_/Q sky130_fd_sc_hd__dfxtp_1
X_7395_ _7395_/CLK _7395_/D vssd1 vssd1 vccd1 vccd1 _7395_/Q sky130_fd_sc_hd__dfxtp_1
X_3627_ _3627_/A vssd1 vssd1 vccd1 vccd1 _7778_/D sky130_fd_sc_hd__clkbuf_1
X_3558_ _3935_/A vssd1 vssd1 vccd1 vccd1 _3558_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3127_ clkbuf_0__3127_/X vssd1 vssd1 vccd1 vccd1 _6469_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6416__482 _6417__483/A vssd1 vssd1 vccd1 vccd1 _7547_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5228_ _5200_/X _5228_/B vssd1 vssd1 vccd1 vccd1 _5228_/X sky130_fd_sc_hd__and2b_1
XFILLER_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5159_ _5187_/A vssd1 vssd1 vccd1 vccd1 _5159_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6491__61 _6492__62/A vssd1 vssd1 vccd1 vccd1 _7606_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__2989_ clkbuf_0__2989_/X vssd1 vssd1 vccd1 vccd1 _6138__351/A sky130_fd_sc_hd__clkbuf_4
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4530_ _4530_/A vssd1 vssd1 vccd1 vccd1 _7429_/D sky130_fd_sc_hd__clkbuf_1
X_4461_ _4461_/A _4461_/B vssd1 vssd1 vccd1 vccd1 _7458_/D sky130_fd_sc_hd__nor2_1
XFILLER_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6200_ _6233_/D _6245_/B _7803_/Q vssd1 vssd1 vccd1 vccd1 _6883_/B sky130_fd_sc_hd__a21o_1
X_7180_ _7180_/CLK _7180_/D vssd1 vssd1 vccd1 vccd1 _7180_/Q sky130_fd_sc_hd__dfxtp_1
X_4392_ _4392_/A vssd1 vssd1 vccd1 vccd1 _7486_/D sky130_fd_sc_hd__clkbuf_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _7394_/Q _7378_/Q _7648_/Q _7640_/Q _5936_/A _5933_/A vssd1 vssd1 vccd1 vccd1
+ _6063_/B sky130_fd_sc_hd__mux4_2
XFILLER_100_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _7016_/A _5022_/B vssd1 vssd1 vccd1 vccd1 _5014_/A sky130_fd_sc_hd__or2_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6964_ _6912_/X _6919_/X _6888_/B vssd1 vssd1 vccd1 vccd1 _6964_/X sky130_fd_sc_hd__a21o_1
XFILLER_53_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6895_ _6870_/Y _6893_/X _6859_/A _6916_/B vssd1 vssd1 vccd1 vccd1 _6919_/A sky130_fd_sc_hd__o211ai_1
X_5846_ _5852_/A vssd1 vssd1 vccd1 vccd1 _5846_/X sky130_fd_sc_hd__buf_1
XFILLER_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5777_ _5789_/A vssd1 vssd1 vccd1 vccd1 _5777_/X sky130_fd_sc_hd__buf_1
XFILLER_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7516_ _7516_/CLK _7516_/D vssd1 vssd1 vccd1 vccd1 _7516_/Q sky130_fd_sc_hd__dfxtp_1
X_4728_ _7468_/Q vssd1 vssd1 vccd1 vccd1 _4728_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4659_ _4659_/A vssd1 vssd1 vccd1 vccd1 _7361_/D sky130_fd_sc_hd__clkbuf_1
X_7447_ _7447_/CLK _7447_/D vssd1 vssd1 vccd1 vccd1 _7447_/Q sky130_fd_sc_hd__dfxtp_1
X_7378_ _7378_/CLK _7378_/D vssd1 vssd1 vccd1 vccd1 _7378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6329_ _6329_/A vssd1 vssd1 vccd1 vccd1 _7477_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__2774_ clkbuf_0__2774_/X vssd1 vssd1 vccd1 vccd1 _5819__279/A sky130_fd_sc_hd__clkbuf_4
X_5798__261 _5799__262/A vssd1 vssd1 vccd1 vccd1 _7278_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6464__520 _6465__521/A vssd1 vssd1 vccd1 vccd1 _7585_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6753__140 _6753__140/A vssd1 vssd1 vccd1 vccd1 _7707_/CLK sky130_fd_sc_hd__inv_2
X_6519__84 _6519__84/A vssd1 vssd1 vccd1 vccd1 _7629_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6837__33 _6838__34/A vssd1 vssd1 vccd1 vccd1 _7775_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_wb_clk_i _7474_/CLK vssd1 vssd1 vccd1 vccd1 _7853_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3961_ _3961_/A vssd1 vssd1 vccd1 vccd1 _7648_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5700_ _5700_/A vssd1 vssd1 vccd1 vccd1 _7211_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6680_ _6679_/X _6661_/X _6595_/A vssd1 vssd1 vccd1 vccd1 _6680_/X sky130_fd_sc_hd__a21bo_1
X_3892_ _3892_/A vssd1 vssd1 vccd1 vccd1 _7695_/D sky130_fd_sc_hd__clkbuf_1
X_5631_ _7406_/Q _5457_/A _5396_/A _6396_/B vssd1 vssd1 vccd1 vccd1 _5631_/X sky130_fd_sc_hd__a31o_1
XFILLER_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5562_ _5676_/B _5463_/Y _5561_/X _5495_/X vssd1 vssd1 vccd1 vccd1 _5562_/X sky130_fd_sc_hd__a22o_1
XFILLER_8_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4513_ _7437_/Q _4227_/X _4515_/S vssd1 vssd1 vccd1 vccd1 _4514_/A sky130_fd_sc_hd__mux2_1
X_7301_ _7301_/CLK _7301_/D vssd1 vssd1 vccd1 vccd1 _7301_/Q sky130_fd_sc_hd__dfxtp_1
X_5493_ _5493_/A _5493_/B _5493_/C _5493_/D vssd1 vssd1 vccd1 vccd1 _5493_/X sky130_fd_sc_hd__or4_2
X_7232_ _7232_/CLK _7232_/D vssd1 vssd1 vccd1 vccd1 _7232_/Q sky130_fd_sc_hd__dfxtp_1
X_4444_ _7457_/Q vssd1 vssd1 vccd1 vccd1 _6024_/A sky130_fd_sc_hd__clkbuf_2
X_6333__417 _6333__417/A vssd1 vssd1 vccd1 vccd1 _7480_/CLK sky130_fd_sc_hd__inv_2
X_4375_ _4578_/A _4578_/B _4523_/B vssd1 vssd1 vccd1 vccd1 _4391_/S sky130_fd_sc_hd__and3_2
X_7163_ _7163_/CLK _7163_/D vssd1 vssd1 vccd1 vccd1 _7163_/Q sky130_fd_sc_hd__dfxtp_1
X_7094_ _7104_/B _7092_/Y _7093_/Y _5245_/B vssd1 vssd1 vccd1 vccd1 _7852_/D sky130_fd_sc_hd__a211oi_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _7412_/Q _7353_/Q _7420_/Q _7401_/Q _5979_/X _5980_/X vssd1 vssd1 vccd1 vccd1
+ _6045_/X sky130_fd_sc_hd__mux4_1
X_6546__105 _6550__109/A vssd1 vssd1 vccd1 vccd1 _7650_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7865__239 vssd1 vssd1 vccd1 vccd1 partID[15] _7865__239/LO sky130_fd_sc_hd__conb_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3111_ clkbuf_0__3111_/X vssd1 vssd1 vccd1 vccd1 _6372__449/A sky130_fd_sc_hd__clkbuf_4
X_6266__382 _6266__382/A vssd1 vssd1 vccd1 vccd1 _7435_/CLK sky130_fd_sc_hd__inv_2
X_6947_ _6943_/X _6939_/X _6883_/Y vssd1 vssd1 vccd1 vccd1 _6947_/X sky130_fd_sc_hd__a21o_1
XFILLER_53_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6878_ _7853_/Q _6878_/B vssd1 vssd1 vccd1 vccd1 _6882_/A sky130_fd_sc_hd__xor2_1
XFILLER_6_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6429__492 _6431__494/A vssd1 vssd1 vccd1 vccd1 _7557_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3309_ clkbuf_0__3309_/X vssd1 vssd1 vccd1 vccd1 _6818__18/A sky130_fd_sc_hd__clkbuf_4
XFILLER_45_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4160_ _4160_/A vssd1 vssd1 vccd1 vccd1 _7568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4091_ _4106_/S vssd1 vssd1 vccd1 vccd1 _4100_/S sky130_fd_sc_hd__buf_2
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7850_ _7853_/CLK _7850_/D vssd1 vssd1 vccd1 vccd1 _7850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6801_ _6832_/A vssd1 vssd1 vccd1 vccd1 _6801_/X sky130_fd_sc_hd__buf_1
XFILLER_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4993_ _5068_/A vssd1 vssd1 vccd1 vccd1 _5004_/A sky130_fd_sc_hd__inv_2
X_7781_ _7781_/CLK _7781_/D vssd1 vssd1 vccd1 vccd1 _7781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6107__326 _6108__327/A vssd1 vssd1 vccd1 vccd1 _7375_/CLK sky130_fd_sc_hd__inv_2
X_3944_ _3944_/A vssd1 vssd1 vccd1 vccd1 _3944_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6663_ _6676_/A vssd1 vssd1 vccd1 vccd1 _6714_/C sky130_fd_sc_hd__clkbuf_2
X_3875_ _3875_/A vssd1 vssd1 vccd1 vccd1 _7702_/D sky130_fd_sc_hd__clkbuf_1
X_5749__222 _5749__222/A vssd1 vssd1 vccd1 vccd1 _7239_/CLK sky130_fd_sc_hd__inv_2
X_5614_ _7517_/Q _7509_/Q _7448_/Q _7440_/Q _4302_/B _4297_/A vssd1 vssd1 vccd1 vccd1
+ _5614_/X sky130_fd_sc_hd__mux4_2
XFILLER_117_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6594_ _6594_/A vssd1 vssd1 vccd1 vccd1 _6602_/B sky130_fd_sc_hd__clkbuf_2
X_5545_ _5455_/X _5529_/X _5544_/X _5497_/X vssd1 vssd1 vccd1 vccd1 _5545_/X sky130_fd_sc_hd__a31o_1
XFILLER_105_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5476_ _5569_/S _5475_/X _5404_/A vssd1 vssd1 vccd1 vccd1 _5476_/X sky130_fd_sc_hd__a21o_1
XFILLER_117_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7215_ _7333_/CLK _7215_/D vssd1 vssd1 vccd1 vccd1 _7215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4427_ _4424_/X _4427_/B _6328_/B vssd1 vssd1 vccd1 vccd1 _4428_/A sky130_fd_sc_hd__and3b_1
X_7146_ _7348_/CLK _7146_/D vssd1 vssd1 vccd1 vccd1 _7146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ _4373_/S vssd1 vssd1 vccd1 vccd1 _4367_/S sky130_fd_sc_hd__buf_2
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7077_ _7077_/A _7077_/B vssd1 vssd1 vccd1 vccd1 _7105_/C sky130_fd_sc_hd__and2_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _7521_/Q vssd1 vssd1 vccd1 vccd1 _5403_/A sky130_fd_sc_hd__buf_2
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6028_ _7590_/Q _7558_/Q _7833_/Q _7534_/Q _5983_/X _5984_/X vssd1 vssd1 vccd1 vccd1
+ _6029_/B sky130_fd_sc_hd__mux4_1
XFILLER_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__2989_ _6136_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2989_/X sky130_fd_sc_hd__clkbuf_16
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3660_ _7827_/Q vssd1 vssd1 vccd1 vccd1 _3660_/X sky130_fd_sc_hd__clkbuf_4
X_7894__221 vssd1 vssd1 vccd1 vccd1 _7894__221/HI partID[5] sky130_fd_sc_hd__conb_1
XFILLER_70_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3591_ _3630_/D _3724_/A _4424_/C _3630_/C vssd1 vssd1 vccd1 vccd1 _4596_/A sky130_fd_sc_hd__and4bb_4
X_5330_ _7026_/A _7154_/Q _5334_/S vssd1 vssd1 vccd1 vccd1 _5331_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3091_ clkbuf_0__3091_/X vssd1 vssd1 vccd1 vccd1 _6307__414/A sky130_fd_sc_hd__clkbuf_4
X_5261_ _5282_/A vssd1 vssd1 vccd1 vccd1 _5274_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_114_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7000_ _6996_/X _6997_/X _7815_/Q vssd1 vssd1 vccd1 vccd1 _7000_/X sky130_fd_sc_hd__a21o_1
X_4212_ _4212_/A vssd1 vssd1 vccd1 vccd1 _7547_/D sky130_fd_sc_hd__clkbuf_1
X_5192_ _7199_/Q _5217_/A _5198_/A vssd1 vssd1 vccd1 vccd1 _5192_/X sky130_fd_sc_hd__and3_1
XFILLER_110_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4143_ _4063_/X _7573_/Q _4147_/S vssd1 vssd1 vccd1 vccd1 _4144_/A sky130_fd_sc_hd__mux2_1
X_6410__477 _6412__479/A vssd1 vssd1 vccd1 vccd1 _7542_/CLK sky130_fd_sc_hd__inv_2
X_4074_ _4046_/X _7602_/Q _4082_/S vssd1 vssd1 vccd1 vccd1 _4075_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7833_ _7833_/CLK _7833_/D vssd1 vssd1 vccd1 vccd1 _7833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7764_ _7764_/CLK _7764_/D vssd1 vssd1 vccd1 vccd1 _7764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6715_ _6713_/X _6714_/X _6690_/A vssd1 vssd1 vccd1 vccd1 _7684_/D sky130_fd_sc_hd__a21oi_1
XFILLER_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4976_ _4976_/A vssd1 vssd1 vccd1 vccd1 _7115_/D sky130_fd_sc_hd__clkbuf_1
X_3927_ _3927_/A _3927_/B _3927_/C vssd1 vssd1 vccd1 vccd1 _4243_/B sky130_fd_sc_hd__or3_4
X_7695_ _7695_/CLK _7695_/D vssd1 vssd1 vccd1 vccd1 _7695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__2774_ _5814_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2774_/X sky130_fd_sc_hd__clkbuf_16
X_3858_ _3858_/A vssd1 vssd1 vccd1 vccd1 _7706_/D sky130_fd_sc_hd__clkbuf_1
X_6734__127 _6736__129/A vssd1 vssd1 vccd1 vccd1 _7693_/CLK sky130_fd_sc_hd__inv_2
X_6577_ _7669_/Q vssd1 vssd1 vccd1 vccd1 _6583_/B sky130_fd_sc_hd__clkbuf_2
X_3789_ _7526_/Q vssd1 vssd1 vccd1 vccd1 _3907_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5528_ _7186_/Q _5453_/X _5527_/X vssd1 vssd1 vccd1 vccd1 _7186_/D sky130_fd_sc_hd__a21o_1
XFILLER_105_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5459_ _7040_/B _5493_/C _7040_/C vssd1 vssd1 vccd1 vccd1 _5459_/X sky130_fd_sc_hd__or3_2
X_6498__67 _6498__67/A vssd1 vssd1 vccd1 vccd1 _7612_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7129_ _7329_/CLK _7129_/D vssd1 vssd1 vccd1 vccd1 _7129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7878__205 vssd1 vssd1 vccd1 vccd1 _7878__205/HI core1Index[5] sky130_fd_sc_hd__conb_1
XFILLER_24_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6279__392 _6281__394/A vssd1 vssd1 vccd1 vccd1 _7445_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_2_0_wb_clk_i _7474_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_61_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4830_ _4845_/S vssd1 vssd1 vccd1 vccd1 _4839_/S sky130_fd_sc_hd__buf_2
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _4722_/X _7295_/Q _4765_/S vssd1 vssd1 vccd1 vccd1 _4762_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3712_ _3941_/A vssd1 vssd1 vccd1 vccd1 _3712_/X sky130_fd_sc_hd__clkbuf_2
X_4692_ _4692_/A vssd1 vssd1 vccd1 vccd1 _7323_/D sky130_fd_sc_hd__clkbuf_1
X_7480_ _7480_/CLK _7480_/D vssd1 vssd1 vccd1 vccd1 _7480_/Q sky130_fd_sc_hd__dfxtp_1
X_3643_ _3570_/X _7771_/Q _3647_/S vssd1 vssd1 vccd1 vccd1 _3644_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3143_ clkbuf_0__3143_/X vssd1 vssd1 vccd1 vccd1 _6531__94/A sky130_fd_sc_hd__clkbuf_4
X_5313_ _5311_/X _7345_/Q _5307_/X _5308_/X _7145_/Q vssd1 vssd1 vccd1 vccd1 _7145_/D
+ sky130_fd_sc_hd__o32a_1
X_3574_ _3947_/A vssd1 vssd1 vccd1 vccd1 _3574_/X sky130_fd_sc_hd__clkbuf_2
X_5244_ _5138_/C _5243_/X _5206_/X vssd1 vssd1 vccd1 vccd1 _5245_/C sky130_fd_sc_hd__a21oi_2
Xclkbuf_0__3111_ _6367_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3111_/X sky130_fd_sc_hd__clkbuf_16
X_5175_ _7193_/Q _5175_/B _5185_/C vssd1 vssd1 vccd1 vccd1 _5175_/X sky130_fd_sc_hd__and3_1
XFILLER_110_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4126_ _4126_/A vssd1 vssd1 vccd1 vccd1 _7581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4057_ _7826_/Q vssd1 vssd1 vccd1 vccd1 _4057_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_24_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7816_ _7818_/CLK _7816_/D vssd1 vssd1 vccd1 vccd1 _7816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7747_ _7747_/CLK _7747_/D vssd1 vssd1 vccd1 vccd1 _7747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4959_ _4221_/X _7166_/Q _4965_/S vssd1 vssd1 vccd1 vccd1 _4960_/A sky130_fd_sc_hd__mux2_1
X_7678_ _7680_/CLK _7678_/D vssd1 vssd1 vccd1 vccd1 _7678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6629_ _7840_/Q _6714_/B vssd1 vssd1 vccd1 vccd1 _6652_/C sky130_fd_sc_hd__xor2_1
X_6159__363 _6160__364/A vssd1 vssd1 vccd1 vccd1 _7415_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3309_ _6814_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3309_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6980_ _6996_/A _6259_/B _6979_/X _6974_/B _6983_/A vssd1 vssd1 vccd1 vccd1 _6980_/X
+ sky130_fd_sc_hd__a311o_1
X_5931_ _6631_/B vssd1 vssd1 vccd1 vccd1 _5931_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5862_ _5036_/A _7327_/Q _5866_/S vssd1 vssd1 vccd1 vccd1 _5863_/A sky130_fd_sc_hd__mux2_1
X_4813_ _4813_/A vssd1 vssd1 vccd1 vccd1 _7274_/D sky130_fd_sc_hd__clkbuf_1
X_7601_ _7601_/CLK _7601_/D vssd1 vssd1 vccd1 vccd1 _7601_/Q sky130_fd_sc_hd__dfxtp_1
X_7532_ _7532_/CLK _7532_/D vssd1 vssd1 vccd1 vccd1 _7532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4744_ _4744_/A vssd1 vssd1 vccd1 vccd1 _7303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4675_ _4675_/A vssd1 vssd1 vccd1 vccd1 _7354_/D sky130_fd_sc_hd__clkbuf_1
X_7463_ _7463_/CLK _7463_/D vssd1 vssd1 vccd1 vccd1 _7463_/Q sky130_fd_sc_hd__dfxtp_1
X_7394_ _7394_/CLK _7394_/D vssd1 vssd1 vccd1 vccd1 _7394_/Q sky130_fd_sc_hd__dfxtp_1
X_3626_ _3574_/X _7778_/Q _3628_/S vssd1 vssd1 vccd1 vccd1 _3627_/A sky130_fd_sc_hd__mux2_1
X_3557_ _7827_/Q vssd1 vssd1 vccd1 vccd1 _3935_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3126_ clkbuf_0__3126_/X vssd1 vssd1 vccd1 vccd1 _6448__508/A sky130_fd_sc_hd__clkbuf_4
X_6276_ _6282_/A vssd1 vssd1 vccd1 vccd1 _6276_/X sky130_fd_sc_hd__buf_1
X_5227_ _7144_/Q _5215_/X _5216_/X _5226_/X vssd1 vssd1 vccd1 vccd1 _5227_/X sky130_fd_sc_hd__o22a_4
X_5800__263 _5801__264/A vssd1 vssd1 vccd1 vccd1 _7280_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5158_ _7120_/Q _5145_/X input28/X _5146_/X _5157_/X vssd1 vssd1 vccd1 vccd1 _5158_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_56_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5089_ _5122_/A vssd1 vssd1 vccd1 vccd1 _5098_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4109_ _4686_/A vssd1 vssd1 vccd1 vccd1 _4865_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6382__457 _6384__459/A vssd1 vssd1 vccd1 vccd1 _7520_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6423__487 _6425__489/A vssd1 vssd1 vccd1 vccd1 _7552_/CLK sky130_fd_sc_hd__inv_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__2988_ clkbuf_0__2988_/X vssd1 vssd1 vccd1 vccd1 _6133__347/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5743__217 _5743__217/A vssd1 vssd1 vccd1 vccd1 _7234_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4460_ _4457_/A _4457_/B _4421_/X vssd1 vssd1 vccd1 vccd1 _4461_/B sky130_fd_sc_hd__o21ai_1
X_4391_ _7486_/Q _3950_/A _4391_/S vssd1 vssd1 vccd1 vccd1 _4392_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6130_ _6130_/A vssd1 vssd1 vccd1 vccd1 _6130_/X sky130_fd_sc_hd__buf_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _7413_/Q _7354_/Q _7421_/Q _7402_/Q _5979_/X _5942_/X vssd1 vssd1 vccd1 vccd1
+ _6061_/X sky130_fd_sc_hd__mux4_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5081_/B vssd1 vssd1 vccd1 vccd1 _5022_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_97_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6963_ _7808_/Q _6969_/B vssd1 vssd1 vccd1 vccd1 _6963_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6894_ _6900_/B vssd1 vssd1 vccd1 vccd1 _6916_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7515_ _7515_/CLK _7515_/D vssd1 vssd1 vccd1 vccd1 _7515_/Q sky130_fd_sc_hd__dfxtp_1
X_4727_ _4727_/A vssd1 vssd1 vccd1 vccd1 _7310_/D sky130_fd_sc_hd__clkbuf_1
X_7446_ _7446_/CLK _7446_/D vssd1 vssd1 vccd1 vccd1 _7446_/Q sky130_fd_sc_hd__dfxtp_1
X_4658_ _4405_/X _7361_/Q _4660_/S vssd1 vssd1 vccd1 vccd1 _4659_/A sky130_fd_sc_hd__mux2_1
X_3609_ _3609_/A vssd1 vssd1 vccd1 vccd1 _7785_/D sky130_fd_sc_hd__clkbuf_1
Xinput90 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _5337_/B sky130_fd_sc_hd__buf_8
X_7377_ _7377_/CLK _7377_/D vssd1 vssd1 vccd1 vccd1 _7377_/Q sky130_fd_sc_hd__dfxtp_1
X_4589_ _4589_/A vssd1 vssd1 vccd1 vccd1 _7400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3109_ clkbuf_0__3109_/X vssd1 vssd1 vccd1 vccd1 _6360__439/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6328_ _7696_/Q _6328_/B _6328_/C _6394_/A vssd1 vssd1 vccd1 vccd1 _6329_/A sky130_fd_sc_hd__and4b_1
XFILLER_1_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__2773_ clkbuf_0__2773_/X vssd1 vssd1 vccd1 vccd1 _5812__273/A sky130_fd_sc_hd__clkbuf_4
XFILLER_107_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6259_ _6259_/A _6259_/B vssd1 vssd1 vccd1 vccd1 _6897_/B sky130_fd_sc_hd__nor2_1
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5807__269 _5807__269/A vssd1 vssd1 vccd1 vccd1 _7286_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3960_ _3935_/X _7648_/Q _3964_/S vssd1 vssd1 vccd1 vccd1 _3961_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3891_ _3784_/X _7695_/Q _3899_/S vssd1 vssd1 vccd1 vccd1 _3892_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5630_ _5455_/X _5628_/X _5629_/X vssd1 vssd1 vccd1 vccd1 _7191_/D sky130_fd_sc_hd__a21o_1
X_5561_ _5492_/Y _5560_/X _5493_/X vssd1 vssd1 vccd1 vccd1 _5561_/X sky130_fd_sc_hd__a21o_1
X_5492_ _5492_/A _5492_/B vssd1 vssd1 vccd1 vccd1 _5492_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4512_ _4512_/A vssd1 vssd1 vccd1 vccd1 _7438_/D sky130_fd_sc_hd__clkbuf_1
X_7300_ _7300_/CLK _7300_/D vssd1 vssd1 vccd1 vccd1 _7300_/Q sky130_fd_sc_hd__dfxtp_1
X_7231_ _7231_/CLK _7231_/D vssd1 vssd1 vccd1 vccd1 _7231_/Q sky130_fd_sc_hd__dfxtp_1
X_4443_ _5998_/A vssd1 vssd1 vccd1 vccd1 _4457_/A sky130_fd_sc_hd__clkbuf_2
X_7162_ _7162_/CLK _7162_/D vssd1 vssd1 vccd1 vccd1 _7162_/Q sky130_fd_sc_hd__dfxtp_1
X_4374_ _4374_/A vssd1 vssd1 vccd1 vccd1 _7494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7093_ _7852_/Q _7104_/B vssd1 vssd1 vccd1 vccd1 _7093_/Y sky130_fd_sc_hd__nor2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6040_/X _6041_/X _6042_/X _6043_/X _5945_/X _4436_/X vssd1 vssd1 vccd1 vccd1
+ _6044_/X sky130_fd_sc_hd__mux4_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6946_ _7803_/Q _6952_/B vssd1 vssd1 vccd1 vccd1 _6946_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_1_0_0__3110_ clkbuf_0__3110_/X vssd1 vssd1 vccd1 vccd1 _6366__444/A sky130_fd_sc_hd__clkbuf_4
X_6877_ _6918_/A _7795_/Q vssd1 vssd1 vccd1 vccd1 _6878_/B sky130_fd_sc_hd__xor2_1
XFILLER_22_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5828_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5828_/X sky130_fd_sc_hd__buf_1
XFILLER_10_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7429_ _7429_/CLK _7429_/D vssd1 vssd1 vccd1 vccd1 _7429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6273__387 _6273__387/A vssd1 vssd1 vccd1 vccd1 _7440_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3308_ clkbuf_0__3308_/X vssd1 vssd1 vccd1 vccd1 _6812__13/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5855__307 _5855__307/A vssd1 vssd1 vccd1 vccd1 _7324_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4090_ _4243_/A _4131_/D vssd1 vssd1 vccd1 vccd1 _4106_/S sky130_fd_sc_hd__or2_2
XFILLER_75_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4992_ _5337_/C _5138_/C _5177_/A vssd1 vssd1 vccd1 vccd1 _5068_/A sky130_fd_sc_hd__nand3_4
X_7780_ _7780_/CLK _7780_/D vssd1 vssd1 vccd1 vccd1 _7780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3943_ _3943_/A vssd1 vssd1 vccd1 vccd1 _7654_/D sky130_fd_sc_hd__clkbuf_1
X_6731_ _6731_/A vssd1 vssd1 vccd1 vccd1 _6731_/X sky130_fd_sc_hd__buf_1
XFILLER_23_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6662_ _6640_/C _6661_/X _7670_/Q vssd1 vssd1 vccd1 vccd1 _6662_/X sky130_fd_sc_hd__a21bo_1
X_3874_ _3820_/X _7702_/Q _3878_/S vssd1 vssd1 vccd1 vccd1 _3875_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5613_ _5613_/A _5613_/B vssd1 vssd1 vccd1 vccd1 _5613_/Y sky130_fd_sc_hd__nand2_1
X_6593_ _6593_/A _6593_/B vssd1 vssd1 vccd1 vccd1 _6686_/B sky130_fd_sc_hd__nand2_2
X_6552__110 _6555__113/A vssd1 vssd1 vccd1 vccd1 _7655_/CLK sky130_fd_sc_hd__inv_2
X_5544_ _6328_/C _5463_/Y _5543_/X _5495_/X vssd1 vssd1 vccd1 vccd1 _5544_/X sky130_fd_sc_hd__a22o_1
XFILLER_8_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5475_ _7511_/Q _7503_/Q _7442_/Q _7434_/Q _4301_/A _5467_/X vssd1 vssd1 vccd1 vccd1
+ _5475_/X sky130_fd_sc_hd__mux4_2
XFILLER_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7214_ _7333_/CLK _7214_/D vssd1 vssd1 vccd1 vccd1 _7214_/Q sky130_fd_sc_hd__dfxtp_1
X_4426_ _4424_/B _4424_/C _4424_/A vssd1 vssd1 vccd1 vccd1 _4427_/B sky130_fd_sc_hd__a21o_1
X_7145_ _7348_/CLK _7145_/D vssd1 vssd1 vccd1 vccd1 _7145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ _4955_/A _4706_/A vssd1 vssd1 vccd1 vccd1 _4373_/S sky130_fd_sc_hd__or2_2
X_7076_ _7076_/A vssd1 vssd1 vccd1 vccd1 _7847_/D sky130_fd_sc_hd__clkbuf_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _7522_/Q vssd1 vssd1 vccd1 vccd1 _5434_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6027_ _7788_/Q _7780_/Q _7772_/Q _7764_/Q _5979_/X _5980_/X vssd1 vssd1 vccd1 vccd1
+ _6027_/X sky130_fd_sc_hd__mux4_2
XFILLER_74_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6831__29 _6831__29/A vssd1 vssd1 vccd1 vccd1 _7771_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2988_ _6130_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2988_/X sky130_fd_sc_hd__clkbuf_16
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _6927_/Y _6928_/X _7014_/A vssd1 vssd1 vccd1 vccd1 _7798_/D sky130_fd_sc_hd__a21oi_1
XFILLER_80_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6477__531 _6478__532/A vssd1 vssd1 vccd1 vccd1 _7596_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3590_ _7092_/A _3588_/X _5239_/A vssd1 vssd1 vccd1 vccd1 _3630_/C sky130_fd_sc_hd__a21oi_1
Xclkbuf_1_1_0__3090_ clkbuf_0__3090_/X vssd1 vssd1 vccd1 vccd1 _6342_/A sky130_fd_sc_hd__clkbuf_4
X_5260_ _7157_/Q _7158_/Q vssd1 vssd1 vccd1 vccd1 _5282_/A sky130_fd_sc_hd__or2b_1
X_4211_ _4173_/X _7547_/Q _4211_/S vssd1 vssd1 vccd1 vccd1 _4212_/A sky130_fd_sc_hd__mux2_1
X_5191_ _7108_/Q vssd1 vssd1 vccd1 vccd1 _5217_/A sky130_fd_sc_hd__clkbuf_2
X_6766__151 _6768__153/A vssd1 vssd1 vccd1 vccd1 _7718_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4142_ _4142_/A vssd1 vssd1 vccd1 vccd1 _7574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6113__331 _6113__331/A vssd1 vssd1 vccd1 vccd1 _7380_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4073_ _4088_/S vssd1 vssd1 vccd1 vccd1 _4082_/S sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_13_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7336_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7832_ _7832_/CLK _7832_/D vssd1 vssd1 vccd1 vccd1 _7832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7763_ _7763_/CLK _7763_/D vssd1 vssd1 vccd1 vccd1 _7763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4975_ _7115_/Q _4399_/A _4979_/S vssd1 vssd1 vccd1 vccd1 _4976_/A sky130_fd_sc_hd__mux2_1
X_3926_ _3926_/A vssd1 vssd1 vccd1 vccd1 _3926_/X sky130_fd_sc_hd__clkbuf_4
X_6714_ _6714_/A _6714_/B _6714_/C vssd1 vssd1 vccd1 vccd1 _6714_/X sky130_fd_sc_hd__or3_1
X_7694_ _7694_/CLK _7694_/D vssd1 vssd1 vccd1 vccd1 _7694_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2773_ _5808_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2773_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_109_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3857_ _3718_/X _7706_/Q _3859_/S vssd1 vssd1 vccd1 vccd1 _3858_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6576_ _6576_/A _6696_/B _6696_/C vssd1 vssd1 vccd1 vccd1 _6588_/B sky130_fd_sc_hd__nand3_1
X_3788_ _7524_/Q _7519_/Q vssd1 vssd1 vccd1 vccd1 _4304_/B sky130_fd_sc_hd__xnor2_2
XFILLER_118_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5527_ _5455_/X _5501_/X _5526_/X _5497_/X vssd1 vssd1 vccd1 vccd1 _5527_/X sky130_fd_sc_hd__a31o_1
XFILLER_117_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5458_ _7204_/Q _7205_/Q _5458_/C _5458_/D vssd1 vssd1 vccd1 vccd1 _7040_/C sky130_fd_sc_hd__or4_2
XFILLER_1_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5389_ _7205_/Q vssd1 vssd1 vccd1 vccd1 _5493_/A sky130_fd_sc_hd__buf_2
X_4409_ _4408_/X _7481_/Q _4409_/S vssd1 vssd1 vccd1 vccd1 _4410_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7128_ _7372_/CLK _7128_/D vssd1 vssd1 vccd1 vccd1 _7128_/Q sky130_fd_sc_hd__dfxtp_1
X_7059_ _7059_/A vssd1 vssd1 vccd1 vccd1 _7842_/D sky130_fd_sc_hd__clkbuf_1
X_5361__192 _5362__193/A vssd1 vssd1 vccd1 vccd1 _7164_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6346__428 _6347__429/A vssd1 vssd1 vccd1 vccd1 _7491_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _4760_/A vssd1 vssd1 vccd1 vccd1 _7296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3711_ _3711_/A vssd1 vssd1 vccd1 vccd1 _7749_/D sky130_fd_sc_hd__clkbuf_1
X_4691_ _4399_/X _7323_/Q _4697_/S vssd1 vssd1 vccd1 vccd1 _4692_/A sky130_fd_sc_hd__mux2_1
X_3642_ _3642_/A vssd1 vssd1 vccd1 vccd1 _7772_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3142_ clkbuf_0__3142_/X vssd1 vssd1 vccd1 vccd1 _6525__89/A sky130_fd_sc_hd__clkbuf_4
X_6361_ _6373_/A vssd1 vssd1 vccd1 vccd1 _6361_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_0__f__3296_ clkbuf_0__3296_/X vssd1 vssd1 vccd1 vccd1 _6751__139/A sky130_fd_sc_hd__clkbuf_16
XFILLER_115_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5312_ _5311_/X _7344_/Q _5307_/X _5308_/X _7144_/Q vssd1 vssd1 vccd1 vccd1 _7144_/D
+ sky130_fd_sc_hd__o32a_1
X_3573_ _7823_/Q vssd1 vssd1 vccd1 vccd1 _3947_/A sky130_fd_sc_hd__buf_2
XFILLER_114_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5243_ _7342_/Q _7341_/Q _7344_/Q _7343_/Q vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__and4_1
Xclkbuf_0__3110_ _6361_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3110_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_114_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5174_ _5236_/B vssd1 vssd1 vccd1 vccd1 _5185_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_68_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4125_ _3832_/X _7581_/Q _4129_/S vssd1 vssd1 vccd1 vccd1 _4126_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5792__257 _5792__257/A vssd1 vssd1 vccd1 vccd1 _7274_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4056_ _4056_/A vssd1 vssd1 vccd1 vccd1 _7608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7815_ _7819_/CLK _7815_/D vssd1 vssd1 vccd1 vccd1 _7815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7746_ _7746_/CLK _7746_/D vssd1 vssd1 vccd1 vccd1 _7746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4958_ _4958_/A vssd1 vssd1 vccd1 vccd1 _7167_/D sky130_fd_sc_hd__clkbuf_1
X_7677_ _7679_/CLK _7677_/D vssd1 vssd1 vccd1 vccd1 _7677_/Q sky130_fd_sc_hd__dfxtp_1
X_4889_ _4811_/X _7242_/Q _4893_/S vssd1 vssd1 vccd1 vccd1 _4890_/A sky130_fd_sc_hd__mux2_1
X_3909_ _3924_/S vssd1 vssd1 vccd1 vccd1 _3918_/S sky130_fd_sc_hd__buf_2
X_6628_ _7684_/Q _6711_/B vssd1 vssd1 vccd1 vccd1 _6714_/B sky130_fd_sc_hd__xor2_1
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6559_ _6573_/A vssd1 vssd1 vccd1 vccd1 _6594_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3308_ _6808_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3308_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_86_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5368__198 _5368__198/A vssd1 vssd1 vccd1 vccd1 _7170_/CLK sky130_fd_sc_hd__inv_2
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5930_ _6394_/A _6328_/C _6714_/A vssd1 vssd1 vccd1 vccd1 _6631_/B sky130_fd_sc_hd__and3_2
XFILLER_18_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5861_ _5861_/A vssd1 vssd1 vccd1 vccd1 _7326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7600_ _7600_/CLK _7600_/D vssd1 vssd1 vccd1 vccd1 _7600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4812_ _4811_/X _7274_/Q _4818_/S vssd1 vssd1 vccd1 vccd1 _4813_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7531_ _7531_/CLK _7531_/D vssd1 vssd1 vccd1 vccd1 _7531_/Q sky130_fd_sc_hd__dfxtp_1
X_4743_ _4722_/X _7303_/Q _4747_/S vssd1 vssd1 vccd1 vccd1 _4744_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7462_ _7462_/CLK _7462_/D vssd1 vssd1 vccd1 vccd1 _7462_/Q sky130_fd_sc_hd__dfxtp_1
X_4674_ _3660_/X _7354_/Q _4678_/S vssd1 vssd1 vccd1 vccd1 _4675_/A sky130_fd_sc_hd__mux2_1
X_6413_ _6413_/A vssd1 vssd1 vccd1 vccd1 _6413_/X sky130_fd_sc_hd__buf_1
X_7393_ _7393_/CLK _7393_/D vssd1 vssd1 vccd1 vccd1 _7393_/Q sky130_fd_sc_hd__dfxtp_1
X_3625_ _3625_/A vssd1 vssd1 vccd1 vccd1 _7779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3556_ _3556_/A vssd1 vssd1 vccd1 vccd1 _7836_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3125_ clkbuf_0__3125_/X vssd1 vssd1 vccd1 vccd1 _6443__504/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5226_ _5217_/X _5226_/B vssd1 vssd1 vccd1 vccd1 _5226_/X sky130_fd_sc_hd__and2b_1
X_5157_ _7187_/Q _5161_/B _5215_/A vssd1 vssd1 vccd1 vccd1 _5157_/X sky130_fd_sc_hd__and3_1
XFILLER_96_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5088_ _5088_/A vssd1 vssd1 vccd1 vccd1 _5088_/X sky130_fd_sc_hd__clkbuf_1
X_4108_ _4194_/A vssd1 vssd1 vccd1 vccd1 _4150_/B sky130_fd_sc_hd__inv_2
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4039_ _4039_/A vssd1 vssd1 vccd1 vccd1 _7614_/D sky130_fd_sc_hd__clkbuf_1
X_7035__54 _7035__54/A vssd1 vssd1 vccd1 vccd1 _7833_/CLK sky130_fd_sc_hd__inv_2
X_6779__161 _6779__161/A vssd1 vssd1 vccd1 vccd1 _7728_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6126__341 _6127__342/A vssd1 vssd1 vccd1 vccd1 _7390_/CLK sky130_fd_sc_hd__inv_2
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7729_ _7729_/CLK _7729_/D vssd1 vssd1 vccd1 vccd1 _7729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6849__43 _6850__44/A vssd1 vssd1 vccd1 vccd1 _7785_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2987_ clkbuf_0__2987_/X vssd1 vssd1 vccd1 vccd1 _6127__342/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6359__438 _6359__438/A vssd1 vssd1 vccd1 vccd1 _7501_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4390_ _4390_/A vssd1 vssd1 vccd1 vccd1 _7487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _6056_/X _6057_/X _6058_/X _6059_/X _5953_/X _5947_/X vssd1 vssd1 vccd1 vccd1
+ _6060_/X sky130_fd_sc_hd__mux4_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _5068_/A vssd1 vssd1 vccd1 vccd1 _5081_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_78_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6962_ _6960_/Y _6961_/X _6954_/X vssd1 vssd1 vccd1 vccd1 _7807_/D sky130_fd_sc_hd__a21oi_1
X_5913_ _5925_/A vssd1 vssd1 vccd1 vccd1 _5913_/X sky130_fd_sc_hd__buf_1
X_6893_ _6893_/A _6893_/B _6893_/C _6892_/X vssd1 vssd1 vccd1 vccd1 _6893_/X sky130_fd_sc_hd__or4b_1
XFILLER_34_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7514_ _7514_/CLK _7514_/D vssd1 vssd1 vccd1 vccd1 _7514_/Q sky130_fd_sc_hd__dfxtp_1
X_4726_ _4725_/X _7310_/Q _4729_/S vssd1 vssd1 vccd1 vccd1 _4727_/A sky130_fd_sc_hd__mux2_1
X_4657_ _4657_/A vssd1 vssd1 vccd1 vccd1 _7362_/D sky130_fd_sc_hd__clkbuf_1
X_7445_ _7445_/CLK _7445_/D vssd1 vssd1 vccd1 vccd1 _7445_/Q sky130_fd_sc_hd__dfxtp_1
X_7376_ _7376_/CLK _7376_/D vssd1 vssd1 vccd1 vccd1 _7376_/Q sky130_fd_sc_hd__dfxtp_1
X_3608_ _3578_/X _7785_/Q _3608_/S vssd1 vssd1 vccd1 vccd1 _3609_/A sky130_fd_sc_hd__mux2_1
Xinput80 wbs_data_i[4] vssd1 vssd1 vccd1 vccd1 _7024_/A sky130_fd_sc_hd__buf_8
Xinput91 wbs_we_i vssd1 vssd1 vccd1 vccd1 _4998_/A sky130_fd_sc_hd__buf_12
X_4588_ _7400_/Q _3941_/A _4588_/S vssd1 vssd1 vccd1 vccd1 _4589_/A sky130_fd_sc_hd__mux2_1
X_6327_ _6327_/A vssd1 vssd1 vccd1 vccd1 _7476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3539_ _3678_/A _3585_/A vssd1 vssd1 vccd1 vccd1 _3927_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_1_0_0__2772_ clkbuf_0__2772_/X vssd1 vssd1 vccd1 vccd1 _5805__267/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6258_ _7812_/Q _7811_/Q vssd1 vssd1 vccd1 vccd1 _6259_/B sky130_fd_sc_hd__nand2_1
X_5209_ _5206_/X _5209_/B vssd1 vssd1 vccd1 vccd1 _5209_/X sky130_fd_sc_hd__and2b_1
XFILLER_103_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6189_ _6189_/A _6888_/B vssd1 vssd1 vccd1 vccd1 _6866_/A sky130_fd_sc_hd__xor2_1
XFILLER_29_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5254__184 _5254__184/A vssd1 vssd1 vccd1 vccd1 _7113_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6471__526 _6471__526/A vssd1 vssd1 vccd1 vccd1 _7591_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6760__146 _6760__146/A vssd1 vssd1 vccd1 vccd1 _7713_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3890_ _3905_/S vssd1 vssd1 vccd1 vccd1 _3899_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5560_ _5550_/X _5553_/X _5556_/X _5559_/X _5404_/X _5602_/S vssd1 vssd1 vccd1 vccd1
+ _5560_/X sky130_fd_sc_hd__mux4_2
XFILLER_117_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5491_ _5491_/A _5493_/D _7040_/C vssd1 vssd1 vccd1 vccd1 _5492_/B sky130_fd_sc_hd__or3_1
X_4511_ _7438_/Q _4224_/X _4515_/S vssd1 vssd1 vccd1 vccd1 _4512_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4442_ _6002_/A vssd1 vssd1 vccd1 vccd1 _5998_/A sky130_fd_sc_hd__clkbuf_2
X_6525__89 _6525__89/A vssd1 vssd1 vccd1 vccd1 _7634_/CLK sky130_fd_sc_hd__inv_2
X_7230_ _7230_/CLK _7230_/D vssd1 vssd1 vccd1 vccd1 _7230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7161_ _7161_/CLK _7161_/D vssd1 vssd1 vccd1 vccd1 _7161_/Q sky130_fd_sc_hd__dfxtp_1
X_4373_ _4173_/X _7494_/Q _4373_/S vssd1 vssd1 vccd1 vccd1 _4374_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7092_ _7092_/A _7092_/B vssd1 vssd1 vccd1 vccd1 _7092_/Y sky130_fd_sc_hd__nand2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6043_ _7757_/Q _7749_/Q _7741_/Q _7655_/Q _6024_/X _5940_/X vssd1 vssd1 vccd1 vccd1
+ _6043_/X sky130_fd_sc_hd__mux4_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6843__38 _6844__39/A vssd1 vssd1 vccd1 vccd1 _7780_/CLK sky130_fd_sc_hd__inv_2
XFILLER_100_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6945_ _6942_/Y _6944_/X _6935_/X vssd1 vssd1 vccd1 vccd1 _7802_/D sky130_fd_sc_hd__a21oi_1
XFILLER_54_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7474_/CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_41_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6876_ _6242_/A _6249_/B _6873_/Y _6874_/X _6875_/X vssd1 vssd1 vccd1 vccd1 _6893_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_50_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5827_ _6269_/A vssd1 vssd1 vccd1 vccd1 _5827_/X sky130_fd_sc_hd__buf_1
XFILLER_10_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5758_ _5758_/A vssd1 vssd1 vccd1 vccd1 _5758_/X sky130_fd_sc_hd__buf_1
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4709_ _4709_/A vssd1 vssd1 vccd1 vccd1 _7316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7428_ _7428_/CLK _7428_/D vssd1 vssd1 vccd1 vccd1 _7428_/Q sky130_fd_sc_hd__dfxtp_1
X_5689_ _5689_/A vssd1 vssd1 vccd1 vccd1 _7206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7359_ _7359_/CLK _7359_/D vssd1 vssd1 vccd1 vccd1 _7359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3307_ clkbuf_0__3307_/X vssd1 vssd1 vccd1 vccd1 _6807__9/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5813__274 _5813__274/A vssd1 vssd1 vccd1 vccd1 _7291_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6436__498 _6437__499/A vssd1 vssd1 vccd1 vccd1 _7563_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4991_ _7108_/Q _5144_/A vssd1 vssd1 vccd1 vccd1 _5177_/A sky130_fd_sc_hd__nor2_4
XFILLER_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3942_ _3941_/X _7654_/Q _3942_/S vssd1 vssd1 vccd1 vccd1 _3943_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6661_ _6684_/A vssd1 vssd1 vccd1 vccd1 _6661_/X sky130_fd_sc_hd__clkbuf_2
X_3873_ _3873_/A vssd1 vssd1 vccd1 vccd1 _7703_/D sky130_fd_sc_hd__clkbuf_1
X_6592_ _6595_/A _6595_/B _6613_/A _7675_/Q vssd1 vssd1 vccd1 vccd1 _6593_/B sky130_fd_sc_hd__a31o_1
X_5612_ _7244_/Q _7175_/Q _7485_/Q _7252_/Q _4297_/A _5427_/X vssd1 vssd1 vccd1 vccd1
+ _5613_/B sky130_fd_sc_hd__mux4_1
XFILLER_31_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5543_ _5492_/Y _5542_/X _5493_/X vssd1 vssd1 vccd1 vccd1 _5543_/X sky130_fd_sc_hd__a21o_1
X_5474_ _5516_/A vssd1 vssd1 vccd1 vccd1 _5569_/S sky130_fd_sc_hd__buf_2
X_7213_ _7333_/CLK _7213_/D vssd1 vssd1 vccd1 vccd1 _7213_/Q sky130_fd_sc_hd__dfxtp_1
X_4425_ _4423_/Y _3973_/B _4424_/X _4131_/A _4421_/X vssd1 vssd1 vccd1 vccd1 _7466_/D
+ sky130_fd_sc_hd__o221a_1
X_7144_ _7348_/CLK _7144_/D vssd1 vssd1 vccd1 vccd1 _7144_/Q sky130_fd_sc_hd__dfxtp_1
X_4356_ _4356_/A vssd1 vssd1 vccd1 vccd1 _7502_/D sky130_fd_sc_hd__clkbuf_1
X_6153__359 _6153__359/A vssd1 vssd1 vccd1 vccd1 _7411_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6816__16 _6818__18/A vssd1 vssd1 vccd1 vccd1 _7758_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7075_ _7070_/X _7075_/B vssd1 vssd1 vccd1 vccd1 _7076_/A sky130_fd_sc_hd__and2b_1
X_4287_ _4287_/A vssd1 vssd1 vccd1 vccd1 _7523_/D sky130_fd_sc_hd__clkbuf_1
X_5756__228 _5757__229/A vssd1 vssd1 vccd1 vccd1 _7245_/CLK sky130_fd_sc_hd__inv_2
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6026_ _6021_/X _6022_/X _6023_/X _6025_/X _5945_/X _4436_/X vssd1 vssd1 vccd1 vccd1
+ _6026_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7869__196 vssd1 vssd1 vccd1 vccd1 _7869__196/HI core0Index[3] sky130_fd_sc_hd__conb_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__2987_ _6124_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2987_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_81_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6928_ _6924_/X _6907_/X _6881_/B vssd1 vssd1 vccd1 vccd1 _6928_/X sky130_fd_sc_hd__a21o_1
X_6859_ _6859_/A _7793_/Q vssd1 vssd1 vccd1 vccd1 _6897_/A sky130_fd_sc_hd__or2_1
XFILLER_50_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4210_ _4210_/A vssd1 vssd1 vccd1 vccd1 _7548_/D sky130_fd_sc_hd__clkbuf_1
X_5190_ _7131_/Q _5187_/X input8/X _5177_/X _5189_/X vssd1 vssd1 vccd1 vccd1 _5190_/X
+ sky130_fd_sc_hd__a221o_4
X_4141_ _4060_/X _7574_/Q _4141_/S vssd1 vssd1 vccd1 vccd1 _4142_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4072_ _4243_/B _4072_/B vssd1 vssd1 vccd1 vccd1 _4088_/S sky130_fd_sc_hd__or2_2
XFILLER_95_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7831_ _7831_/CLK _7831_/D vssd1 vssd1 vccd1 vccd1 _7831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7762_ _7762_/CLK _7762_/D vssd1 vssd1 vccd1 vccd1 _7762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4974_ _4974_/A vssd1 vssd1 vccd1 vccd1 _7116_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6713_ _6679_/A _6684_/A _7684_/Q vssd1 vssd1 vccd1 vccd1 _6713_/X sky130_fd_sc_hd__a21bo_1
X_7693_ _7693_/CLK _7693_/D vssd1 vssd1 vccd1 vccd1 _7693_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2772_ _5802_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2772_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_32_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3925_ _3925_/A vssd1 vssd1 vccd1 vccd1 _7661_/D sky130_fd_sc_hd__clkbuf_1
X_6773__156 _6773__156/A vssd1 vssd1 vccd1 vccd1 _7723_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3856_ _3856_/A vssd1 vssd1 vccd1 vccd1 _7707_/D sky130_fd_sc_hd__clkbuf_1
X_6120__336 _6122__338/A vssd1 vssd1 vccd1 vccd1 _7385_/CLK sky130_fd_sc_hd__inv_2
X_6575_ _6696_/B _6696_/C _6576_/A vssd1 vssd1 vccd1 vccd1 _6588_/A sky130_fd_sc_hd__a21o_1
X_3787_ _7523_/Q _7518_/Q vssd1 vssd1 vccd1 vccd1 _3787_/X sky130_fd_sc_hd__or2b_1
XFILLER_118_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5526_ _7528_/Q _5463_/Y _5525_/X _5495_/X vssd1 vssd1 vccd1 vccd1 _5526_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5457_ _5457_/A vssd1 vssd1 vccd1 vccd1 _5457_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4408_ _4408_/A vssd1 vssd1 vccd1 vccd1 _4408_/X sky130_fd_sc_hd__buf_2
XFILLER_87_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5388_ _5388_/A vssd1 vssd1 vccd1 vccd1 _7040_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_101_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7127_ _7329_/CLK _7127_/D vssd1 vssd1 vccd1 vccd1 _7127_/Q sky130_fd_sc_hd__dfxtp_1
X_4339_ _4767_/A _4505_/C vssd1 vssd1 vccd1 vccd1 _4355_/S sky130_fd_sc_hd__nand2_4
XFILLER_101_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7058_ _7048_/X _7058_/B vssd1 vssd1 vccd1 vccd1 _7059_/A sky130_fd_sc_hd__and2b_1
XFILLER_59_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6009_ _6099_/A _6009_/B vssd1 vssd1 vccd1 vccd1 _6009_/X sky130_fd_sc_hd__or2_1
XFILLER_74_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6286__398 _6286__398/A vssd1 vssd1 vccd1 vccd1 _7451_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _3709_/X _7749_/Q _3713_/S vssd1 vssd1 vccd1 vccd1 _3711_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4690_ _4690_/A vssd1 vssd1 vccd1 vccd1 _7324_/D sky130_fd_sc_hd__clkbuf_1
X_3641_ _3566_/X _7772_/Q _3641_/S vssd1 vssd1 vccd1 vccd1 _3642_/A sky130_fd_sc_hd__mux2_1
X_3572_ _3572_/A vssd1 vssd1 vccd1 vccd1 _7832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3141_ clkbuf_0__3141_/X vssd1 vssd1 vccd1 vccd1 _6519__84/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5311_ _7070_/A vssd1 vssd1 vccd1 vccd1 _5311_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5242_ _7070_/A vssd1 vssd1 vccd1 vccd1 _5245_/B sky130_fd_sc_hd__clkbuf_4
X_5173_ _5187_/A vssd1 vssd1 vccd1 vccd1 _5173_/X sky130_fd_sc_hd__buf_2
XFILLER_96_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4124_ _4124_/A vssd1 vssd1 vccd1 vccd1 _7582_/D sky130_fd_sc_hd__clkbuf_1
Xinput1 caravel_uart_rx vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4055_ _4054_/X _7608_/Q _4061_/S vssd1 vssd1 vccd1 vccd1 _4056_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6306__413 _6306__413/A vssd1 vssd1 vccd1 vccd1 _7466_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7814_ _7819_/CLK _7814_/D vssd1 vssd1 vccd1 vccd1 _7814_/Q sky130_fd_sc_hd__dfxtp_1
X_7745_ _7745_/CLK _7745_/D vssd1 vssd1 vccd1 vccd1 _7745_/Q sky130_fd_sc_hd__dfxtp_1
X_4957_ _4213_/X _7167_/Q _4965_/S vssd1 vssd1 vccd1 vccd1 _4958_/A sky130_fd_sc_hd__mux2_1
X_7676_ _7680_/CLK _7676_/D vssd1 vssd1 vccd1 vccd1 _7676_/Q sky130_fd_sc_hd__dfxtp_1
X_4888_ _4888_/A vssd1 vssd1 vccd1 vccd1 _7243_/D sky130_fd_sc_hd__clkbuf_1
X_3908_ _4919_/B _4706_/A vssd1 vssd1 vccd1 vccd1 _3924_/S sky130_fd_sc_hd__or2_2
X_6627_ _6189_/A _6708_/B _6612_/Y _6616_/X _6626_/X vssd1 vssd1 vccd1 vccd1 _6652_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_20_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3839_ _7468_/Q vssd1 vssd1 vccd1 vccd1 _4417_/A sky130_fd_sc_hd__buf_2
X_6558_ _7672_/Q _7671_/Q _7670_/Q _7669_/Q vssd1 vssd1 vccd1 vccd1 _6573_/A sky130_fd_sc_hd__and4_1
XFILLER_105_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5509_ _7690_/Q _7279_/Q _7162_/Q _7271_/Q _5472_/A _5508_/X vssd1 vssd1 vccd1 vccd1
+ _5509_/X sky130_fd_sc_hd__mux4_1
X_6352__433 _6353__434/A vssd1 vssd1 vccd1 vccd1 _7496_/CLK sky130_fd_sc_hd__inv_2
X_6489_ _6507_/A vssd1 vssd1 vccd1 vccd1 _6489_/X sky130_fd_sc_hd__buf_1
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3307_ _6802_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3307_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_79_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7884__211 vssd1 vssd1 vccd1 vccd1 _7884__211/HI manufacturerID[3] sky130_fd_sc_hd__conb_1
XFILLER_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2452_ clkbuf_0__2452_/X vssd1 vssd1 vccd1 vccd1 _5739__214/A sky130_fd_sc_hd__clkbuf_16
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6166__369 _6166__369/A vssd1 vssd1 vccd1 vccd1 _7421_/CLK sky130_fd_sc_hd__inv_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5769__238 _5769__238/A vssd1 vssd1 vccd1 vccd1 _7255_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5860_ _5033_/A hold2/A _5866_/S vssd1 vssd1 vccd1 vccd1 _5861_/A sky130_fd_sc_hd__mux2_1
X_4811_ _7473_/Q vssd1 vssd1 vccd1 vccd1 _4811_/X sky130_fd_sc_hd__buf_2
XFILLER_33_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7530_ _7855_/CLK _7530_/D vssd1 vssd1 vccd1 vccd1 _7530_/Q sky130_fd_sc_hd__dfxtp_1
X_4742_ _4742_/A vssd1 vssd1 vccd1 vccd1 _7304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4673_ _4673_/A vssd1 vssd1 vccd1 vccd1 _7355_/D sky130_fd_sc_hd__clkbuf_1
X_7461_ _7461_/CLK _7461_/D vssd1 vssd1 vccd1 vccd1 _7461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3624_ _3570_/X _7779_/Q _3628_/S vssd1 vssd1 vccd1 vccd1 _3625_/A sky130_fd_sc_hd__mux2_1
X_7392_ _7392_/CLK _7392_/D vssd1 vssd1 vccd1 vccd1 _7392_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3124_ clkbuf_0__3124_/X vssd1 vssd1 vccd1 vccd1 _6435__497/A sky130_fd_sc_hd__clkbuf_4
X_3555_ _3554_/X _7836_/Q _3567_/S vssd1 vssd1 vccd1 vccd1 _3556_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5225_ _7143_/Q _5215_/X _5216_/X _5224_/X vssd1 vssd1 vccd1 vccd1 _5225_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5156_ _7119_/Q _5145_/X input25/X _5146_/X _5155_/X vssd1 vssd1 vccd1 vccd1 _5156_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_96_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5087_ _5087_/A _5087_/B vssd1 vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__and2_1
XFILLER_111_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4107_ _4107_/A vssd1 vssd1 vccd1 vccd1 _7587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4038_ _3941_/X _7614_/Q _4038_/S vssd1 vssd1 vccd1 vccd1 _4039_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _7588_/Q _7556_/Q _7831_/Q _7532_/Q _6002_/A _5956_/X vssd1 vssd1 vccd1 vccd1
+ _5990_/B sky130_fd_sc_hd__mux4_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7728_ _7728_/CLK _7728_/D vssd1 vssd1 vccd1 vccd1 _7728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7659_ _7687_/CLK _7659_/D vssd1 vssd1 vccd1 vccd1 _7659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2986_ clkbuf_0__2986_/X vssd1 vssd1 vccd1 vccd1 _6122__338/A sky130_fd_sc_hd__clkbuf_4
XFILLER_4_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput190 _5170_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[7] sky130_fd_sc_hd__buf_2
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5010_ _7105_/A vssd1 vssd1 vccd1 vccd1 _7016_/A sky130_fd_sc_hd__buf_6
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6961_ _6912_/X _6919_/X _6195_/B vssd1 vssd1 vccd1 vccd1 _6961_/X sky130_fd_sc_hd__a21o_1
X_5912_ _6117_/A vssd1 vssd1 vccd1 vccd1 _5912_/X sky130_fd_sc_hd__buf_1
X_6892_ _6972_/A _6892_/B _6892_/C _6892_/D vssd1 vssd1 vccd1 vccd1 _6892_/X sky130_fd_sc_hd__and4_1
XFILLER_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7513_ _7513_/CLK _7513_/D vssd1 vssd1 vccd1 vccd1 _7513_/Q sky130_fd_sc_hd__dfxtp_1
X_4725_ _7469_/Q vssd1 vssd1 vccd1 vccd1 _4725_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4656_ _4402_/X _7362_/Q _4660_/S vssd1 vssd1 vccd1 vccd1 _4657_/A sky130_fd_sc_hd__mux2_1
X_7444_ _7444_/CLK _7444_/D vssd1 vssd1 vccd1 vccd1 _7444_/Q sky130_fd_sc_hd__dfxtp_1
X_4587_ _4587_/A vssd1 vssd1 vccd1 vccd1 _7401_/D sky130_fd_sc_hd__clkbuf_1
X_7375_ _7375_/CLK _7375_/D vssd1 vssd1 vccd1 vccd1 _7375_/Q sky130_fd_sc_hd__dfxtp_1
X_3607_ _3607_/A vssd1 vssd1 vccd1 vccd1 _7786_/D sky130_fd_sc_hd__clkbuf_1
Xinput81 wbs_data_i[5] vssd1 vssd1 vccd1 vccd1 _7026_/A sky130_fd_sc_hd__buf_8
Xinput70 wbs_data_i[24] vssd1 vssd1 vccd1 vccd1 _5066_/A sky130_fd_sc_hd__buf_4
XFILLER_115_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6326_ _6326_/A _6326_/B _7030_/B vssd1 vssd1 vccd1 vccd1 _6327_/A sky130_fd_sc_hd__and3_1
X_3538_ _7465_/Q _5932_/A _4448_/B _4424_/B vssd1 vssd1 vccd1 vccd1 _3545_/B sky130_fd_sc_hd__o211ai_1
Xclkbuf_1_1_0__3107_ clkbuf_0__3107_/X vssd1 vssd1 vccd1 vccd1 _6349__430/A sky130_fd_sc_hd__clkbuf_4
XFILLER_107_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2771_ clkbuf_0__2771_/X vssd1 vssd1 vccd1 vccd1 _5801__264/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6257_ _7813_/Q vssd1 vssd1 vccd1 vccd1 _6259_/A sky130_fd_sc_hd__inv_2
X_5208_ _7136_/Q _5199_/X _5204_/X _5207_/X vssd1 vssd1 vccd1 vccd1 _5208_/X sky130_fd_sc_hd__o22a_4
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6188_ _7808_/Q _6188_/B vssd1 vssd1 vccd1 vccd1 _6888_/B sky130_fd_sc_hd__xnor2_2
X_5139_ _5139_/A vssd1 vssd1 vccd1 vccd1 _5139_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5839__294 _5839__294/A vssd1 vssd1 vccd1 vccd1 _7311_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_8_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7839_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6365__443 _6366__444/A vssd1 vssd1 vccd1 vccd1 _7506_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4510_ _4510_/A vssd1 vssd1 vccd1 vccd1 _7439_/D sky130_fd_sc_hd__clkbuf_1
X_5490_ _5602_/S _5470_/X _5477_/X _5489_/X vssd1 vssd1 vccd1 vccd1 _5490_/X sky130_fd_sc_hd__a31o_1
XFILLER_117_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4441_ _5936_/A vssd1 vssd1 vccd1 vccd1 _6002_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7160_ _7160_/CLK _7160_/D vssd1 vssd1 vccd1 vccd1 _7160_/Q sky130_fd_sc_hd__dfxtp_1
X_6111_ _6111_/A vssd1 vssd1 vccd1 vccd1 _6111_/X sky130_fd_sc_hd__buf_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4372_ _4372_/A vssd1 vssd1 vccd1 vccd1 _7495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7091_ _7105_/C vssd1 vssd1 vccd1 vccd1 _7104_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6042_ _7725_/Q _7709_/Q _7428_/Q _7490_/Q _5935_/X _5974_/X vssd1 vssd1 vccd1 vccd1
+ _6042_/X sky130_fd_sc_hd__mux4_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6944_ _6943_/X _6939_/X _6873_/B vssd1 vssd1 vccd1 vccd1 _6944_/X sky130_fd_sc_hd__a21o_1
XFILLER_81_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6875_ _7844_/Q _6249_/B _6247_/B _6249_/A vssd1 vssd1 vccd1 vccd1 _6875_/X sky130_fd_sc_hd__a2bb2o_1
X_5826_ _6300_/A vssd1 vssd1 vccd1 vccd1 _5826_/X sky130_fd_sc_hd__buf_1
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4708_ _4705_/X _7316_/Q _4720_/S vssd1 vssd1 vccd1 vccd1 _4709_/A sky130_fd_sc_hd__mux2_1
X_7427_ _7427_/CLK _7427_/D vssd1 vssd1 vccd1 vccd1 _7427_/Q sky130_fd_sc_hd__dfxtp_1
X_5688_ _7206_/Q _5092_/A _5692_/S vssd1 vssd1 vccd1 vccd1 _5689_/A sky130_fd_sc_hd__mux2_1
X_4639_ _4639_/A vssd1 vssd1 vccd1 vccd1 _7378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7358_ _7358_/CLK _7358_/D vssd1 vssd1 vccd1 vccd1 _7358_/Q sky130_fd_sc_hd__dfxtp_1
X_7289_ _7289_/CLK _7289_/D vssd1 vssd1 vccd1 vccd1 _7289_/Q sky130_fd_sc_hd__dfxtp_1
X_6309_ _6309_/A vssd1 vssd1 vccd1 vccd1 _7468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3306_ clkbuf_0__3306_/X vssd1 vssd1 vccd1 vccd1 _6814_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6139__352 _6141__354/A vssd1 vssd1 vccd1 vccd1 _7401_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6530__93 _6531__94/A vssd1 vssd1 vccd1 vccd1 _7638_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4990_ _5149_/A vssd1 vssd1 vccd1 vccd1 _5144_/A sky130_fd_sc_hd__inv_2
XFILLER_91_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3941_ _3941_/A vssd1 vssd1 vccd1 vccd1 _3941_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_16_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6660_ _6583_/B _6711_/D _6659_/Y _5996_/A vssd1 vssd1 vccd1 vccd1 _7669_/D sky130_fd_sc_hd__o211a_1
X_3872_ _3816_/X _7703_/Q _3878_/S vssd1 vssd1 vccd1 vccd1 _3873_/A sky130_fd_sc_hd__mux2_1
X_6591_ _7675_/Q _6595_/A _6595_/B _6613_/A vssd1 vssd1 vccd1 vccd1 _6593_/A sky130_fd_sc_hd__nand4_1
X_5611_ _5609_/X _5610_/X _5611_/S vssd1 vssd1 vccd1 vccd1 _5611_/X sky130_fd_sc_hd__mux2_2
XFILLER_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5542_ _5532_/X _5535_/X _5538_/X _5541_/X _5404_/X _5602_/S vssd1 vssd1 vccd1 vccd1
+ _5542_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5473_ _7238_/Q _7169_/Q _7479_/Q _7246_/Q _5472_/X _5427_/X vssd1 vssd1 vccd1 vccd1
+ _5473_/X sky130_fd_sc_hd__mux4_1
X_7212_ _7333_/CLK _7212_/D vssd1 vssd1 vccd1 vccd1 _7212_/Q sky130_fd_sc_hd__dfxtp_1
X_4424_ _4424_/A _4424_/B _4424_/C vssd1 vssd1 vccd1 vccd1 _4424_/X sky130_fd_sc_hd__and3_1
X_7143_ _7344_/CLK _7143_/D vssd1 vssd1 vccd1 vccd1 _7143_/Q sky130_fd_sc_hd__dfxtp_1
X_4355_ _4173_/X _7502_/Q _4355_/S vssd1 vssd1 vccd1 vccd1 _4356_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7074_ _5031_/A _7847_/Q _7074_/S vssd1 vssd1 vccd1 vccd1 _7075_/B sky130_fd_sc_hd__mux2_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4286_ _6394_/C _4286_/B _4286_/C vssd1 vssd1 vccd1 vccd1 _4287_/A sky130_fd_sc_hd__and3_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6025_ _7756_/Q _7748_/Q _7740_/Q _7654_/Q _6024_/X _5940_/X vssd1 vssd1 vccd1 vccd1
+ _6025_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2986_ _6118_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2986_/X sky130_fd_sc_hd__clkbuf_16
X_6927_ _7798_/Q _6933_/B vssd1 vssd1 vccd1 vccd1 _6927_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6789_ _6795_/A vssd1 vssd1 vccd1 vccd1 _6789_/X sky130_fd_sc_hd__buf_1
XFILLER_10_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5373__202 _5374__203/A vssd1 vssd1 vccd1 vccd1 _7174_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6503__71 _6504__72/A vssd1 vssd1 vccd1 vccd1 _7616_/CLK sky130_fd_sc_hd__inv_2
X_4140_ _4140_/A vssd1 vssd1 vccd1 vccd1 _7575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4071_ _4071_/A vssd1 vssd1 vccd1 vccd1 _7603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6821__20 _6822__21/A vssd1 vssd1 vccd1 vccd1 _7762_/CLK sky130_fd_sc_hd__inv_2
X_7830_ _7830_/CLK _7830_/D vssd1 vssd1 vccd1 vccd1 _7830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7761_ _7761_/CLK _7761_/D vssd1 vssd1 vccd1 vccd1 _7761_/Q sky130_fd_sc_hd__dfxtp_1
X_4973_ _7116_/Q _4393_/A _4979_/S vssd1 vssd1 vccd1 vccd1 _4974_/A sky130_fd_sc_hd__mux2_1
X_6712_ _6710_/X _6711_/Y _6690_/X vssd1 vssd1 vccd1 vccd1 _7683_/D sky130_fd_sc_hd__a21oi_1
X_7692_ _7692_/CLK _7692_/D vssd1 vssd1 vccd1 vccd1 _7692_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2771_ _5796_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2771_/X sky130_fd_sc_hd__clkbuf_16
X_3924_ _3840_/X _7661_/Q _3924_/S vssd1 vssd1 vccd1 vccd1 _3925_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6643_ _6731_/A vssd1 vssd1 vccd1 vccd1 _6643_/X sky130_fd_sc_hd__buf_1
X_3855_ _3715_/X _7707_/Q _3859_/S vssd1 vssd1 vccd1 vccd1 _3856_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6574_ _6602_/A _6621_/B _6621_/C _7678_/Q vssd1 vssd1 vccd1 vccd1 _6696_/C sky130_fd_sc_hd__a31o_1
X_3786_ _7523_/Q vssd1 vssd1 vccd1 vccd1 _4285_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7680_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5525_ _5492_/Y _5524_/X _5493_/X vssd1 vssd1 vccd1 vccd1 _5525_/X sky130_fd_sc_hd__a21o_1
X_5762__233 _5762__233/A vssd1 vssd1 vccd1 vccd1 _7250_/CLK sky130_fd_sc_hd__inv_2
X_5456_ _7405_/Q vssd1 vssd1 vccd1 vccd1 _6326_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4407_ _4407_/A vssd1 vssd1 vccd1 vccd1 _7482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5387_ _5446_/A vssd1 vssd1 vccd1 vccd1 _5682_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7126_ _7372_/CLK _7126_/D vssd1 vssd1 vccd1 vccd1 _7126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4338_ _4338_/A vssd1 vssd1 vccd1 vccd1 _7510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7057_ _5042_/A _6189_/A _7067_/S vssd1 vssd1 vccd1 vccd1 _7058_/B sky130_fd_sc_hd__mux2_1
X_4269_ _7528_/Q _7529_/Q _6308_/B vssd1 vssd1 vccd1 vccd1 _4270_/B sky130_fd_sc_hd__o21ai_1
XFILLER_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6008_ _7589_/Q _7557_/Q _7832_/Q _7533_/Q _5983_/X _5984_/X vssd1 vssd1 vccd1 vccd1
+ _6009_/B sky130_fd_sc_hd__mux4_1
XFILLER_67_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3640_ _3640_/A vssd1 vssd1 vccd1 vccd1 _7773_/D sky130_fd_sc_hd__clkbuf_1
X_3571_ _3570_/X _7832_/Q _3579_/S vssd1 vssd1 vccd1 vccd1 _3572_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3140_ clkbuf_0__3140_/X vssd1 vssd1 vccd1 vccd1 _6538_/A sky130_fd_sc_hd__clkbuf_4
X_5310_ _5303_/X _7343_/Q _5307_/X _5308_/X _7143_/Q vssd1 vssd1 vccd1 vccd1 _7143_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5241_ _5269_/A vssd1 vssd1 vccd1 vccd1 _7070_/A sky130_fd_sc_hd__clkbuf_4
X_5172_ _7125_/Q _5159_/X input33/X _5163_/X _5171_/X vssd1 vssd1 vccd1 vccd1 _5172_/X
+ sky130_fd_sc_hd__a221o_4
X_4123_ _3828_/X _7582_/Q _4123_/S vssd1 vssd1 vccd1 vccd1 _4124_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput2 caravel_wb_ack_i vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4054_ _7827_/Q vssd1 vssd1 vccd1 vccd1 _4054_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5833__289 _5833__289/A vssd1 vssd1 vccd1 vccd1 _7306_/CLK sky130_fd_sc_hd__inv_2
X_7813_ _7819_/CLK _7813_/D vssd1 vssd1 vccd1 vccd1 _7813_/Q sky130_fd_sc_hd__dfxtp_1
X_7744_ _7744_/CLK _7744_/D vssd1 vssd1 vccd1 vccd1 _7744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4956_ _4971_/S vssd1 vssd1 vccd1 vccd1 _4965_/S sky130_fd_sc_hd__buf_2
X_7675_ _7680_/CLK _7675_/D vssd1 vssd1 vccd1 vccd1 _7675_/Q sky130_fd_sc_hd__dfxtp_1
X_4887_ _4808_/X _7243_/Q _4893_/S vssd1 vssd1 vccd1 vccd1 _4888_/A sky130_fd_sc_hd__mux2_1
X_3907_ _7527_/Q _3907_/B _4111_/A vssd1 vssd1 vccd1 vccd1 _4706_/A sky130_fd_sc_hd__or3b_2
X_6626_ _6619_/X _6620_/Y _6623_/X _6624_/Y _6625_/X vssd1 vssd1 vccd1 vccd1 _6626_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3838_ _3838_/A vssd1 vssd1 vccd1 vccd1 _7714_/D sky130_fd_sc_hd__clkbuf_1
X_6557_ _7687_/Q _7660_/Q _6725_/D _7659_/Q vssd1 vssd1 vccd1 vccd1 _6630_/A sky130_fd_sc_hd__a31oi_2
XFILLER_20_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3769_ _3703_/X _7727_/Q _3775_/S vssd1 vssd1 vccd1 vccd1 _3770_/A sky130_fd_sc_hd__mux2_1
X_5508_ _5518_/A vssd1 vssd1 vccd1 vccd1 _5508_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3306_ _6801_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3306_/X sky130_fd_sc_hd__clkbuf_16
X_5439_ _5439_/A _5491_/A vssd1 vssd1 vccd1 vccd1 _5462_/D sky130_fd_sc_hd__or2_1
XFILLER_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7109_ _7109_/CLK _7109_/D vssd1 vssd1 vccd1 vccd1 _7109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4810_ _4810_/A vssd1 vssd1 vccd1 vccd1 _7275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4719_/X _7304_/Q _4741_/S vssd1 vssd1 vccd1 vccd1 _4742_/A sky130_fd_sc_hd__mux2_1
X_4672_ _3657_/X _7355_/Q _4678_/S vssd1 vssd1 vccd1 vccd1 _4673_/A sky130_fd_sc_hd__mux2_1
X_7460_ _7460_/CLK _7460_/D vssd1 vssd1 vccd1 vccd1 _7460_/Q sky130_fd_sc_hd__dfxtp_1
X_3623_ _3623_/A vssd1 vssd1 vccd1 vccd1 _7780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7391_ _7391_/CLK _7391_/D vssd1 vssd1 vccd1 vccd1 _7391_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3123_ clkbuf_0__3123_/X vssd1 vssd1 vccd1 vccd1 _6428__491/A sky130_fd_sc_hd__clkbuf_4
X_3554_ _3932_/A vssd1 vssd1 vccd1 vccd1 _3554_/X sky130_fd_sc_hd__buf_2
X_6342_ _6342_/A vssd1 vssd1 vccd1 vccd1 _6342_/X sky130_fd_sc_hd__buf_1
XFILLER_115_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5224_ _5217_/X _5224_/B vssd1 vssd1 vccd1 vccd1 _5224_/X sky130_fd_sc_hd__and2b_1
XFILLER_103_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5155_ _7186_/Q _5161_/B _5215_/A vssd1 vssd1 vccd1 vccd1 _5155_/X sky130_fd_sc_hd__and3_1
XFILLER_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5086_ _5086_/A vssd1 vssd1 vccd1 vccd1 _5086_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4106_ _4069_/X _7587_/Q _4106_/S vssd1 vssd1 vccd1 vccd1 _4107_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4037_ _4037_/A vssd1 vssd1 vccd1 vccd1 _7615_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _7786_/Q _7778_/Q _7770_/Q _7762_/Q _4446_/A _5954_/X vssd1 vssd1 vccd1 vccd1
+ _5988_/X sky130_fd_sc_hd__mux4_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__2769_ clkbuf_0__2769_/X vssd1 vssd1 vccd1 vccd1 _5794__259/A sky130_fd_sc_hd__clkbuf_4
X_7727_ _7727_/CLK _7727_/D vssd1 vssd1 vccd1 vccd1 _7727_/Q sky130_fd_sc_hd__dfxtp_1
X_4939_ _4213_/X _7175_/Q _4947_/S vssd1 vssd1 vccd1 vccd1 _4940_/A sky130_fd_sc_hd__mux2_1
X_7658_ _7658_/CLK _7658_/D vssd1 vssd1 vccd1 vccd1 _7658_/Q sky130_fd_sc_hd__dfxtp_1
X_6609_ _7682_/Q _6609_/B vssd1 vssd1 vccd1 vccd1 _6708_/B sky130_fd_sc_hd__xnor2_1
X_7589_ _7589_/CLK _7589_/D vssd1 vssd1 vccd1 vccd1 _7589_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__2985_ clkbuf_0__2985_/X vssd1 vssd1 vccd1 vccd1 _6130_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_opt_1_0_wb_clk_i _7826_/CLK vssd1 vssd1 vccd1 vccd1 _6481_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_4_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6786__167 _6788__169/A vssd1 vssd1 vccd1 vccd1 _7734_/CLK sky130_fd_sc_hd__inv_2
X_6172__374 _6172__374/A vssd1 vssd1 vccd1 vccd1 _7426_/CLK sky130_fd_sc_hd__inv_2
Xoutput180 _5227_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[27] sky130_fd_sc_hd__buf_2
Xoutput191 _5172_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[8] sky130_fd_sc_hd__buf_2
X_6133__347 _6133__347/A vssd1 vssd1 vccd1 vccd1 _7396_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5775__243 _5775__243/A vssd1 vssd1 vccd1 vccd1 _7260_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6441__502 _6442__503/A vssd1 vssd1 vccd1 vccd1 _7567_/CLK sky130_fd_sc_hd__inv_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6398__467 _6400__469/A vssd1 vssd1 vccd1 vccd1 _7532_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6537__99 _6537__99/A vssd1 vssd1 vccd1 vccd1 _7644_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6855__48 _6855__48/A vssd1 vssd1 vccd1 vccd1 _7790_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6960_ _7807_/Q _6969_/B vssd1 vssd1 vccd1 vccd1 _6960_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6891_ _7846_/Q _6883_/Y _6884_/Y _7849_/Q _6890_/X vssd1 vssd1 vccd1 vccd1 _6892_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2777_ clkbuf_0__2777_/X vssd1 vssd1 vccd1 vccd1 _5852_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7512_ _7512_/CLK _7512_/D vssd1 vssd1 vccd1 vccd1 _7512_/Q sky130_fd_sc_hd__dfxtp_1
X_4724_ _4724_/A vssd1 vssd1 vccd1 vccd1 _7311_/D sky130_fd_sc_hd__clkbuf_1
X_4655_ _4655_/A vssd1 vssd1 vccd1 vccd1 _7363_/D sky130_fd_sc_hd__clkbuf_1
X_7443_ _7443_/CLK _7443_/D vssd1 vssd1 vccd1 vccd1 _7443_/Q sky130_fd_sc_hd__dfxtp_1
X_7374_ _7374_/CLK _7374_/D vssd1 vssd1 vccd1 vccd1 _7374_/Q sky130_fd_sc_hd__dfxtp_1
X_4586_ _7401_/Q _3938_/A _4588_/S vssd1 vssd1 vccd1 vccd1 _4587_/A sky130_fd_sc_hd__mux2_1
X_3606_ _3574_/X _7786_/Q _3608_/S vssd1 vssd1 vccd1 vccd1 _3607_/A sky130_fd_sc_hd__mux2_1
Xinput82 wbs_data_i[6] vssd1 vssd1 vccd1 vccd1 _7028_/A sky130_fd_sc_hd__buf_8
Xinput60 wbs_data_i[15] vssd1 vssd1 vccd1 vccd1 _5047_/A sky130_fd_sc_hd__buf_6
Xinput71 wbs_data_i[25] vssd1 vssd1 vccd1 vccd1 _5069_/A sky130_fd_sc_hd__buf_4
XFILLER_115_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3106_ clkbuf_0__3106_/X vssd1 vssd1 vccd1 vccd1 _6343__425/A sky130_fd_sc_hd__clkbuf_4
X_6325_ _6325_/A _6325_/B vssd1 vssd1 vccd1 vccd1 _7030_/B sky130_fd_sc_hd__nor2_4
X_3537_ _7464_/Q _7463_/Q _7462_/Q vssd1 vssd1 vccd1 vccd1 _4424_/B sky130_fd_sc_hd__and3_1
Xclkbuf_1_0_0__2770_ clkbuf_0__2770_/X vssd1 vssd1 vccd1 vccd1 _5814_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6256_ _6859_/A _6900_/B vssd1 vssd1 vccd1 vccd1 _6978_/A sky130_fd_sc_hd__nor2_1
X_5207_ _5206_/X _5207_/B vssd1 vssd1 vccd1 vccd1 _5207_/X sky130_fd_sc_hd__and2b_1
XFILLER_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6187_ _5661_/X _6869_/A _6869_/B vssd1 vssd1 vccd1 vccd1 _6191_/A sky130_fd_sc_hd__nand3b_1
X_5138_ _5337_/C _7342_/Q _5138_/C _5138_/D vssd1 vssd1 vccd1 vccd1 _5139_/A sky130_fd_sc_hd__and4_1
XFILLER_57_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5069_ _5069_/A _5077_/B vssd1 vssd1 vccd1 vccd1 _5070_/A sky130_fd_sc_hd__or2_1
XFILLER_16_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6406__474 _6406__474/A vssd1 vssd1 vccd1 vccd1 _7539_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4440_ _7458_/Q vssd1 vssd1 vccd1 vccd1 _5936_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6828__26 _6828__26/A vssd1 vssd1 vccd1 vccd1 _7768_/CLK sky130_fd_sc_hd__inv_2
X_4371_ _4170_/X _7495_/Q _4373_/S vssd1 vssd1 vccd1 vccd1 _4372_/A sky130_fd_sc_hd__mux2_1
X_7090_ _7090_/A vssd1 vssd1 vccd1 vccd1 _7851_/D sky130_fd_sc_hd__clkbuf_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6041_ _7575_/Q _7385_/Q _7733_/Q _7631_/Q _6002_/X _4450_/A vssd1 vssd1 vccd1 vccd1
+ _6041_/X sky130_fd_sc_hd__mux4_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6448__508 _6448__508/A vssd1 vssd1 vccd1 vccd1 _7573_/CLK sky130_fd_sc_hd__inv_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6943_ _6943_/A vssd1 vssd1 vccd1 vccd1 _6943_/X sky130_fd_sc_hd__clkbuf_2
X_6874_ _7845_/Q _6247_/B _6195_/B _7842_/Q vssd1 vssd1 vccd1 vccd1 _6874_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_10_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5687_ _5687_/A vssd1 vssd1 vccd1 vccd1 _7205_/D sky130_fd_sc_hd__clkbuf_1
X_4707_ _4729_/S vssd1 vssd1 vccd1 vccd1 _4720_/S sky130_fd_sc_hd__buf_2
X_4638_ _3660_/X _7378_/Q _4642_/S vssd1 vssd1 vccd1 vccd1 _4639_/A sky130_fd_sc_hd__mux2_1
X_7426_ _7426_/CLK _7426_/D vssd1 vssd1 vccd1 vccd1 _7426_/Q sky130_fd_sc_hd__dfxtp_1
X_4569_ _4569_/A vssd1 vssd1 vccd1 vccd1 _7412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7357_ _7357_/CLK _7357_/D vssd1 vssd1 vccd1 vccd1 _7357_/Q sky130_fd_sc_hd__dfxtp_1
X_7288_ _7288_/CLK _7288_/D vssd1 vssd1 vccd1 vccd1 _7288_/Q sky130_fd_sc_hd__dfxtp_1
X_6308_ _7814_/Q _6308_/B vssd1 vssd1 vccd1 vccd1 _6309_/A sky130_fd_sc_hd__and2_1
X_6239_ _7804_/Q _7803_/Q vssd1 vssd1 vccd1 vccd1 _6245_/C sky130_fd_sc_hd__and2_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3305_ clkbuf_0__3305_/X vssd1 vssd1 vccd1 vccd1 _6798__177/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6291__402 _6292__403/A vssd1 vssd1 vccd1 vccd1 _7455_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6515__80 _6516__81/A vssd1 vssd1 vccd1 vccd1 _7625_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3940_ _3940_/A vssd1 vssd1 vccd1 vccd1 _7655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3871_ _3871_/A vssd1 vssd1 vccd1 vccd1 _7704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6590_ _7673_/Q vssd1 vssd1 vccd1 vccd1 _6595_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5610_ _7586_/Q _7570_/Q _7554_/Q _7546_/Q _5486_/X _5426_/X vssd1 vssd1 vccd1 vccd1
+ _5610_/X sky130_fd_sc_hd__mux4_1
X_5541_ _5539_/X _5540_/X _5578_/S vssd1 vssd1 vccd1 vccd1 _5541_/X sky130_fd_sc_hd__mux2_1
X_6454__512 _6455__513/A vssd1 vssd1 vccd1 vccd1 _7577_/CLK sky130_fd_sc_hd__inv_2
X_7211_ _5246_/A _7211_/D vssd1 vssd1 vccd1 vccd1 _7211_/Q sky130_fd_sc_hd__dfxtp_1
X_5472_ _5472_/A vssd1 vssd1 vccd1 vccd1 _5472_/X sky130_fd_sc_hd__buf_6
X_4423_ _4431_/B vssd1 vssd1 vccd1 vccd1 _4423_/Y sky130_fd_sc_hd__inv_2
X_7142_ _7344_/CLK _7142_/D vssd1 vssd1 vccd1 vccd1 _7142_/Q sky130_fd_sc_hd__dfxtp_1
X_4354_ _4354_/A vssd1 vssd1 vccd1 vccd1 _7503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7073_ _7073_/A vssd1 vssd1 vccd1 vccd1 _7846_/D sky130_fd_sc_hd__clkbuf_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6024_ _6024_/A vssd1 vssd1 vccd1 vccd1 _6024_/X sky130_fd_sc_hd__clkbuf_4
X_4285_ _4285_/A _4285_/B vssd1 vssd1 vccd1 vccd1 _4286_/C sky130_fd_sc_hd__or2_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6743__132 _6743__132/A vssd1 vssd1 vccd1 vccd1 _7699_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ _6923_/Y _6925_/X _7014_/A vssd1 vssd1 vccd1 vccd1 _7797_/D sky130_fd_sc_hd__a21oi_1
Xclkbuf_0__2985_ _6117_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2985_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_81_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6857_ _6857_/A vssd1 vssd1 vccd1 vccd1 _6857_/X sky130_fd_sc_hd__buf_1
XFILLER_80_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5808_ _5820_/A vssd1 vssd1 vccd1 vccd1 _5808_/X sky130_fd_sc_hd__buf_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7409_ _7409_/CLK _7409_/D vssd1 vssd1 vccd1 vccd1 _7409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_40 _4054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4070_ _4069_/X _7603_/Q _4070_/S vssd1 vssd1 vccd1 vccd1 _4071_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7760_ _7760_/CLK _7760_/D vssd1 vssd1 vccd1 vccd1 _7760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4972_ _4972_/A vssd1 vssd1 vccd1 vccd1 _7160_/D sky130_fd_sc_hd__clkbuf_1
X_6711_ _6711_/A _6711_/B _6711_/C _6711_/D vssd1 vssd1 vccd1 vccd1 _6711_/Y sky130_fd_sc_hd__nand4_1
X_7691_ _7691_/CLK _7691_/D vssd1 vssd1 vccd1 vccd1 _7691_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2770_ _5795_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2770_/X sky130_fd_sc_hd__clkbuf_16
X_3923_ _3923_/A vssd1 vssd1 vccd1 vccd1 _7662_/D sky130_fd_sc_hd__clkbuf_1
X_3854_ _3854_/A vssd1 vssd1 vccd1 vccd1 _7708_/D sky130_fd_sc_hd__clkbuf_1
X_6298__408 _6298__408/A vssd1 vssd1 vccd1 vccd1 _7461_/CLK sky130_fd_sc_hd__inv_2
X_6573_ _6573_/A vssd1 vssd1 vccd1 vccd1 _6621_/B sky130_fd_sc_hd__clkbuf_2
X_3785_ _7524_/Q vssd1 vssd1 vccd1 vccd1 _4194_/A sky130_fd_sc_hd__clkbuf_2
X_6378__454 _6378__454/A vssd1 vssd1 vccd1 vccd1 _7517_/CLK sky130_fd_sc_hd__inv_2
X_5524_ _5505_/X _5511_/X _5517_/X _5523_/X _4291_/A _5602_/S vssd1 vssd1 vccd1 vccd1
+ _5524_/X sky130_fd_sc_hd__mux4_2
XFILLER_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5455_ _5634_/B vssd1 vssd1 vccd1 vccd1 _5455_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4406_ _4405_/X _7482_/Q _4409_/S vssd1 vssd1 vccd1 vccd1 _4407_/A sky130_fd_sc_hd__mux2_1
X_7125_ _7331_/CLK _7125_/D vssd1 vssd1 vccd1 vccd1 _7125_/Q sky130_fd_sc_hd__dfxtp_1
X_5386_ _7405_/Q vssd1 vssd1 vccd1 vccd1 _5463_/A sky130_fd_sc_hd__inv_2
XFILLER_113_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4337_ _4173_/X _7510_/Q _4337_/S vssd1 vssd1 vccd1 vccd1 _4338_/A sky130_fd_sc_hd__mux2_1
X_7056_ _7056_/A vssd1 vssd1 vccd1 vccd1 _7841_/D sky130_fd_sc_hd__clkbuf_1
X_4268_ _6310_/A vssd1 vssd1 vccd1 vccd1 _6308_/B sky130_fd_sc_hd__clkbuf_2
X_6007_ _7459_/Q vssd1 vssd1 vccd1 vccd1 _6099_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_39_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4199_ _4155_/X _7553_/Q _4205_/S vssd1 vssd1 vccd1 vccd1 _4200_/A sky130_fd_sc_hd__mux2_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _7003_/A vssd1 vssd1 vccd1 vccd1 _6909_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5739__214 _5739__214/A vssd1 vssd1 vccd1 vccd1 _7231_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7861__235 vssd1 vssd1 vccd1 vccd1 partID[8] _7861__235/LO sky130_fd_sc_hd__conb_1
XFILLER_33_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3570_ _3944_/A vssd1 vssd1 vccd1 vccd1 _3570_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _5338_/A vssd1 vssd1 vccd1 vccd1 _5269_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5171_ _7192_/Q _5175_/B _5171_/C vssd1 vssd1 vccd1 vccd1 _5171_/X sky130_fd_sc_hd__and3_1
XFILLER_84_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4122_ _4122_/A vssd1 vssd1 vccd1 vccd1 _7583_/D sky130_fd_sc_hd__clkbuf_1
X_4053_ _4053_/A vssd1 vssd1 vccd1 vccd1 _7609_/D sky130_fd_sc_hd__clkbuf_1
Xinput3 caravel_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7812_ _7812_/CLK _7812_/D vssd1 vssd1 vccd1 vccd1 _7812_/Q sky130_fd_sc_hd__dfxtp_1
X_7743_ _7743_/CLK _7743_/D vssd1 vssd1 vccd1 vccd1 _7743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4955_ _4955_/A _4955_/B vssd1 vssd1 vccd1 vccd1 _4971_/S sky130_fd_sc_hd__or2_2
X_3906_ _3906_/A vssd1 vssd1 vccd1 vccd1 _7688_/D sky130_fd_sc_hd__clkbuf_1
X_7674_ _7680_/CLK _7674_/D vssd1 vssd1 vccd1 vccd1 _7674_/Q sky130_fd_sc_hd__dfxtp_1
X_4886_ _4886_/A vssd1 vssd1 vccd1 vccd1 _7244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6625_ _6615_/A _6615_/B _7844_/Q vssd1 vssd1 vccd1 vccd1 _6625_/X sky130_fd_sc_hd__a21bo_1
XFILLER_20_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3837_ _3836_/X _7714_/Q _3841_/S vssd1 vssd1 vccd1 vccd1 _3838_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6556_ _7686_/Q _7685_/Q vssd1 vssd1 vccd1 vccd1 _6725_/D sky130_fd_sc_hd__and2_1
X_3768_ _3768_/A vssd1 vssd1 vccd1 vccd1 _7728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5507_ _7295_/Q _7287_/Q _7263_/Q _7111_/Q _5481_/X _5506_/X vssd1 vssd1 vccd1 vccd1
+ _5507_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_0__3305_ _6795_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3305_/X sky130_fd_sc_hd__clkbuf_16
X_3699_ _4028_/A _3928_/B vssd1 vssd1 vccd1 vccd1 _3722_/S sky130_fd_sc_hd__or2_2
XFILLER_10_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5438_ _7205_/Q vssd1 vssd1 vccd1 vccd1 _5439_/A sky130_fd_sc_hd__clkinv_2
X_7108_ _7331_/CLK _7108_/D vssd1 vssd1 vccd1 vccd1 _7108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6400__469 _6400__469/A vssd1 vssd1 vccd1 vccd1 _7534_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4740_/A vssd1 vssd1 vccd1 vccd1 _7305_/D sky130_fd_sc_hd__clkbuf_1
X_4671_ _4671_/A vssd1 vssd1 vccd1 vccd1 _7356_/D sky130_fd_sc_hd__clkbuf_1
X_7390_ _7390_/CLK _7390_/D vssd1 vssd1 vccd1 vccd1 _7390_/Q sky130_fd_sc_hd__dfxtp_1
X_3622_ _3566_/X _7780_/Q _3622_/S vssd1 vssd1 vccd1 vccd1 _3623_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3122_ clkbuf_0__3122_/X vssd1 vssd1 vccd1 vccd1 _6425__489/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3553_ _7828_/Q vssd1 vssd1 vccd1 vccd1 _3932_/A sky130_fd_sc_hd__clkbuf_4
X_5223_ _7142_/Q _5215_/X _5216_/X _5222_/X vssd1 vssd1 vccd1 vccd1 _5223_/X sky130_fd_sc_hd__o22a_4
XFILLER_102_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5154_ _7118_/Q _5145_/X input14/X _5146_/X _5153_/X vssd1 vssd1 vccd1 vccd1 _5154_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4105_ _4105_/A vssd1 vssd1 vccd1 vccd1 _7588_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5085_ _5085_/A _5087_/B vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__and2_1
XFILLER_110_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4036_ _3938_/X _7615_/Q _4038_/S vssd1 vssd1 vccd1 vccd1 _4037_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5987_ _5978_/X _5981_/X _5986_/X _5964_/X vssd1 vssd1 vccd1 vccd1 _5987_/X sky130_fd_sc_hd__o211a_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__2768_ clkbuf_0__2768_/X vssd1 vssd1 vccd1 vccd1 _5788__254/A sky130_fd_sc_hd__clkbuf_4
X_7726_ _7726_/CLK _7726_/D vssd1 vssd1 vccd1 vccd1 _7726_/Q sky130_fd_sc_hd__dfxtp_1
X_4938_ _4953_/S vssd1 vssd1 vccd1 vccd1 _4947_/S sky130_fd_sc_hd__buf_2
XFILLER_33_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7657_ _7657_/CLK _7657_/D vssd1 vssd1 vccd1 vccd1 _7657_/Q sky130_fd_sc_hd__dfxtp_1
X_4869_ _7251_/Q _4399_/A _4875_/S vssd1 vssd1 vccd1 vccd1 _4870_/A sky130_fd_sc_hd__mux2_1
X_6608_ _6566_/X _6567_/Y _6588_/X _6601_/Y _6607_/X vssd1 vssd1 vccd1 vccd1 _6630_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_115_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7588_ _7588_/CLK _7588_/D vssd1 vssd1 vccd1 vccd1 _7588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5809__270 _5813__274/A vssd1 vssd1 vccd1 vccd1 _7287_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__2984_ clkbuf_0__2984_/X vssd1 vssd1 vccd1 vccd1 _6116__334/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput170 _5205_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[18] sky130_fd_sc_hd__buf_2
XFILLER_0_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput192 _5176_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[9] sky130_fd_sc_hd__buf_2
Xoutput181 _5229_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[28] sky130_fd_sc_hd__buf_2
XFILLER_87_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__3130_ clkbuf_0__3130_/X vssd1 vssd1 vccd1 vccd1 _6465__521/A sky130_fd_sc_hd__clkbuf_16
XFILLER_109_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6890_ _7850_/Q _6890_/B vssd1 vssd1 vccd1 vccd1 _6890_/X sky130_fd_sc_hd__xor2_1
XFILLER_46_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__2776_ clkbuf_0__2776_/X vssd1 vssd1 vccd1 vccd1 _6269_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4723_ _4722_/X _7311_/Q _4729_/S vssd1 vssd1 vccd1 vccd1 _4724_/A sky130_fd_sc_hd__mux2_1
X_7511_ _7511_/CLK _7511_/D vssd1 vssd1 vccd1 vccd1 _7511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7442_ _7442_/CLK _7442_/D vssd1 vssd1 vccd1 vccd1 _7442_/Q sky130_fd_sc_hd__dfxtp_1
X_4654_ _4399_/X _7363_/Q _4660_/S vssd1 vssd1 vccd1 vccd1 _4655_/A sky130_fd_sc_hd__mux2_1
X_4585_ _4585_/A vssd1 vssd1 vccd1 vccd1 _7402_/D sky130_fd_sc_hd__clkbuf_1
X_7373_ _7373_/CLK _7373_/D vssd1 vssd1 vccd1 vccd1 _7373_/Q sky130_fd_sc_hd__dfxtp_1
X_3605_ _3605_/A vssd1 vssd1 vccd1 vccd1 _7787_/D sky130_fd_sc_hd__clkbuf_1
Xinput50 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _5098_/A sky130_fd_sc_hd__buf_6
Xinput61 wbs_data_i[16] vssd1 vssd1 vccd1 vccd1 _5049_/A sky130_fd_sc_hd__buf_4
Xinput72 wbs_data_i[26] vssd1 vssd1 vccd1 vccd1 _5071_/A sky130_fd_sc_hd__buf_4
X_7874__201 vssd1 vssd1 vccd1 vccd1 _7874__201/HI core1Index[1] sky130_fd_sc_hd__conb_1
Xclkbuf_0__2452_ _5383_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2452_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3536_ _7466_/Q _7461_/Q vssd1 vssd1 vccd1 vccd1 _4448_/B sky130_fd_sc_hd__xnor2_2
Xclkbuf_1_1_0__3105_ clkbuf_0__3105_/X vssd1 vssd1 vccd1 vccd1 _6341__424/A sky130_fd_sc_hd__clkbuf_4
Xinput83 wbs_data_i[7] vssd1 vssd1 vccd1 vccd1 _7030_/A sky130_fd_sc_hd__buf_8
X_6324_ _6324_/A _6396_/A vssd1 vssd1 vccd1 vccd1 _7475_/D sky130_fd_sc_hd__nor2_1
X_6255_ _7793_/Q vssd1 vssd1 vccd1 vccd1 _6900_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5206_ _5217_/A vssd1 vssd1 vccd1 vccd1 _5206_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6186_ _7808_/Q _6188_/B _7809_/Q vssd1 vssd1 vccd1 vccd1 _6869_/B sky130_fd_sc_hd__a21o_1
X_5137_ _5177_/A vssd1 vssd1 vccd1 vccd1 _5138_/D sky130_fd_sc_hd__buf_6
X_5068_ _5068_/A vssd1 vssd1 vccd1 vccd1 _5077_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4019_ _4019_/A vssd1 vssd1 vccd1 vccd1 _7623_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7709_ _7709_/CLK _7709_/D vssd1 vssd1 vccd1 vccd1 _7709_/Q sky130_fd_sc_hd__dfxtp_1
X_6792__172 _6792__172/A vssd1 vssd1 vccd1 vccd1 _7739_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6372__449 _6372__449/A vssd1 vssd1 vccd1 vccd1 _7512_/CLK sky130_fd_sc_hd__inv_2
X_4370_ _4370_/A vssd1 vssd1 vccd1 vccd1 _7496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _7623_/Q _7615_/Q _7607_/Q _7599_/Q _5933_/X _5998_/X vssd1 vssd1 vccd1 vccd1
+ _6040_/X sky130_fd_sc_hd__mux4_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6942_ _7802_/Q _6952_/B vssd1 vssd1 vccd1 vccd1 _6942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7687_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6873_ _7847_/Q _6873_/B vssd1 vssd1 vccd1 vccd1 _6873_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5686_ _5493_/A _5090_/A _5692_/S vssd1 vssd1 vccd1 vccd1 _5687_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4706_ _4706_/A _4847_/B vssd1 vssd1 vccd1 vccd1 _4729_/S sky130_fd_sc_hd__or2_4
X_4637_ _4637_/A vssd1 vssd1 vccd1 vccd1 _7379_/D sky130_fd_sc_hd__clkbuf_1
X_7425_ _7425_/CLK _7425_/D vssd1 vssd1 vccd1 vccd1 _7425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4568_ _4253_/X _7412_/Q _4570_/S vssd1 vssd1 vccd1 vccd1 _4569_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7356_ _7356_/CLK _7356_/D vssd1 vssd1 vccd1 vccd1 _7356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3519_ _7224_/Q _7225_/Q _7215_/Q _7214_/Q vssd1 vssd1 vccd1 vccd1 _3520_/B sky130_fd_sc_hd__or4b_1
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7287_ _7287_/CLK _7287_/D vssd1 vssd1 vccd1 vccd1 _7287_/Q sky130_fd_sc_hd__dfxtp_1
X_4499_ _4411_/X _7443_/Q _4503_/S vssd1 vssd1 vccd1 vccd1 _4500_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6238_ _6238_/A _6238_/B _6238_/C _6238_/D vssd1 vssd1 vccd1 vccd1 _6253_/B sky130_fd_sc_hd__and4_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3304_ clkbuf_0__3304_/X vssd1 vssd1 vccd1 vccd1 _6794__174/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6799__178 _6800__179/A vssd1 vssd1 vccd1 vccd1 _7745_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3870_ _3784_/X _7704_/Q _3878_/S vssd1 vssd1 vccd1 vccd1 _3871_/A sky130_fd_sc_hd__mux2_1
X_5788__254 _5788__254/A vssd1 vssd1 vccd1 vccd1 _7271_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5540_ _7179_/Q _7360_/Q _7716_/Q _7256_/Q _5520_/X _5521_/X vssd1 vssd1 vccd1 vccd1
+ _5540_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5471_ _7519_/Q vssd1 vssd1 vccd1 vccd1 _5472_/A sky130_fd_sc_hd__clkbuf_4
X_4422_ _7467_/Q _7476_/Q _3927_/B _4421_/X vssd1 vssd1 vccd1 vccd1 _7467_/D sky130_fd_sc_hd__o211a_1
X_7210_ _7826_/CLK _7210_/D vssd1 vssd1 vccd1 vccd1 _7210_/Q sky130_fd_sc_hd__dfxtp_1
X_7141_ _7344_/CLK _7141_/D vssd1 vssd1 vccd1 vccd1 _7141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4353_ _4170_/X _7503_/Q _4355_/S vssd1 vssd1 vccd1 vccd1 _4354_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7072_ _7070_/X _7072_/B vssd1 vssd1 vccd1 vccd1 _7073_/A sky130_fd_sc_hd__and2b_1
X_4284_ _4284_/A _4284_/B vssd1 vssd1 vccd1 vccd1 _7524_/D sky130_fd_sc_hd__nor2_1
XFILLER_100_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6023_ _7724_/Q _7708_/Q _7427_/Q _7489_/Q _5939_/X _5974_/X vssd1 vssd1 vccd1 vccd1
+ _6023_/X sky130_fd_sc_hd__mux4_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6925_ _6924_/X _6907_/X _6880_/B vssd1 vssd1 vccd1 vccd1 _6925_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__2984_ _6111_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2984_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_62_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3999_ _3938_/X _7631_/Q _4001_/S vssd1 vssd1 vccd1 vccd1 _4000_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5669_ _7839_/Q _5679_/A _7407_/Q _5672_/D vssd1 vssd1 vccd1 vccd1 _5669_/X sky130_fd_sc_hd__and4_1
X_7408_ _7408_/CLK _7408_/D vssd1 vssd1 vccd1 vccd1 _7408_/Q sky130_fd_sc_hd__dfxtp_1
X_7339_ _7339_/CLK _7339_/D vssd1 vssd1 vccd1 vccd1 _7339_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_30 _5087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_41 _4213_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5380__208 _5381__209/A vssd1 vssd1 vccd1 vccd1 _7180_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4971_ _4239_/X _7160_/Q _4971_/S vssd1 vssd1 vccd1 vccd1 _4972_/A sky130_fd_sc_hd__mux2_1
X_6710_ _6679_/A _6684_/X _7683_/Q vssd1 vssd1 vccd1 vccd1 _6710_/X sky130_fd_sc_hd__a21bo_1
XFILLER_17_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7690_ _7690_/CLK _7690_/D vssd1 vssd1 vccd1 vccd1 _7690_/Q sky130_fd_sc_hd__dfxtp_1
X_3922_ _3836_/X _7662_/Q _3924_/S vssd1 vssd1 vccd1 vccd1 _3923_/A sky130_fd_sc_hd__mux2_1
X_6641_ _6641_/A vssd1 vssd1 vccd1 vccd1 _7660_/D sky130_fd_sc_hd__clkbuf_1
X_3853_ _3712_/X _7708_/Q _3853_/S vssd1 vssd1 vccd1 vccd1 _3854_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6572_ _6613_/A _6613_/B _6621_/D vssd1 vssd1 vccd1 vccd1 _6696_/B sky130_fd_sc_hd__nand3_1
X_3784_ _4393_/A vssd1 vssd1 vccd1 vccd1 _3784_/X sky130_fd_sc_hd__buf_2
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5523_ _5519_/X _5522_/X _5578_/S vssd1 vssd1 vccd1 vccd1 _5523_/X sky130_fd_sc_hd__mux2_1
X_5454_ _7040_/A vssd1 vssd1 vccd1 vccd1 _5634_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4405_ _4405_/A vssd1 vssd1 vccd1 vccd1 _4405_/X sky130_fd_sc_hd__buf_2
X_7124_ _7331_/CLK _7124_/D vssd1 vssd1 vccd1 vccd1 _7124_/Q sky130_fd_sc_hd__dfxtp_1
X_5803__265 _5805__267/A vssd1 vssd1 vccd1 vccd1 _7282_/CLK sky130_fd_sc_hd__inv_2
X_4336_ _4336_/A vssd1 vssd1 vccd1 vccd1 _7511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7055_ _7048_/X _7055_/B vssd1 vssd1 vccd1 vccd1 _7056_/A sky130_fd_sc_hd__and2b_1
X_4267_ _4267_/A vssd1 vssd1 vccd1 vccd1 _7531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6006_ _7787_/Q _7779_/Q _7771_/Q _7763_/Q _5979_/X _5980_/X vssd1 vssd1 vccd1 vccd1
+ _6006_/X sky130_fd_sc_hd__mux4_1
XFILLER_86_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_31_wb_clk_i _7474_/CLK vssd1 vssd1 vccd1 vccd1 _7802_/CLK sky130_fd_sc_hd__clkbuf_16
X_4198_ _4198_/A vssd1 vssd1 vccd1 vccd1 _7554_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__2451_ clkbuf_0__2451_/X vssd1 vssd1 vccd1 vccd1 _5758_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6908_ _6916_/B _6907_/X _6904_/C _6916_/A vssd1 vssd1 vccd1 vccd1 _6908_/X sky130_fd_sc_hd__a31o_1
XFILLER_24_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6839_ _6845_/A vssd1 vssd1 vccd1 vccd1 _6839_/X sky130_fd_sc_hd__buf_1
XFILLER_50_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5170_ _7124_/Q _5159_/X input32/X _5163_/X _5169_/X vssd1 vssd1 vccd1 vccd1 _5170_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4121_ _3824_/X _7583_/Q _4123_/S vssd1 vssd1 vccd1 vccd1 _4122_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4052_ _4051_/X _7609_/Q _4061_/S vssd1 vssd1 vccd1 vccd1 _4053_/A sky130_fd_sc_hd__mux2_1
Xinput4 caravel_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7811_ _7812_/CLK _7811_/D vssd1 vssd1 vccd1 vccd1 _7811_/Q sky130_fd_sc_hd__dfxtp_1
X_7742_ _7742_/CLK _7742_/D vssd1 vssd1 vccd1 vccd1 _7742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4954_ _4954_/A vssd1 vssd1 vccd1 vccd1 _7168_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3905_ _3840_/X _7688_/Q _3905_/S vssd1 vssd1 vccd1 vccd1 _3906_/A sky130_fd_sc_hd__mux2_1
X_7673_ _7680_/CLK _7673_/D vssd1 vssd1 vccd1 vccd1 _7673_/Q sky130_fd_sc_hd__dfxtp_1
X_4885_ _4803_/X _7244_/Q _4893_/S vssd1 vssd1 vccd1 vccd1 _4886_/A sky130_fd_sc_hd__mux2_1
X_6624_ _6699_/B _6699_/C _6249_/A vssd1 vssd1 vccd1 vccd1 _6624_/Y sky130_fd_sc_hd__a21oi_1
X_3836_ _4414_/A vssd1 vssd1 vccd1 vccd1 _3836_/X sky130_fd_sc_hd__buf_2
X_3767_ _3698_/X _7728_/Q _3775_/S vssd1 vssd1 vccd1 vccd1 _3768_/A sky130_fd_sc_hd__mux2_1
X_5506_ _5521_/A vssd1 vssd1 vccd1 vccd1 _5506_/X sky130_fd_sc_hd__buf_4
X_3698_ _3926_/A vssd1 vssd1 vccd1 vccd1 _3698_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3304_ _6789_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3304_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_10_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5437_ _5437_/A vssd1 vssd1 vccd1 vccd1 _6396_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5299_ _5307_/A vssd1 vssd1 vccd1 vccd1 _5299_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7107_ _7107_/A vssd1 vssd1 vccd1 vccd1 _7855_/D sky130_fd_sc_hd__clkbuf_1
X_4319_ _4319_/A vssd1 vssd1 vccd1 vccd1 _7518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6467__523 _6468__524/A vssd1 vssd1 vccd1 vccd1 _7588_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6494__64 _6494__64/A vssd1 vssd1 vccd1 vccd1 _7609_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6756__143 _6757__144/A vssd1 vssd1 vccd1 vccd1 _7710_/CLK sky130_fd_sc_hd__inv_2
X_5257__185 _5259__187/A vssd1 vssd1 vccd1 vccd1 _7114_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7891__218 vssd1 vssd1 vccd1 vccd1 _7891__218/HI manufacturerID[10] sky130_fd_sc_hd__conb_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4670_ _3649_/X _7356_/Q _4678_/S vssd1 vssd1 vccd1 vccd1 _4671_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3621_ _3621_/A vssd1 vssd1 vccd1 vccd1 _7781_/D sky130_fd_sc_hd__clkbuf_1
X_3552_ _3552_/A vssd1 vssd1 vccd1 vccd1 _7837_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3121_ clkbuf_0__3121_/X vssd1 vssd1 vccd1 vccd1 _6432_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5222_ _5217_/X _5222_/B vssd1 vssd1 vccd1 vccd1 _5222_/X sky130_fd_sc_hd__and2b_1
X_6549__108 _6550__109/A vssd1 vssd1 vccd1 vccd1 _7653_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5153_ _7185_/Q _5161_/B _5215_/A vssd1 vssd1 vccd1 vccd1 _5153_/X sky130_fd_sc_hd__and3_1
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4104_ _4066_/X _7588_/Q _4106_/S vssd1 vssd1 vccd1 vccd1 _4105_/A sky130_fd_sc_hd__mux2_1
X_5084_ _5084_/A vssd1 vssd1 vccd1 vccd1 _5084_/X sky130_fd_sc_hd__clkbuf_1
X_5915__311 _5916__312/A vssd1 vssd1 vccd1 vccd1 _7352_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4035_ _4035_/A vssd1 vssd1 vccd1 vccd1 _7616_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5986_ _6079_/A _5986_/B vssd1 vssd1 vccd1 vccd1 _5986_/X sky130_fd_sc_hd__or2_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__2767_ clkbuf_0__2767_/X vssd1 vssd1 vccd1 vccd1 _5779__246/A sky130_fd_sc_hd__clkbuf_4
X_7725_ _7725_/CLK _7725_/D vssd1 vssd1 vccd1 vccd1 _7725_/Q sky130_fd_sc_hd__dfxtp_1
X_4937_ _4937_/A _4937_/B vssd1 vssd1 vccd1 vccd1 _4953_/S sky130_fd_sc_hd__nand2_2
X_7656_ _7656_/CLK _7656_/D vssd1 vssd1 vccd1 vccd1 _7656_/Q sky130_fd_sc_hd__dfxtp_1
X_4868_ _4868_/A vssd1 vssd1 vccd1 vccd1 _7252_/D sky130_fd_sc_hd__clkbuf_1
X_6607_ _5584_/X _6686_/B _6604_/X _6605_/Y _6606_/Y vssd1 vssd1 vccd1 vccd1 _6607_/X
+ sky130_fd_sc_hd__o2111a_1
X_3819_ _7473_/Q vssd1 vssd1 vccd1 vccd1 _4402_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7587_ _7587_/CLK _7587_/D vssd1 vssd1 vccd1 vccd1 _7587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4799_ _4725_/X _7278_/Q _4801_/S vssd1 vssd1 vccd1 vccd1 _4800_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2983_ clkbuf_0__2983_/X vssd1 vssd1 vccd1 vccd1 _6108__327/A sky130_fd_sc_hd__clkbuf_4
X_6538_ _6538_/A vssd1 vssd1 vccd1 vccd1 _6538_/X sky130_fd_sc_hd__buf_1
XFILLER_21_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6469_ _6469_/A vssd1 vssd1 vccd1 vccd1 _6469_/X sky130_fd_sc_hd__buf_1
Xoutput160 _5238_/X vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
Xoutput171 _5208_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[19] sky130_fd_sc_hd__buf_2
Xoutput182 _5231_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[29] sky130_fd_sc_hd__buf_2
XFILLER_102_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5782__249 _5782__249/A vssd1 vssd1 vccd1 vccd1 _7266_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6730__124 _6730__124/A vssd1 vssd1 vccd1 vccd1 _7690_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5840_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5840_/X sky130_fd_sc_hd__buf_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5771_ _5771_/A vssd1 vssd1 vccd1 vccd1 _5771_/X sky130_fd_sc_hd__buf_1
XFILLER_21_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4722_ _7470_/Q vssd1 vssd1 vccd1 vccd1 _4722_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7510_ _7510_/CLK _7510_/D vssd1 vssd1 vccd1 vccd1 _7510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7441_ _7441_/CLK _7441_/D vssd1 vssd1 vccd1 vccd1 _7441_/Q sky130_fd_sc_hd__dfxtp_1
Xinput40 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 _5109_/A sky130_fd_sc_hd__buf_4
X_4653_ _4653_/A vssd1 vssd1 vccd1 vccd1 _7364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4584_ _7402_/Q _3935_/A _4588_/S vssd1 vssd1 vccd1 vccd1 _4585_/A sky130_fd_sc_hd__mux2_1
X_7372_ _7372_/CLK _7372_/D vssd1 vssd1 vccd1 vccd1 _7372_/Q sky130_fd_sc_hd__dfxtp_1
X_3604_ _3570_/X _7787_/Q _3608_/S vssd1 vssd1 vccd1 vccd1 _3605_/A sky130_fd_sc_hd__mux2_1
Xinput51 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 _5101_/A sky130_fd_sc_hd__buf_4
Xinput62 wbs_data_i[17] vssd1 vssd1 vccd1 vccd1 _5051_/A sky130_fd_sc_hd__buf_4
Xinput73 wbs_data_i[27] vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__buf_4
Xclkbuf_0__2451_ _5382_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2451_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1_0__3104_ clkbuf_0__3104_/X vssd1 vssd1 vccd1 vccd1 _6333__417/A sky130_fd_sc_hd__clkbuf_4
X_3535_ _3535_/A vssd1 vssd1 vccd1 vccd1 _5932_/A sky130_fd_sc_hd__clkbuf_2
Xinput84 wbs_data_i[8] vssd1 vssd1 vccd1 vccd1 _5031_/A sky130_fd_sc_hd__buf_6
X_6323_ _7821_/Q vssd1 vssd1 vccd1 vccd1 _6324_/A sky130_fd_sc_hd__inv_2
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6254_ _7794_/Q vssd1 vssd1 vccd1 vccd1 _6859_/A sky130_fd_sc_hd__inv_2
X_5205_ _7135_/Q _5199_/X _5201_/X _5204_/X vssd1 vssd1 vccd1 vccd1 _5205_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6185_ _6251_/B vssd1 vssd1 vccd1 vccd1 _6869_/A sky130_fd_sc_hd__clkbuf_2
X_5136_ _5136_/A vssd1 vssd1 vccd1 vccd1 _5136_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5067_ _5067_/A vssd1 vssd1 vccd1 vccd1 _5067_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4018_ _3938_/X _7623_/Q _4020_/S vssd1 vssd1 vccd1 vccd1 _4019_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5969_ _6737_/S vssd1 vssd1 vccd1 vccd1 _6723_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7708_ _7708_/CLK _7708_/D vssd1 vssd1 vccd1 vccd1 _7708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7639_ _7639_/CLK _7639_/D vssd1 vssd1 vccd1 vccd1 _7639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6527__90 _6529__92/A vssd1 vssd1 vccd1 vccd1 _7635_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7897__224 vssd1 vssd1 vccd1 vccd1 _7897__224/HI partID[12] sky130_fd_sc_hd__conb_1
XFILLER_117_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6941_ _6938_/Y _6940_/X _6935_/X vssd1 vssd1 vccd1 vccd1 _7801_/D sky130_fd_sc_hd__a21oi_1
XFILLER_47_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6872_ _6872_/A _6872_/B vssd1 vssd1 vccd1 vccd1 _6893_/A sky130_fd_sc_hd__xnor2_1
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5685_ _5685_/A vssd1 vssd1 vccd1 vccd1 _7204_/D sky130_fd_sc_hd__clkbuf_1
X_4705_ _7475_/Q vssd1 vssd1 vccd1 vccd1 _4705_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4636_ _3657_/X _7379_/Q _4642_/S vssd1 vssd1 vccd1 vccd1 _4637_/A sky130_fd_sc_hd__mux2_1
X_7424_ _7424_/CLK _7424_/D vssd1 vssd1 vccd1 vccd1 _7424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7355_ _7355_/CLK _7355_/D vssd1 vssd1 vccd1 vccd1 _7355_/Q sky130_fd_sc_hd__dfxtp_1
X_4567_ _4567_/A vssd1 vssd1 vccd1 vccd1 _7413_/D sky130_fd_sc_hd__clkbuf_1
X_3518_ _7216_/Q _7217_/Q _7212_/Q _7213_/Q vssd1 vssd1 vccd1 vccd1 _5399_/C sky130_fd_sc_hd__or4_1
XFILLER_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4498_ _4498_/A vssd1 vssd1 vccd1 vccd1 _7444_/D sky130_fd_sc_hd__clkbuf_1
X_7286_ _7286_/CLK _7286_/D vssd1 vssd1 vccd1 vccd1 _7286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6237_ _6872_/A _6873_/B _6235_/Y _6236_/X vssd1 vssd1 vccd1 vccd1 _6238_/D sky130_fd_sc_hd__o22a_1
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _5119_/A vssd1 vssd1 vccd1 vccd1 _5119_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6099_ _6099_/A _6099_/B vssd1 vssd1 vccd1 vccd1 _6099_/X sky130_fd_sc_hd__or2_1
Xclkbuf_1_0_0__3303_ clkbuf_0__3303_/X vssd1 vssd1 vccd1 vccd1 _6787__168/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3234_ clkbuf_0__3234_/X vssd1 vssd1 vccd1 vccd1 _6651__121/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5470_ _5590_/A _5465_/X _5469_/X vssd1 vssd1 vccd1 vccd1 _5470_/X sky130_fd_sc_hd__a21o_1
X_5829__285 _5830__286/A vssd1 vssd1 vccd1 vccd1 _7302_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4421_ _6328_/B vssd1 vssd1 vccd1 vccd1 _4421_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7140_ _7344_/CLK _7140_/D vssd1 vssd1 vccd1 vccd1 _7140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4352_ _4352_/A vssd1 vssd1 vccd1 vccd1 _7504_/D sky130_fd_sc_hd__clkbuf_1
X_7071_ _5033_/A _7846_/Q _7074_/S vssd1 vssd1 vccd1 vccd1 _7072_/B sky130_fd_sc_hd__mux2_1
X_6521__85 _6525__89/A vssd1 vssd1 vccd1 vccd1 _7630_/CLK sky130_fd_sc_hd__inv_2
X_4283_ _4150_/B _4286_/B _4280_/A vssd1 vssd1 vccd1 vccd1 _4284_/B sky130_fd_sc_hd__a21o_1
XFILLER_98_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6022_ _7574_/Q _7384_/Q _7732_/Q _7630_/Q _6002_/X _4450_/A vssd1 vssd1 vccd1 vccd1
+ _6022_/X sky130_fd_sc_hd__mux4_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6461__518 _6462__519/A vssd1 vssd1 vccd1 vccd1 _7583_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6924_ _6943_/A vssd1 vssd1 vccd1 vccd1 _6924_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__2983_ _6105_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2983_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_82_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3998_ _3998_/A vssd1 vssd1 vccd1 vccd1 _7632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__2449_ clkbuf_0__2449_/X vssd1 vssd1 vccd1 vccd1 _5375__204/A sky130_fd_sc_hd__clkbuf_4
X_5668_ _5668_/A vssd1 vssd1 vccd1 vccd1 _7199_/D sky130_fd_sc_hd__clkbuf_1
X_7407_ _7407_/CLK _7407_/D vssd1 vssd1 vccd1 vccd1 _7407_/Q sky130_fd_sc_hd__dfxtp_1
X_6750__138 _6751__139/A vssd1 vssd1 vccd1 vccd1 _7705_/CLK sky130_fd_sc_hd__inv_2
X_4619_ _4619_/A vssd1 vssd1 vccd1 vccd1 _7387_/D sky130_fd_sc_hd__clkbuf_1
X_5599_ _7585_/Q _7569_/Q _7553_/Q _7545_/Q _5427_/A _5472_/X vssd1 vssd1 vccd1 vccd1
+ _5599_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7338_ _7339_/CLK _7338_/D vssd1 vssd1 vccd1 vccd1 _7338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7269_ _7269_/CLK _7269_/D vssd1 vssd1 vccd1 vccd1 _7269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_31 _5094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_20 _5156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_42 _4803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3148_ clkbuf_0__3148_/X vssd1 vssd1 vccd1 vccd1 _6555__113/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4970_ _4970_/A vssd1 vssd1 vccd1 vccd1 _7161_/D sky130_fd_sc_hd__clkbuf_1
X_3921_ _3921_/A vssd1 vssd1 vccd1 vccd1 _7663_/D sky130_fd_sc_hd__clkbuf_1
X_6640_ _6723_/A _6640_/B _6640_/C vssd1 vssd1 vccd1 vccd1 _6641_/A sky130_fd_sc_hd__and3_1
X_3852_ _3852_/A vssd1 vssd1 vccd1 vccd1 _7709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6571_ _7678_/Q _6602_/A vssd1 vssd1 vccd1 vccd1 _6621_/D sky130_fd_sc_hd__and2_1
X_3783_ _7475_/Q vssd1 vssd1 vccd1 vccd1 _4393_/A sky130_fd_sc_hd__buf_2
X_5522_ _7512_/Q _7504_/Q _7443_/Q _7435_/Q _5520_/X _5521_/X vssd1 vssd1 vccd1 vccd1
+ _5522_/X sky130_fd_sc_hd__mux4_2
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5453_ _5453_/A vssd1 vssd1 vccd1 vccd1 _5453_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5250__180 _5252__182/A vssd1 vssd1 vccd1 vccd1 _7109_/CLK sky130_fd_sc_hd__inv_2
X_4404_ _4404_/A vssd1 vssd1 vccd1 vccd1 _7483_/D sky130_fd_sc_hd__clkbuf_1
X_7123_ _7372_/CLK _7123_/D vssd1 vssd1 vccd1 vccd1 _7123_/Q sky130_fd_sc_hd__dfxtp_1
X_4335_ _4170_/X _7511_/Q _4337_/S vssd1 vssd1 vccd1 vccd1 _4336_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7054_ _5044_/A _5661_/X _7067_/S vssd1 vssd1 vccd1 vccd1 _7055_/B sky130_fd_sc_hd__mux2_1
X_4266_ _4265_/X _7531_/Q _4266_/S vssd1 vssd1 vccd1 vccd1 _4267_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6005_ _6016_/A vssd1 vssd1 vccd1 vccd1 _6005_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2450_ clkbuf_0__2450_/X vssd1 vssd1 vccd1 vccd1 _5381__209/A sky130_fd_sc_hd__clkbuf_4
X_4197_ _4149_/X _7554_/Q _4205_/S vssd1 vssd1 vccd1 vccd1 _4198_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2998_ clkbuf_0__2998_/X vssd1 vssd1 vccd1 vccd1 _6177__378/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6168__370 _6169__371/A vssd1 vssd1 vccd1 vccd1 _7422_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ _6939_/A vssd1 vssd1 vccd1 vccd1 _6907_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6542__103 _6543__104/A vssd1 vssd1 vccd1 vccd1 _7648_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4120_ _4120_/A vssd1 vssd1 vccd1 vccd1 _7584_/D sky130_fd_sc_hd__clkbuf_1
X_4051_ _7828_/Q vssd1 vssd1 vccd1 vccd1 _4051_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 caravel_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7810_ _7812_/CLK _7810_/D vssd1 vssd1 vccd1 vccd1 _7810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7741_ _7741_/CLK _7741_/D vssd1 vssd1 vccd1 vccd1 _7741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4953_ _4239_/X _7168_/Q _4953_/S vssd1 vssd1 vccd1 vccd1 _4954_/A sky130_fd_sc_hd__mux2_1
X_7672_ _7845_/CLK _7672_/D vssd1 vssd1 vccd1 vccd1 _7672_/Q sky130_fd_sc_hd__dfxtp_1
X_3904_ _3904_/A vssd1 vssd1 vccd1 vccd1 _7689_/D sky130_fd_sc_hd__clkbuf_1
X_6623_ _7845_/Q _6699_/B _6699_/C vssd1 vssd1 vccd1 vccd1 _6623_/X sky130_fd_sc_hd__and3_1
X_4884_ _4899_/S vssd1 vssd1 vccd1 vccd1 _4893_/S sky130_fd_sc_hd__buf_2
X_3835_ _7469_/Q vssd1 vssd1 vccd1 vccd1 _4414_/A sky130_fd_sc_hd__buf_2
XFILLER_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3766_ _3781_/S vssd1 vssd1 vccd1 vccd1 _3775_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5505_ _5503_/X _5504_/X _5569_/S vssd1 vssd1 vccd1 vccd1 _5505_/X sky130_fd_sc_hd__mux2_1
X_3697_ _3697_/A vssd1 vssd1 vccd1 vccd1 _7753_/D sky130_fd_sc_hd__clkbuf_1
X_5436_ _5436_/A _5446_/B vssd1 vssd1 vccd1 vccd1 _5437_/A sky130_fd_sc_hd__or2_1
Xclkbuf_0__3303_ _6783_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3303_/X sky130_fd_sc_hd__clkbuf_16
X_6391__464 _6391__464/A vssd1 vssd1 vccd1 vccd1 _7527_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3234_ _6649_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3234_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_113_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5298_ _5295_/X _7336_/Q _5291_/X _5292_/X _7136_/Q vssd1 vssd1 vccd1 vccd1 _7136_/D
+ sky130_fd_sc_hd__o32a_1
X_7106_ _7106_/A _7106_/B _7106_/C vssd1 vssd1 vccd1 vccd1 _7107_/A sky130_fd_sc_hd__or3_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4318_ _4312_/B _4318_/B _6394_/C vssd1 vssd1 vccd1 vccd1 _4319_/A sky130_fd_sc_hd__and3b_1
X_4249_ _4249_/A vssd1 vssd1 vccd1 vccd1 _7537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5851__304 _5851__304/A vssd1 vssd1 vccd1 vccd1 _7321_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3620_ _3562_/X _7781_/Q _3622_/S vssd1 vssd1 vccd1 vccd1 _3621_/A sky130_fd_sc_hd__mux2_1
X_3551_ _3505_/X _7837_/Q _3567_/S vssd1 vssd1 vccd1 vccd1 _3552_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3120_ clkbuf_0__3120_/X vssd1 vssd1 vccd1 vccd1 _6417__483/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6270_ _6282_/A vssd1 vssd1 vccd1 vccd1 _6270_/X sky130_fd_sc_hd__buf_1
X_5221_ _7141_/Q _5215_/X _5216_/X _5220_/X vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__o22a_4
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5152_ _7117_/Q _5145_/X input3/X _5146_/X _5151_/X vssd1 vssd1 vccd1 vccd1 _5152_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4103_ _4103_/A vssd1 vssd1 vccd1 vccd1 _7589_/D sky130_fd_sc_hd__clkbuf_1
X_5083_ _5083_/A _5087_/B vssd1 vssd1 vccd1 vccd1 _5084_/A sky130_fd_sc_hd__and2_1
XFILLER_84_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4034_ _3935_/X _7616_/Q _4038_/S vssd1 vssd1 vccd1 vccd1 _4035_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5985_ _7390_/Q _7374_/Q _7644_/Q _7636_/Q _5983_/X _5984_/X vssd1 vssd1 vccd1 vccd1
+ _5986_/B sky130_fd_sc_hd__mux4_1
X_7724_ _7724_/CLK _7724_/D vssd1 vssd1 vccd1 vccd1 _7724_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4936_ _4936_/A vssd1 vssd1 vccd1 vccd1 _7176_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7655_ _7655_/CLK _7655_/D vssd1 vssd1 vccd1 vccd1 _7655_/Q sky130_fd_sc_hd__dfxtp_1
X_4867_ _7252_/Q _4393_/A _4875_/S vssd1 vssd1 vccd1 vccd1 _4868_/A sky130_fd_sc_hd__mux2_1
X_6606_ _5565_/X _6606_/B _6606_/C vssd1 vssd1 vccd1 vccd1 _6606_/Y sky130_fd_sc_hd__nand3b_1
X_3818_ _3818_/A vssd1 vssd1 vccd1 vccd1 _7719_/D sky130_fd_sc_hd__clkbuf_1
X_7586_ _7586_/CLK _7586_/D vssd1 vssd1 vccd1 vccd1 _7586_/Q sky130_fd_sc_hd__dfxtp_1
X_4798_ _4798_/A vssd1 vssd1 vccd1 vccd1 _7279_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3749_ _3749_/A vssd1 vssd1 vccd1 vccd1 _7736_/D sky130_fd_sc_hd__clkbuf_1
Xoutput150 _5028_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[6] sky130_fd_sc_hd__buf_2
Xoutput161 _5152_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[0] sky130_fd_sc_hd__buf_2
X_5419_ _7520_/Q vssd1 vssd1 vccd1 vccd1 _5590_/A sky130_fd_sc_hd__buf_2
XFILLER_114_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput172 _5154_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[1] sky130_fd_sc_hd__buf_2
Xoutput183 _5156_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[2] sky130_fd_sc_hd__buf_2
XFILLER_99_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3148_ _6551_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3148_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_48_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5816__276 _5818__278/A vssd1 vssd1 vccd1 vccd1 _7293_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _4721_/A vssd1 vssd1 vccd1 vccd1 _7312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6555__113 _6555__113/A vssd1 vssd1 vccd1 vccd1 _7658_/CLK sky130_fd_sc_hd__inv_2
X_7440_ _7440_/CLK _7440_/D vssd1 vssd1 vccd1 vccd1 _7440_/Q sky130_fd_sc_hd__dfxtp_1
X_4652_ _4393_/X _7364_/Q _4660_/S vssd1 vssd1 vccd1 vccd1 _4653_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput30 caravel_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_2
X_3603_ _3603_/A vssd1 vssd1 vccd1 vccd1 _7788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4583_ _4583_/A vssd1 vssd1 vccd1 vccd1 _7403_/D sky130_fd_sc_hd__clkbuf_1
X_7371_ _7372_/CLK _7371_/D vssd1 vssd1 vccd1 vccd1 _7371_/Q sky130_fd_sc_hd__dfxtp_1
Xinput52 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 _5103_/A sky130_fd_sc_hd__buf_4
Xinput41 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 _5112_/A sky130_fd_sc_hd__buf_4
Xinput63 wbs_data_i[18] vssd1 vssd1 vccd1 vccd1 _5053_/A sky130_fd_sc_hd__buf_4
Xclkbuf_0__2450_ _5376_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2450_/X sky130_fd_sc_hd__clkbuf_16
X_3534_ _7460_/Q vssd1 vssd1 vccd1 vccd1 _3535_/A sky130_fd_sc_hd__inv_2
Xinput85 wbs_data_i[9] vssd1 vssd1 vccd1 vccd1 _5033_/A sky130_fd_sc_hd__buf_6
Xinput74 wbs_data_i[28] vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__buf_4
X_6322_ _6322_/A vssd1 vssd1 vccd1 vccd1 _7474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6253_ _6253_/A _6253_/B _6253_/C _6993_/A vssd1 vssd1 vccd1 vccd1 _6260_/A sky130_fd_sc_hd__and4_1
XFILLER_115_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5204_ _5204_/A vssd1 vssd1 vccd1 vccd1 _5204_/X sky130_fd_sc_hd__buf_2
XFILLER_69_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6184_ _7809_/Q _7808_/Q _6188_/B vssd1 vssd1 vccd1 vccd1 _6251_/B sky130_fd_sc_hd__nand3_1
X_5135_ _7341_/Q _5142_/B vssd1 vssd1 vccd1 vccd1 _5136_/A sky130_fd_sc_hd__and2_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5066_ _5066_/A _5066_/B vssd1 vssd1 vccd1 vccd1 _5067_/A sky130_fd_sc_hd__or2_1
X_4017_ _4017_/A vssd1 vssd1 vccd1 vccd1 _7624_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6803__5 _6803__5/A vssd1 vssd1 vccd1 vccd1 _7747_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5968_ _5015_/A _3588_/X _5269_/A vssd1 vssd1 vccd1 vccd1 _6737_/S sky130_fd_sc_hd__a21oi_4
X_7707_ _7707_/CLK _7707_/D vssd1 vssd1 vccd1 vccd1 _7707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4919_ _4919_/A _4919_/B vssd1 vssd1 vccd1 vccd1 _4935_/S sky130_fd_sc_hd__or2_2
X_5899_ _5899_/A vssd1 vssd1 vccd1 vccd1 _7343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7638_ _7638_/CLK _7638_/D vssd1 vssd1 vccd1 vccd1 _7638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7569_ _7569_/CLK _7569_/D vssd1 vssd1 vccd1 vccd1 _7569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6769__154 _6769__154/A vssd1 vssd1 vccd1 vccd1 _7721_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116__334 _6116__334/A vssd1 vssd1 vccd1 vccd1 _7383_/CLK sky130_fd_sc_hd__inv_2
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6940_ _6924_/X _6939_/X _6872_/B vssd1 vssd1 vccd1 vccd1 _6940_/X sky130_fd_sc_hd__a21o_1
X_6871_ _6871_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _6872_/B sky130_fd_sc_hd__nand2_1
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6162__365 _6163__366/A vssd1 vssd1 vccd1 vccd1 _7417_/CLK sky130_fd_sc_hd__inv_2
X_4704_ _4704_/A vssd1 vssd1 vccd1 vccd1 _7317_/D sky130_fd_sc_hd__clkbuf_1
X_5684_ _5462_/A _5087_/A _5692_/S vssd1 vssd1 vccd1 vccd1 _5685_/A sky130_fd_sc_hd__mux2_1
X_4635_ _4635_/A vssd1 vssd1 vccd1 vccd1 _7380_/D sky130_fd_sc_hd__clkbuf_1
X_7423_ _7423_/CLK _7423_/D vssd1 vssd1 vccd1 vccd1 _7423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4566_ _4250_/X _7413_/Q _4570_/S vssd1 vssd1 vccd1 vccd1 _4567_/A sky130_fd_sc_hd__mux2_1
X_7354_ _7354_/CLK _7354_/D vssd1 vssd1 vccd1 vccd1 _7354_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7840_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3517_ _7218_/Q _7219_/Q _5446_/A _3517_/D vssd1 vssd1 vccd1 vccd1 _5458_/C sky130_fd_sc_hd__or4_4
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4497_ _4408_/X _7444_/Q _4497_/S vssd1 vssd1 vccd1 vccd1 _4498_/A sky130_fd_sc_hd__mux2_1
X_7285_ _7285_/CLK _7285_/D vssd1 vssd1 vccd1 vccd1 _7285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6236_ _7849_/Q _6871_/A _6871_/B vssd1 vssd1 vccd1 vccd1 _6236_/X sky130_fd_sc_hd__and3_1
X_6167_ _6167_/A vssd1 vssd1 vccd1 vccd1 _6167_/X sky130_fd_sc_hd__buf_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _7333_/Q _5120_/B vssd1 vssd1 vccd1 vccd1 _5119_/A sky130_fd_sc_hd__and2_1
XFILLER_111_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ _7594_/Q _7562_/Q _7837_/Q _7538_/Q _5983_/X _5984_/X vssd1 vssd1 vccd1 vccd1
+ _6099_/B sky130_fd_sc_hd__mux4_1
Xclkbuf_1_0_0__3302_ clkbuf_0__3302_/X vssd1 vssd1 vccd1 vccd1 _6779__161/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5049_ _5049_/A _5055_/B vssd1 vssd1 vccd1 vccd1 _5050_/A sky130_fd_sc_hd__or2_1
XFILLER_72_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3233_ clkbuf_0__3233_/X vssd1 vssd1 vccd1 vccd1 _6648__119/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5928__322 _5929__323/A vssd1 vssd1 vccd1 vccd1 _7363_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7857__231 vssd1 vssd1 vccd1 vccd1 partID[0] _7857__231/LO sky130_fd_sc_hd__conb_1
XFILLER_4_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4420_ _4578_/A vssd1 vssd1 vccd1 vccd1 _6328_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_8_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4351_ _4167_/X _7504_/Q _4355_/S vssd1 vssd1 vccd1 vccd1 _4352_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7070_ _7070_/A vssd1 vssd1 vccd1 vccd1 _7070_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4282_ _4731_/C _4284_/A _4281_/Y vssd1 vssd1 vccd1 vccd1 _7525_/D sky130_fd_sc_hd__o21a_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ _7622_/Q _7614_/Q _7606_/Q _7598_/Q _5933_/X _5998_/X vssd1 vssd1 vccd1 vccd1
+ _6021_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6923_ _7797_/Q _6933_/B vssd1 vssd1 vccd1 vccd1 _6923_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3997_ _3935_/X _7632_/Q _4001_/S vssd1 vssd1 vccd1 vccd1 _3998_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5736_ _5736_/A vssd1 vssd1 vccd1 vccd1 _7227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5667_ _5667_/A _5667_/B vssd1 vssd1 vccd1 vccd1 _5668_/A sky130_fd_sc_hd__or2_1
Xclkbuf_1_1_0__2448_ clkbuf_0__2448_/X vssd1 vssd1 vccd1 vccd1 _5368__198/A sky130_fd_sc_hd__clkbuf_4
X_4618_ _3657_/X _7387_/Q _4624_/S vssd1 vssd1 vccd1 vccd1 _4619_/A sky130_fd_sc_hd__mux2_1
X_7406_ _7855_/CLK _7406_/D vssd1 vssd1 vccd1 vccd1 _7406_/Q sky130_fd_sc_hd__dfxtp_1
X_5598_ _7182_/Q _7363_/Q _7719_/Q _7259_/Q _5427_/A _5472_/X vssd1 vssd1 vccd1 vccd1
+ _5598_/X sky130_fd_sc_hd__mux4_1
X_7337_ _7339_/CLK _7337_/D vssd1 vssd1 vccd1 vccd1 _7337_/Q sky130_fd_sc_hd__dfxtp_1
X_4549_ _4549_/A vssd1 vssd1 vccd1 vccd1 _7421_/D sky130_fd_sc_hd__clkbuf_1
X_7268_ _7268_/CLK _7268_/D vssd1 vssd1 vccd1 vccd1 _7268_/Q sky130_fd_sc_hd__dfxtp_1
X_6219_ _6879_/A _6879_/B _7095_/B vssd1 vssd1 vccd1 vccd1 _6219_/Y sky130_fd_sc_hd__a21oi_1
X_7199_ _7838_/CLK _7199_/D vssd1 vssd1 vccd1 vccd1 _7199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_10 _4233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_32 _5098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_43 _4817_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_21 _5162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3147_ clkbuf_0__3147_/X vssd1 vssd1 vccd1 vccd1 _6548__107/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5835__290 _5839__294/A vssd1 vssd1 vccd1 vccd1 _7307_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3920_ _3832_/X _7663_/Q _3924_/S vssd1 vssd1 vccd1 vccd1 _3921_/A sky130_fd_sc_hd__mux2_1
X_3851_ _3709_/X _7709_/Q _3853_/S vssd1 vssd1 vccd1 vccd1 _3852_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6570_ _7677_/Q vssd1 vssd1 vccd1 vccd1 _6602_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3782_ _3782_/A vssd1 vssd1 vccd1 vccd1 _7721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5521_ _5521_/A vssd1 vssd1 vccd1 vccd1 _5521_/X sky130_fd_sc_hd__clkbuf_4
X_5452_ _7092_/B vssd1 vssd1 vccd1 vccd1 _5453_/A sky130_fd_sc_hd__clkbuf_2
X_4403_ _4402_/X _7483_/Q _4409_/S vssd1 vssd1 vccd1 vccd1 _4404_/A sky130_fd_sc_hd__mux2_1
X_5383_ _5758_/A vssd1 vssd1 vccd1 vccd1 _5383_/X sky130_fd_sc_hd__buf_1
XFILLER_113_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7122_ _7372_/CLK _7122_/D vssd1 vssd1 vccd1 vccd1 _7122_/Q sky130_fd_sc_hd__dfxtp_1
X_4334_ _4334_/A vssd1 vssd1 vccd1 vccd1 _7512_/D sky130_fd_sc_hd__clkbuf_1
X_7053_ _7053_/A vssd1 vssd1 vccd1 vccd1 _7840_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6004_ _5999_/X _6000_/X _6001_/X _6003_/X _5945_/X _5947_/X vssd1 vssd1 vccd1 vccd1
+ _6004_/X sky130_fd_sc_hd__mux4_2
X_4265_ _7822_/Q vssd1 vssd1 vccd1 vccd1 _4265_/X sky130_fd_sc_hd__buf_2
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4196_ _4211_/S vssd1 vssd1 vccd1 vccd1 _4205_/S sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__2997_ clkbuf_0__2997_/X vssd1 vssd1 vccd1 vccd1 _6169__371/A sky130_fd_sc_hd__clkbuf_4
X_6812__13 _6812__13/A vssd1 vssd1 vccd1 vccd1 _7755_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6129__344 _6129__344/A vssd1 vssd1 vccd1 vccd1 _7393_/CLK sky130_fd_sc_hd__inv_2
X_6906_ _6906_/A vssd1 vssd1 vccd1 vccd1 _7793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5719_ _7220_/Q _7335_/Q _5725_/S vssd1 vssd1 vccd1 vccd1 _5720_/A sky130_fd_sc_hd__mux2_1
X_6699_ _6711_/A _6699_/B _6699_/C _6705_/D vssd1 vssd1 vccd1 vccd1 _6699_/X sky130_fd_sc_hd__and4_1
XFILLER_40_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6646__117 _6648__119/A vssd1 vssd1 vccd1 vccd1 _7664_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4050_ _4050_/A vssd1 vssd1 vccd1 vccd1 _7610_/D sky130_fd_sc_hd__clkbuf_1
Xinput6 caravel_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__2782_ clkbuf_0__2782_/X vssd1 vssd1 vccd1 vccd1 _5911__309/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7740_ _7740_/CLK _7740_/D vssd1 vssd1 vccd1 vccd1 _7740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4952_ _4952_/A vssd1 vssd1 vccd1 vccd1 _7169_/D sky130_fd_sc_hd__clkbuf_1
X_7671_ _7845_/CLK _7671_/D vssd1 vssd1 vccd1 vccd1 _7671_/Q sky130_fd_sc_hd__dfxtp_1
X_3903_ _3836_/X _7689_/Q _3905_/S vssd1 vssd1 vccd1 vccd1 _3904_/A sky130_fd_sc_hd__mux2_1
X_4883_ _4883_/A _4937_/B vssd1 vssd1 vccd1 vccd1 _4899_/S sky130_fd_sc_hd__nand2_2
X_6622_ _6594_/A _6569_/A _6621_/D _7679_/Q vssd1 vssd1 vccd1 vccd1 _6699_/C sky130_fd_sc_hd__a31o_1
XFILLER_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3834_ _3834_/A vssd1 vssd1 vccd1 vccd1 _7715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3765_ _4596_/A _4523_/B vssd1 vssd1 vccd1 vccd1 _3781_/S sky130_fd_sc_hd__nand2_2
X_3696_ _3578_/X _7753_/Q _3696_/S vssd1 vssd1 vccd1 vccd1 _3697_/A sky130_fd_sc_hd__mux2_1
X_5504_ _7303_/Q _7231_/Q _7699_/Q _7319_/Q _5426_/A _4300_/A vssd1 vssd1 vccd1 vccd1
+ _5504_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_0__3302_ _6777_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3302_/X sky130_fd_sc_hd__clkbuf_16
X_5435_ _7207_/Q _5435_/B _7206_/Q vssd1 vssd1 vccd1 vccd1 _5446_/B sky130_fd_sc_hd__or3b_1
Xclkbuf_0__3233_ _6643_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3233_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_113_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5297_ _5295_/X _7335_/Q _5291_/X _5292_/X _7135_/Q vssd1 vssd1 vccd1 vccd1 _7135_/D
+ sky130_fd_sc_hd__o32a_1
X_7105_ _7105_/A _7105_/B _7105_/C vssd1 vssd1 vccd1 vccd1 _7106_/C sky130_fd_sc_hd__and3_1
X_4317_ _7530_/Q _5396_/A _4305_/A vssd1 vssd1 vccd1 vccd1 _4318_/B sky130_fd_sc_hd__a21o_1
X_4248_ _4247_/X _7537_/Q _4257_/S vssd1 vssd1 vccd1 vccd1 _4249_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4179_ _4179_/A vssd1 vssd1 vccd1 vccd1 _7562_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6474__529 _6474__529/A vssd1 vssd1 vccd1 vccd1 _7594_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6763__149 _6763__149/A vssd1 vssd1 vccd1 vccd1 _7716_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6368__445 _6372__449/A vssd1 vssd1 vccd1 vccd1 _7508_/CLK sky130_fd_sc_hd__inv_2
X_6110__329 _6110__329/A vssd1 vssd1 vccd1 vccd1 _7378_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3550_ _3579_/S vssd1 vssd1 vccd1 vccd1 _3567_/S sky130_fd_sc_hd__buf_2
X_5220_ _5217_/X _5220_/B vssd1 vssd1 vccd1 vccd1 _5220_/X sky130_fd_sc_hd__and2b_1
XFILLER_111_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5151_ _7184_/Q _5161_/B _5215_/A vssd1 vssd1 vccd1 vccd1 _5151_/X sky130_fd_sc_hd__and3_1
X_5082_ _5082_/A vssd1 vssd1 vccd1 vccd1 _5082_/X sky130_fd_sc_hd__clkbuf_1
X_4102_ _4063_/X _7589_/Q _4106_/S vssd1 vssd1 vccd1 vccd1 _4103_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4033_ _4033_/A vssd1 vssd1 vccd1 vccd1 _7617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2765_ clkbuf_0__2765_/X vssd1 vssd1 vccd1 vccd1 _5769__238/A sky130_fd_sc_hd__clkbuf_4
X_5984_ _6031_/A vssd1 vssd1 vccd1 vccd1 _5984_/X sky130_fd_sc_hd__clkbuf_4
X_7723_ _7723_/CLK _7723_/D vssd1 vssd1 vccd1 vccd1 _7723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4935_ _4239_/X _7176_/Q _4935_/S vssd1 vssd1 vccd1 vccd1 _4936_/A sky130_fd_sc_hd__mux2_1
X_7654_ _7654_/CLK _7654_/D vssd1 vssd1 vccd1 vccd1 _7654_/Q sky130_fd_sc_hd__dfxtp_1
X_4866_ _4881_/S vssd1 vssd1 vccd1 vccd1 _4875_/S sky130_fd_sc_hd__buf_2
X_6605_ _6605_/A _6693_/B _6693_/C vssd1 vssd1 vccd1 vccd1 _6605_/Y sky130_fd_sc_hd__nand3_1
X_3817_ _3816_/X _7719_/Q _3829_/S vssd1 vssd1 vccd1 vccd1 _3818_/A sky130_fd_sc_hd__mux2_1
X_7585_ _7585_/CLK _7585_/D vssd1 vssd1 vccd1 vccd1 _7585_/Q sky130_fd_sc_hd__dfxtp_1
X_4797_ _4722_/X _7279_/Q _4801_/S vssd1 vssd1 vccd1 vccd1 _4798_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3317_ clkbuf_0__3317_/X vssd1 vssd1 vccd1 vccd1 _6858__50/A sky130_fd_sc_hd__clkbuf_4
X_3748_ _3698_/X _7736_/Q _3756_/S vssd1 vssd1 vccd1 vccd1 _3749_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5922__317 _5924__319/A vssd1 vssd1 vccd1 vccd1 _7358_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3679_ _4009_/B _3745_/A _4009_/A vssd1 vssd1 vccd1 vccd1 _3928_/B sky130_fd_sc_hd__or3b_2
Xoutput140 _5072_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[26] sky130_fd_sc_hd__buf_2
Xoutput151 _5030_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[7] sky130_fd_sc_hd__buf_2
X_5418_ _7237_/Q _7168_/Q _7478_/Q _7245_/Q _4297_/A _4305_/A vssd1 vssd1 vccd1 vccd1
+ _5418_/X sky130_fd_sc_hd__mux4_1
XFILLER_102_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5349_ _7659_/Q vssd1 vssd1 vccd1 vccd1 _6668_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_87_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput184 _5233_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[30] sky130_fd_sc_hd__buf_2
Xoutput162 _5180_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[10] sky130_fd_sc_hd__buf_2
Xoutput173 _5210_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[20] sky130_fd_sc_hd__buf_2
XFILLER_0_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3147_ _6545_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3147_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7019_ _7019_/A vssd1 vssd1 vccd1 vccd1 _7823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4719_/X _7312_/Q _4720_/S vssd1 vssd1 vccd1 vccd1 _4721_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4651_ _4666_/S vssd1 vssd1 vccd1 vccd1 _4660_/S sky130_fd_sc_hd__buf_2
Xinput31 caravel_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_2
Xinput20 caravel_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 _5222_/B sky130_fd_sc_hd__clkbuf_1
X_3602_ _3566_/X _7788_/Q _3602_/S vssd1 vssd1 vccd1 vccd1 _3603_/A sky130_fd_sc_hd__mux2_1
X_4582_ _7403_/Q _3932_/A _4588_/S vssd1 vssd1 vccd1 vccd1 _4583_/A sky130_fd_sc_hd__mux2_1
X_7370_ _7838_/CLK _7370_/D vssd1 vssd1 vccd1 vccd1 _7370_/Q sky130_fd_sc_hd__dfxtp_1
Xinput42 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 _5114_/A sky130_fd_sc_hd__buf_4
Xinput53 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 _5337_/C sky130_fd_sc_hd__buf_8
Xinput64 wbs_data_i[19] vssd1 vssd1 vccd1 vccd1 _5055_/A sky130_fd_sc_hd__buf_4
X_3533_ _4447_/B _4447_/C _4448_/C vssd1 vssd1 vccd1 vccd1 _3545_/A sky130_fd_sc_hd__mux2_1
Xinput75 wbs_data_i[29] vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__buf_4
Xinput86 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 _5318_/A sky130_fd_sc_hd__buf_8
X_6321_ _7820_/Q _6394_/C vssd1 vssd1 vccd1 vccd1 _6322_/A sky130_fd_sc_hd__and2_1
XFILLER_115_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6252_ _7840_/Q _6972_/A vssd1 vssd1 vccd1 vccd1 _6993_/A sky130_fd_sc_hd__xor2_1
X_5203_ _5216_/A vssd1 vssd1 vccd1 vccd1 _5204_/A sky130_fd_sc_hd__buf_2
X_6183_ _7807_/Q _6228_/B _6197_/A _6192_/C vssd1 vssd1 vccd1 vccd1 _6188_/B sky130_fd_sc_hd__and4_1
X_5134_ _5134_/A vssd1 vssd1 vccd1 vccd1 _5134_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5065_ _5065_/A vssd1 vssd1 vccd1 vccd1 _5065_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4016_ _3935_/X _7624_/Q _4020_/S vssd1 vssd1 vccd1 vccd1 _4017_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7881__208 vssd1 vssd1 vccd1 vccd1 _7881__208/HI manufacturerID[0] sky130_fd_sc_hd__conb_1
X_5967_ _5932_/X _5948_/X _5993_/A _5966_/X vssd1 vssd1 vccd1 vccd1 _5967_/X sky130_fd_sc_hd__a211o_2
X_7706_ _7706_/CLK _7706_/D vssd1 vssd1 vccd1 vccd1 _7706_/Q sky130_fd_sc_hd__dfxtp_1
X_4918_ _4918_/A vssd1 vssd1 vccd1 vccd1 _7229_/D sky130_fd_sc_hd__clkbuf_1
X_5898_ _7343_/Q _5071_/A _5902_/S vssd1 vssd1 vccd1 vccd1 _5899_/A sky130_fd_sc_hd__mux2_1
X_7637_ _7637_/CLK _7637_/D vssd1 vssd1 vccd1 vccd1 _7637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4849_ _4803_/X _7260_/Q _4857_/S vssd1 vssd1 vccd1 vccd1 _4850_/A sky130_fd_sc_hd__mux2_1
X_7568_ _7568_/CLK _7568_/D vssd1 vssd1 vccd1 vccd1 _7568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7499_ _7499_/CLK _7499_/D vssd1 vssd1 vccd1 vccd1 _7499_/Q sky130_fd_sc_hd__dfxtp_1
X_5822__281 _5824__283/A vssd1 vssd1 vccd1 vccd1 _7298_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6533__95 _6535__97/A vssd1 vssd1 vccd1 vccd1 _7640_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6870_ _7840_/Q _6870_/B vssd1 vssd1 vccd1 vccd1 _6870_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6776__159 _6776__159/A vssd1 vssd1 vccd1 vccd1 _7726_/CLK sky130_fd_sc_hd__inv_2
X_5752_ _5758_/A vssd1 vssd1 vccd1 vccd1 _5752_/X sky130_fd_sc_hd__buf_1
X_4703_ _4417_/X _7317_/Q _4703_/S vssd1 vssd1 vccd1 vccd1 _4704_/A sky130_fd_sc_hd__mux2_1
X_6123__339 _6123__339/A vssd1 vssd1 vccd1 vccd1 _7388_/CLK sky130_fd_sc_hd__inv_2
X_5683_ _5727_/A vssd1 vssd1 vccd1 vccd1 _5692_/S sky130_fd_sc_hd__buf_2
X_7422_ _7422_/CLK _7422_/D vssd1 vssd1 vccd1 vccd1 _7422_/Q sky130_fd_sc_hd__dfxtp_1
X_4634_ _3649_/X _7380_/Q _4642_/S vssd1 vssd1 vccd1 vccd1 _4635_/A sky130_fd_sc_hd__mux2_1
X_4565_ _4565_/A vssd1 vssd1 vccd1 vccd1 _7414_/D sky130_fd_sc_hd__clkbuf_1
X_7353_ _7353_/CLK _7353_/D vssd1 vssd1 vccd1 vccd1 _7353_/Q sky130_fd_sc_hd__dfxtp_1
X_3516_ _7220_/Q _7221_/Q _7222_/Q _7223_/Q vssd1 vssd1 vccd1 vccd1 _3517_/D sky130_fd_sc_hd__or4_1
X_6819__19 _6819__19/A vssd1 vssd1 vccd1 vccd1 _7761_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4496_ _4496_/A vssd1 vssd1 vccd1 vccd1 _7445_/D sky130_fd_sc_hd__clkbuf_1
X_7284_ _7284_/CLK _7284_/D vssd1 vssd1 vccd1 vccd1 _7284_/Q sky130_fd_sc_hd__dfxtp_1
X_6235_ _6871_/A _6871_/B _7849_/Q vssd1 vssd1 vccd1 vccd1 _6235_/Y sky130_fd_sc_hd__a21oi_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _5117_/A vssd1 vssd1 vccd1 vccd1 _5117_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6097_ _7792_/Q _7784_/Q _7776_/Q _7768_/Q _6031_/X _5980_/X vssd1 vssd1 vccd1 vccd1
+ _6097_/X sky130_fd_sc_hd__mux4_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5048_ _5048_/A vssd1 vssd1 vccd1 vccd1 _5048_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3301_ clkbuf_0__3301_/X vssd1 vssd1 vccd1 vccd1 _6776__159/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6999_ _7815_/Q _6995_/X _6998_/X _6909_/X vssd1 vssd1 vccd1 vccd1 _7814_/D sky130_fd_sc_hd__o211a_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4350_ _4350_/A vssd1 vssd1 vccd1 vccd1 _7505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4281_ _4731_/C _4284_/A _6396_/A vssd1 vssd1 vccd1 vccd1 _4281_/Y sky130_fd_sc_hd__a21oi_1
X_6020_ _7367_/Q _5931_/X _6019_/X _5996_/X vssd1 vssd1 vccd1 vccd1 _7367_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6922_ _6918_/Y _6920_/X _7014_/A vssd1 vssd1 vccd1 vccd1 _7796_/D sky130_fd_sc_hd__a21oi_1
XFILLER_81_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3996_ _3996_/A vssd1 vssd1 vccd1 vccd1 _7633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5735_ _5735_/A _5735_/B _5735_/C vssd1 vssd1 vccd1 vccd1 _5736_/A sky130_fd_sc_hd__and3_1
X_5666_ _7840_/Q _5649_/X _5638_/A _7199_/Q _7105_/B vssd1 vssd1 vccd1 vccd1 _5667_/B
+ sky130_fd_sc_hd__a32o_1
Xclkbuf_1_1_0__2447_ clkbuf_0__2447_/X vssd1 vssd1 vccd1 vccd1 _5363__194/A sky130_fd_sc_hd__clkbuf_4
X_4617_ _4617_/A vssd1 vssd1 vccd1 vccd1 _7388_/D sky130_fd_sc_hd__clkbuf_1
X_7405_ _7839_/CLK _7405_/D vssd1 vssd1 vccd1 vccd1 _7405_/Q sky130_fd_sc_hd__dfxtp_1
X_5597_ _5466_/X _5596_/X _5404_/A vssd1 vssd1 vccd1 vccd1 _5597_/X sky130_fd_sc_hd__a21o_1
X_7336_ _7336_/CLK _7336_/D vssd1 vssd1 vccd1 vccd1 _7336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4548_ _4250_/X _7421_/Q _4552_/S vssd1 vssd1 vccd1 vccd1 _4549_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4479_ _4408_/X _7452_/Q _4479_/S vssd1 vssd1 vccd1 vccd1 _4480_/A sky130_fd_sc_hd__mux2_1
X_7267_ _7267_/CLK _7267_/D vssd1 vssd1 vccd1 vccd1 _7267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6218_ _7853_/Q _6879_/A _6879_/B vssd1 vssd1 vccd1 vccd1 _6218_/X sky130_fd_sc_hd__and3_1
X_7198_ _7840_/CLK _7198_/D vssd1 vssd1 vccd1 vccd1 _7198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_22 _5085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6149_ _6149_/A vssd1 vssd1 vccd1 vccd1 _7407_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_33 _5337_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7887__214 vssd1 vssd1 vccd1 vccd1 _7887__214/HI manufacturerID[6] sky130_fd_sc_hd__conb_1
XINSDIODE2_11 _4803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_44 _7100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3146_ clkbuf_0__3146_/X vssd1 vssd1 vccd1 vccd1 _6551_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3850_ _3850_/A vssd1 vssd1 vccd1 vccd1 _7710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3781_ _3721_/X _7721_/Q _3781_/S vssd1 vssd1 vccd1 vccd1 _3782_/A sky130_fd_sc_hd__mux2_1
X_5520_ _5520_/A vssd1 vssd1 vccd1 vccd1 _5520_/X sky130_fd_sc_hd__clkbuf_4
X_5451_ _7855_/Q _5394_/Y _5442_/Y _5450_/X vssd1 vssd1 vccd1 vccd1 _7184_/D sky130_fd_sc_hd__a211o_1
XFILLER_8_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4402_ _4402_/A vssd1 vssd1 vccd1 vccd1 _4402_/X sky130_fd_sc_hd__buf_2
X_5382_ _5382_/A vssd1 vssd1 vccd1 vccd1 _5382_/X sky130_fd_sc_hd__buf_1
XFILLER_99_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7121_ _7154_/CLK _7121_/D vssd1 vssd1 vccd1 vccd1 _7121_/Q sky130_fd_sc_hd__dfxtp_1
X_4333_ _4167_/X _7512_/Q _4337_/S vssd1 vssd1 vccd1 vccd1 _4334_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7052_ _7048_/X _7052_/B vssd1 vssd1 vccd1 vccd1 _7053_/A sky130_fd_sc_hd__and2b_1
X_4264_ _4264_/A vssd1 vssd1 vccd1 vccd1 _7532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6003_ _7573_/Q _7383_/Q _7731_/Q _7629_/Q _6002_/X _4465_/X vssd1 vssd1 vccd1 vccd1
+ _6003_/X sky130_fd_sc_hd__mux4_1
X_4195_ _4937_/A _4217_/B vssd1 vssd1 vccd1 vccd1 _4211_/S sky130_fd_sc_hd__nand2_4
Xclkbuf_1_1_0__2996_ clkbuf_0__2996_/X vssd1 vssd1 vccd1 vccd1 _6166__369/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6905_ _7003_/A _6905_/B _6905_/C vssd1 vssd1 vccd1 vccd1 _6906_/A sky130_fd_sc_hd__and3_1
XFILLER_63_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3979_ _7640_/Q _3660_/X _3983_/S vssd1 vssd1 vccd1 vccd1 _3980_/A sky130_fd_sc_hd__mux2_1
X_5718_ _5718_/A vssd1 vssd1 vccd1 vccd1 _7219_/D sky130_fd_sc_hd__clkbuf_1
X_6402__470 _6404__472/A vssd1 vssd1 vccd1 vccd1 _7535_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6698_ _6656_/X _6658_/X _7679_/Q vssd1 vssd1 vccd1 vccd1 _6698_/Y sky130_fd_sc_hd__a21boi_1
X_5649_ _5649_/A vssd1 vssd1 vccd1 vccd1 _5649_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6175__376 _6178__379/A vssd1 vssd1 vccd1 vccd1 _7428_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7319_ _7319_/CLK _7319_/D vssd1 vssd1 vccd1 vccd1 _7319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5778__245 _5779__246/A vssd1 vssd1 vccd1 vccd1 _7262_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3129_ clkbuf_0__3129_/X vssd1 vssd1 vccd1 vccd1 _6462__519/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput7 caravel_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__2781_ clkbuf_0__2781_/X vssd1 vssd1 vccd1 vccd1 _5849__302/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4951_ _4236_/X _7169_/Q _4953_/S vssd1 vssd1 vccd1 vccd1 _4952_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7670_ _7845_/CLK _7670_/D vssd1 vssd1 vccd1 vccd1 _7670_/Q sky130_fd_sc_hd__dfxtp_1
X_3902_ _3902_/A vssd1 vssd1 vccd1 vccd1 _7690_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4882_ _4882_/A vssd1 vssd1 vccd1 vccd1 _7245_/D sky130_fd_sc_hd__clkbuf_1
X_6621_ _7679_/Q _6621_/B _6621_/C _6621_/D vssd1 vssd1 vccd1 vccd1 _6699_/B sky130_fd_sc_hd__nand4_1
X_3833_ _3832_/X _7715_/Q _3841_/S vssd1 vssd1 vccd1 vccd1 _3834_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3764_ _4009_/B _4614_/C _4614_/A vssd1 vssd1 vccd1 vccd1 _4523_/B sky130_fd_sc_hd__and3b_2
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3695_ _3695_/A vssd1 vssd1 vccd1 vccd1 _7754_/D sky130_fd_sc_hd__clkbuf_1
X_5503_ _7663_/Q _7496_/Q _7451_/Q _7311_/Q _5502_/X _5416_/A vssd1 vssd1 vccd1 vccd1
+ _5503_/X sky130_fd_sc_hd__mux4_1
X_6483_ _6501_/A vssd1 vssd1 vccd1 vccd1 _6483_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__3301_ _6771_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3301_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_10_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5434_ _5434_/A _5434_/B vssd1 vssd1 vccd1 vccd1 _5434_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7104_ _7104_/A _7104_/B vssd1 vssd1 vccd1 vccd1 _7106_/B sky130_fd_sc_hd__nor2_1
XFILLER_114_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5296_ _5295_/X _7334_/Q _5291_/X _5292_/X _7134_/Q vssd1 vssd1 vccd1 vccd1 _7134_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_99_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4316_ _4316_/A _4316_/B vssd1 vssd1 vccd1 vccd1 _7519_/D sky130_fd_sc_hd__nor2_1
XFILLER_101_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4247_ _7828_/Q vssd1 vssd1 vccd1 vccd1 _4247_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4178_ _4046_/X _7562_/Q _4186_/S vssd1 vssd1 vccd1 vccd1 _4179_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7826_/CLK
+ sky130_fd_sc_hd__clkbuf_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7799_ _7799_/CLK _7799_/D vssd1 vssd1 vccd1 vccd1 _7799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6485__56 _6486__57/A vssd1 vssd1 vccd1 vccd1 _7601_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6409__476 _6409__476/A vssd1 vssd1 vccd1 vccd1 _7541_/CLK sky130_fd_sc_hd__inv_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5150_ _5236_/B vssd1 vssd1 vccd1 vccd1 _5215_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5081_ _5081_/A _5081_/B vssd1 vssd1 vccd1 vccd1 _5082_/A sky130_fd_sc_hd__or2_1
XFILLER_110_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4101_ _4101_/A vssd1 vssd1 vccd1 vccd1 _7590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4032_ _3932_/X _7617_/Q _4038_/S vssd1 vssd1 vccd1 vccd1 _4033_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5983_ _7458_/Q vssd1 vssd1 vccd1 vccd1 _5983_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__2764_ clkbuf_0__2764_/X vssd1 vssd1 vccd1 vccd1 _5789_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7722_ _7722_/CLK _7722_/D vssd1 vssd1 vccd1 vccd1 _7722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4934_ _4934_/A vssd1 vssd1 vccd1 vccd1 _7177_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_19_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7684_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_7653_ _7653_/CLK _7653_/D vssd1 vssd1 vccd1 vccd1 _7653_/Q sky130_fd_sc_hd__dfxtp_1
X_4865_ _4865_/A _4865_/B _4937_/B vssd1 vssd1 vccd1 vccd1 _4881_/S sky130_fd_sc_hd__and3_2
X_6604_ _6693_/B _6693_/C _6605_/A vssd1 vssd1 vccd1 vccd1 _6604_/X sky130_fd_sc_hd__a21o_1
X_4796_ _4796_/A vssd1 vssd1 vccd1 vccd1 _7280_/D sky130_fd_sc_hd__clkbuf_1
X_7584_ _7584_/CLK _7584_/D vssd1 vssd1 vccd1 vccd1 _7584_/Q sky130_fd_sc_hd__dfxtp_1
X_3816_ _4399_/A vssd1 vssd1 vccd1 vccd1 _3816_/X sky130_fd_sc_hd__buf_2
XFILLER_20_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3316_ clkbuf_0__3316_/X vssd1 vssd1 vccd1 vccd1 _6855__48/A sky130_fd_sc_hd__clkbuf_4
X_3747_ _3762_/S vssd1 vssd1 vccd1 vccd1 _3756_/S sky130_fd_sc_hd__buf_2
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3678_ _3678_/A _3724_/A _3927_/B _3927_/C vssd1 vssd1 vccd1 vccd1 _4131_/D sky130_fd_sc_hd__or4_4
Xoutput141 _5074_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[27] sky130_fd_sc_hd__buf_2
Xoutput130 _5052_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[17] sky130_fd_sc_hd__buf_2
Xoutput152 _5032_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[8] sky130_fd_sc_hd__buf_2
X_5417_ _7510_/Q _7502_/Q _7441_/Q _7433_/Q _5413_/X _5416_/X vssd1 vssd1 vccd1 vccd1
+ _5417_/X sky130_fd_sc_hd__mux4_1
X_5348_ _7687_/Q _5348_/B vssd1 vssd1 vccd1 vccd1 _5348_/X sky130_fd_sc_hd__and2b_1
Xoutput163 _5182_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[11] sky130_fd_sc_hd__buf_2
Xoutput185 _5235_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[31] sky130_fd_sc_hd__buf_2
Xoutput174 _5212_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[21] sky130_fd_sc_hd__buf_2
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3146_ _6544_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3146_/X sky130_fd_sc_hd__clkbuf_16
X_5279_ _5278_/X _7156_/Q _5274_/X _5275_/X _7124_/Q vssd1 vssd1 vccd1 vccd1 _7124_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_87_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7018_ _7100_/A _7024_/B vssd1 vssd1 vccd1 vccd1 _7019_/A sky130_fd_sc_hd__and2_1
XFILLER_47_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6480__534 _6480__534/A vssd1 vssd1 vccd1 vccd1 _7599_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6374__450 _6376__452/A vssd1 vssd1 vccd1 vccd1 _7513_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4650_ _4919_/A _4955_/A vssd1 vssd1 vccd1 vccd1 _4666_/S sky130_fd_sc_hd__or2_4
Xinput21 caravel_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 _5224_/B sky130_fd_sc_hd__clkbuf_1
Xinput10 caravel_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_1
X_3601_ _3601_/A vssd1 vssd1 vccd1 vccd1 _7789_/D sky130_fd_sc_hd__clkbuf_1
Xinput32 caravel_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__buf_2
X_4581_ _4581_/A vssd1 vssd1 vccd1 vccd1 _7404_/D sky130_fd_sc_hd__clkbuf_1
Xinput54 wbs_data_i[0] vssd1 vssd1 vccd1 vccd1 _7105_/A sky130_fd_sc_hd__buf_4
Xinput43 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 _5149_/A sky130_fd_sc_hd__buf_4
X_6320_ _6320_/A vssd1 vssd1 vccd1 vccd1 _7473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3532_ _3678_/A _7458_/Q vssd1 vssd1 vccd1 vccd1 _4448_/C sky130_fd_sc_hd__xnor2_2
Xinput65 wbs_data_i[1] vssd1 vssd1 vccd1 vccd1 _5015_/A sky130_fd_sc_hd__buf_6
Xinput87 wbs_sel_i[1] vssd1 vssd1 vccd1 vccd1 _5856_/A sky130_fd_sc_hd__buf_8
Xinput76 wbs_data_i[2] vssd1 vssd1 vccd1 vccd1 _3805_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6251_ _7810_/Q _6251_/B vssd1 vssd1 vccd1 vccd1 _6972_/A sky130_fd_sc_hd__xor2_2
X_5202_ _7202_/Q _5200_/A _5187_/A vssd1 vssd1 vccd1 vccd1 _5216_/A sky130_fd_sc_hd__a21o_1
XFILLER_88_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6182_ _7806_/Q _7805_/Q _7804_/Q _7803_/Q vssd1 vssd1 vccd1 vccd1 _6192_/C sky130_fd_sc_hd__and4_1
X_5133_ _7340_/Q _5142_/B vssd1 vssd1 vccd1 vccd1 _5134_/A sky130_fd_sc_hd__and2_1
XFILLER_111_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5064_ _5064_/A _5066_/B vssd1 vssd1 vccd1 vccd1 _5065_/A sky130_fd_sc_hd__or2_1
XFILLER_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4015_ _4015_/A vssd1 vssd1 vccd1 vccd1 _7625_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__2816_ clkbuf_0__2816_/X vssd1 vssd1 vccd1 vccd1 _6104__324/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5966_ _5960_/X _5965_/X _4452_/A vssd1 vssd1 vccd1 vccd1 _5966_/X sky130_fd_sc_hd__o21a_1
X_5897_ _5897_/A vssd1 vssd1 vccd1 vccd1 _7342_/D sky130_fd_sc_hd__clkbuf_1
X_7705_ _7705_/CLK _7705_/D vssd1 vssd1 vccd1 vccd1 _7705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4917_ _4826_/X _7229_/Q _4917_/S vssd1 vssd1 vccd1 vccd1 _4918_/A sky130_fd_sc_hd__mux2_1
X_7636_ _7636_/CLK _7636_/D vssd1 vssd1 vccd1 vccd1 _7636_/Q sky130_fd_sc_hd__dfxtp_1
X_4848_ _4863_/S vssd1 vssd1 vccd1 vccd1 _4857_/S sky130_fd_sc_hd__buf_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7567_ _7567_/CLK _7567_/D vssd1 vssd1 vccd1 vccd1 _7567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4779_ _4722_/X _7287_/Q _4783_/S vssd1 vssd1 vccd1 vccd1 _4780_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7498_ _7498_/CLK _7498_/D vssd1 vssd1 vccd1 vccd1 _7498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3129_ _6457_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3129_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_75_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5820_ _5820_/A vssd1 vssd1 vccd1 vccd1 _5820_/X sky130_fd_sc_hd__buf_1
XFILLER_34_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4702_ _4702_/A vssd1 vssd1 vccd1 vccd1 _7318_/D sky130_fd_sc_hd__clkbuf_1
X_7421_ _7421_/CLK _7421_/D vssd1 vssd1 vccd1 vccd1 _7421_/Q sky130_fd_sc_hd__dfxtp_1
X_5682_ _5682_/A _5682_/B _5682_/C vssd1 vssd1 vccd1 vccd1 _5727_/A sky130_fd_sc_hd__and3_4
X_4633_ _4648_/S vssd1 vssd1 vccd1 vccd1 _4642_/S sky130_fd_sc_hd__buf_2
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2394_ clkbuf_0__2394_/X vssd1 vssd1 vccd1 vccd1 _5357__189/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4564_ _4247_/X _7414_/Q _4570_/S vssd1 vssd1 vccd1 vccd1 _4565_/A sky130_fd_sc_hd__mux2_1
X_7352_ _7352_/CLK _7352_/D vssd1 vssd1 vccd1 vccd1 _7352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3515_ _7227_/Q _7226_/Q vssd1 vssd1 vccd1 vccd1 _5446_/A sky130_fd_sc_hd__nor2_4
X_7283_ _7283_/CLK _7283_/D vssd1 vssd1 vccd1 vccd1 _7283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6234_ _6933_/A _6930_/A _6245_/A _7801_/Q vssd1 vssd1 vccd1 vccd1 _6871_/B sky130_fd_sc_hd__a31o_1
X_4495_ _4405_/X _7445_/Q _4497_/S vssd1 vssd1 vccd1 vccd1 _4496_/A sky130_fd_sc_hd__mux2_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _7332_/Q _5120_/B vssd1 vssd1 vccd1 vccd1 _5117_/A sky130_fd_sc_hd__and2_1
X_6096_ _5978_/X _6093_/X _6095_/X _5964_/A vssd1 vssd1 vccd1 vccd1 _6096_/X sky130_fd_sc_hd__o211a_1
XFILLER_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5047_ _5047_/A _5055_/B vssd1 vssd1 vccd1 vccd1 _5048_/A sky130_fd_sc_hd__or2_1
Xclkbuf_1_0_0__3300_ clkbuf_0__3300_/X vssd1 vssd1 vccd1 vccd1 _6783_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_34_wb_clk_i _7474_/CLK vssd1 vssd1 vccd1 vccd1 _7819_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6998_ _6996_/X _6997_/X _7814_/Q vssd1 vssd1 vccd1 vccd1 _6998_/X sky130_fd_sc_hd__a21o_1
X_5949_ _7838_/Q _5949_/B vssd1 vssd1 vccd1 vccd1 _5950_/A sky130_fd_sc_hd__nand2_1
XFILLER_40_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7619_ _7619_/CLK _7619_/D vssd1 vssd1 vccd1 vccd1 _7619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6506__74 _6506__74/A vssd1 vssd1 vccd1 vccd1 _7619_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4280_ _4280_/A vssd1 vssd1 vccd1 vccd1 _6396_/A sky130_fd_sc_hd__buf_2
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6782__164 _6782__164/A vssd1 vssd1 vccd1 vccd1 _7731_/CLK sky130_fd_sc_hd__inv_2
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6824__23 _6825__24/A vssd1 vssd1 vccd1 vccd1 _7765_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6387__460 _6391__464/A vssd1 vssd1 vccd1 vccd1 _7523_/CLK sky130_fd_sc_hd__inv_2
X_6921_ _6954_/A vssd1 vssd1 vccd1 vccd1 _7014_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6783_ _6783_/A vssd1 vssd1 vccd1 vccd1 _6783_/X sky130_fd_sc_hd__buf_1
X_3995_ _3932_/X _7633_/Q _4001_/S vssd1 vssd1 vccd1 vccd1 _3996_/A sky130_fd_sc_hd__mux2_1
X_5847__300 _5849__302/A vssd1 vssd1 vccd1 vccd1 _7317_/CLK sky130_fd_sc_hd__inv_2
X_5734_ _4998_/A _5457_/X _5493_/C _5634_/B vssd1 vssd1 vccd1 vccd1 _5735_/C sky130_fd_sc_hd__o211ai_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5665_ _5665_/A vssd1 vssd1 vccd1 vccd1 _7198_/D sky130_fd_sc_hd__clkbuf_1
X_7404_ _7404_/CLK _7404_/D vssd1 vssd1 vccd1 vccd1 _7404_/Q sky130_fd_sc_hd__dfxtp_1
X_4616_ _3649_/X _7388_/Q _4624_/S vssd1 vssd1 vccd1 vccd1 _4617_/A sky130_fd_sc_hd__mux2_1
X_7335_ _7336_/CLK _7335_/D vssd1 vssd1 vccd1 vccd1 _7335_/Q sky130_fd_sc_hd__dfxtp_1
X_5596_ _7516_/Q _7508_/Q _7447_/Q _7439_/Q _5486_/X _5426_/X vssd1 vssd1 vccd1 vccd1
+ _5596_/X sky130_fd_sc_hd__mux4_2
X_4547_ _4547_/A vssd1 vssd1 vccd1 vccd1 _7422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7266_ _7266_/CLK _7266_/D vssd1 vssd1 vccd1 vccd1 _7266_/Q sky130_fd_sc_hd__dfxtp_1
X_4478_ _4478_/A vssd1 vssd1 vccd1 vccd1 _7453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7197_ _7329_/CLK _7197_/D vssd1 vssd1 vccd1 vccd1 _7197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6217_ _6918_/A _7795_/Q _7797_/Q vssd1 vssd1 vccd1 vccd1 _6879_/B sky130_fd_sc_hd__a21o_1
X_6148_ _7407_/Q _5874_/A _6148_/S vssd1 vssd1 vccd1 vccd1 _6149_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_23 _5085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_12 _5122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_34 _5036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _6079_/A _6079_/B vssd1 vssd1 vccd1 vccd1 _6079_/X sky130_fd_sc_hd__or2_1
XINSDIODE2_45 _7100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3145_ clkbuf_0__3145_/X vssd1 vssd1 vccd1 vccd1 _6543__104/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3780_ _3780_/A vssd1 vssd1 vccd1 vccd1 _7722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5450_ _7184_/Q _7092_/B _5647_/A vssd1 vssd1 vccd1 vccd1 _5450_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4401_ _4401_/A vssd1 vssd1 vccd1 vccd1 _7484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7120_ _7687_/CLK _7120_/D vssd1 vssd1 vccd1 vccd1 _7120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5842__296 _5843__297/A vssd1 vssd1 vccd1 vccd1 _7313_/CLK sky130_fd_sc_hd__inv_2
X_4332_ _4332_/A vssd1 vssd1 vccd1 vccd1 _7513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7051_ _5047_/A _7840_/Q _7067_/S vssd1 vssd1 vccd1 vccd1 _7052_/B sky130_fd_sc_hd__mux2_1
X_4263_ _4262_/X _7532_/Q _4266_/S vssd1 vssd1 vccd1 vccd1 _4264_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6002_ _6002_/A vssd1 vssd1 vccd1 vccd1 _6002_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4194_ _4194_/A _4194_/B _4865_/A vssd1 vssd1 vccd1 vccd1 _4937_/A sky130_fd_sc_hd__and3_4
Xclkbuf_1_1_0__2995_ clkbuf_0__2995_/X vssd1 vssd1 vccd1 vccd1 _6158__362/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6904_ _6916_/B _6939_/A _6904_/C vssd1 vssd1 vccd1 vccd1 _6905_/C sky130_fd_sc_hd__nand3_1
XFILLER_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3978_ _3978_/A vssd1 vssd1 vccd1 vccd1 _7641_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5717_ _7219_/Q _7334_/Q _5725_/S vssd1 vssd1 vccd1 vccd1 _5718_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6697_ _6695_/X _6696_/Y _6690_/X vssd1 vssd1 vccd1 vccd1 _7678_/D sky130_fd_sc_hd__a21oi_1
X_5648_ _7844_/Q vssd1 vssd1 vccd1 vccd1 _6242_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5579_ _5569_/X _5572_/X _5575_/X _5578_/X _4291_/A _7522_/Q vssd1 vssd1 vccd1 vccd1
+ _5579_/X sky130_fd_sc_hd__mux4_2
XFILLER_117_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7318_ _7318_/CLK _7318_/D vssd1 vssd1 vccd1 vccd1 _7318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7249_ _7249_/CLK _7249_/D vssd1 vssd1 vccd1 vccd1 _7249_/Q sky130_fd_sc_hd__dfxtp_1
X_6500__69 _6500__69/A vssd1 vssd1 vccd1 vccd1 _7614_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3128_ clkbuf_0__3128_/X vssd1 vssd1 vccd1 vccd1 _6455__513/A sky130_fd_sc_hd__clkbuf_4
X_6338__421 _6339__422/A vssd1 vssd1 vccd1 vccd1 _7484_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 caravel_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2780_ clkbuf_0__2780_/X vssd1 vssd1 vccd1 vccd1 _5845__299/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4950_ _4950_/A vssd1 vssd1 vccd1 vccd1 _7170_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3901_ _3832_/X _7690_/Q _3905_/S vssd1 vssd1 vccd1 vccd1 _3902_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4881_ _7245_/Q _4417_/A _4881_/S vssd1 vssd1 vccd1 vccd1 _4882_/A sky130_fd_sc_hd__mux2_1
X_6620_ _6705_/B _6705_/C _7843_/Q vssd1 vssd1 vccd1 vccd1 _6620_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3832_ _4411_/A vssd1 vssd1 vccd1 vccd1 _3832_/X sky130_fd_sc_hd__buf_2
XFILLER_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6551_ _6551_/A vssd1 vssd1 vccd1 vccd1 _6551_/X sky130_fd_sc_hd__buf_1
X_3763_ _3763_/A vssd1 vssd1 vccd1 vccd1 _7729_/D sky130_fd_sc_hd__clkbuf_1
X_5502_ _5520_/A vssd1 vssd1 vccd1 vccd1 _5502_/X sky130_fd_sc_hd__buf_6
X_3694_ _3574_/X _7754_/Q _3696_/S vssd1 vssd1 vccd1 vccd1 _3695_/A sky130_fd_sc_hd__mux2_1
X_6482_ _6739_/A vssd1 vssd1 vccd1 vccd1 _6482_/X sky130_fd_sc_hd__buf_1
XFILLER_106_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3300_ _6770_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3300_/X sky130_fd_sc_hd__clkbuf_16
X_5433_ _5429_/X _5432_/X _5433_/S vssd1 vssd1 vccd1 vccd1 _5434_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5364_ _5376_/A vssd1 vssd1 vccd1 vccd1 _5364_/X sky130_fd_sc_hd__buf_1
X_7103_ _7855_/Q vssd1 vssd1 vccd1 vccd1 _7104_/A sky130_fd_sc_hd__inv_2
X_4315_ _4312_/A _4312_/B _6308_/B vssd1 vssd1 vccd1 vccd1 _4316_/B sky130_fd_sc_hd__o21ai_1
XFILLER_114_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5295_ _5303_/A vssd1 vssd1 vccd1 vccd1 _5295_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4246_ _4246_/A vssd1 vssd1 vccd1 vccd1 _7538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4177_ _4192_/S vssd1 vssd1 vccd1 vccd1 _4186_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7798_ _7853_/CLK _7798_/D vssd1 vssd1 vccd1 vccd1 _7798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5784__250 _5785__251/A vssd1 vssd1 vccd1 vccd1 _7267_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5080_ _5080_/A vssd1 vssd1 vccd1 vccd1 _5080_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4100_ _4060_/X _7590_/Q _4100_/S vssd1 vssd1 vccd1 vccd1 _4101_/A sky130_fd_sc_hd__mux2_1
X_7872__199 vssd1 vssd1 vccd1 vccd1 _7872__199/HI core0Index[6] sky130_fd_sc_hd__conb_1
XFILLER_110_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4031_ _4031_/A vssd1 vssd1 vccd1 vccd1 _7618_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5982_ _6095_/A vssd1 vssd1 vccd1 vccd1 _6079_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2763_ clkbuf_0__2763_/X vssd1 vssd1 vccd1 vccd1 _5763__234/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7721_ _7721_/CLK _7721_/D vssd1 vssd1 vccd1 vccd1 _7721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4933_ _4236_/X _7177_/Q _4935_/S vssd1 vssd1 vccd1 vccd1 _4934_/A sky130_fd_sc_hd__mux2_1
X_7652_ _7652_/CLK _7652_/D vssd1 vssd1 vccd1 vccd1 _7652_/Q sky130_fd_sc_hd__dfxtp_1
X_4864_ _4864_/A vssd1 vssd1 vccd1 vccd1 _7253_/D sky130_fd_sc_hd__clkbuf_1
X_6603_ _6613_/A _6613_/B _6602_/A vssd1 vssd1 vccd1 vccd1 _6693_/C sky130_fd_sc_hd__a21o_1
X_7583_ _7583_/CLK _7583_/D vssd1 vssd1 vccd1 vccd1 _7583_/Q sky130_fd_sc_hd__dfxtp_1
X_4795_ _4719_/X _7280_/Q _4795_/S vssd1 vssd1 vccd1 vccd1 _4796_/A sky130_fd_sc_hd__mux2_1
X_3815_ _7474_/Q vssd1 vssd1 vccd1 vccd1 _4399_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0__3315_ clkbuf_0__3315_/X vssd1 vssd1 vccd1 vccd1 _6848__42/A sky130_fd_sc_hd__clkbuf_4
X_3746_ _4131_/A _4424_/A _3991_/C _4028_/A vssd1 vssd1 vccd1 vccd1 _3762_/S sky130_fd_sc_hd__or4_4
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3677_ _3677_/A vssd1 vssd1 vccd1 vccd1 _7761_/D sky130_fd_sc_hd__clkbuf_1
X_5416_ _5416_/A vssd1 vssd1 vccd1 vccd1 _5416_/X sky130_fd_sc_hd__buf_4
Xoutput142 _5076_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[28] sky130_fd_sc_hd__buf_2
Xoutput131 _5054_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[18] sky130_fd_sc_hd__buf_2
Xoutput120 _5104_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[9] sky130_fd_sc_hd__buf_2
X_6396_ _6396_/A _6396_/B vssd1 vssd1 vccd1 vccd1 _7530_/D sky130_fd_sc_hd__nor2_1
Xoutput153 _5034_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[9] sky130_fd_sc_hd__buf_2
X_5347_ _7365_/Q _7366_/Q _7367_/Q _7368_/Q _6718_/A _7686_/Q vssd1 vssd1 vccd1 vccd1
+ _5348_/B sky130_fd_sc_hd__mux4_1
Xoutput175 _5214_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[22] sky130_fd_sc_hd__buf_2
Xoutput186 _5158_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[3] sky130_fd_sc_hd__buf_2
Xoutput164 _5184_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[12] sky130_fd_sc_hd__buf_2
Xclkbuf_0__3145_ _6538_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3145_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5278_ _5303_/A vssd1 vssd1 vccd1 vccd1 _5278_/X sky130_fd_sc_hd__clkbuf_2
X_7017_ _7017_/A vssd1 vssd1 vccd1 vccd1 _7822_/D sky130_fd_sc_hd__clkbuf_1
X_4229_ _4229_/A vssd1 vssd1 vccd1 vccd1 _7543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6490__60 _6494__64/A vssd1 vssd1 vccd1 vccd1 _7605_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6415__481 _6418__484/A vssd1 vssd1 vccd1 vccd1 _7546_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 caravel_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 _5226_/B sky130_fd_sc_hd__clkbuf_1
Xinput11 caravel_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
X_3600_ _3562_/X _7789_/Q _3602_/S vssd1 vssd1 vccd1 vccd1 _3601_/A sky130_fd_sc_hd__mux2_1
X_4580_ _7404_/Q _3926_/A _4588_/S vssd1 vssd1 vccd1 vccd1 _4581_/A sky130_fd_sc_hd__mux2_1
Xinput33 caravel_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_2
X_3531_ _3585_/A _7457_/Q vssd1 vssd1 vccd1 vccd1 _4447_/C sky130_fd_sc_hd__and2b_1
Xinput44 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__buf_4
Xinput55 wbs_data_i[10] vssd1 vssd1 vccd1 vccd1 _5036_/A sky130_fd_sc_hd__buf_6
Xinput88 wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 _5874_/A sky130_fd_sc_hd__buf_8
Xinput66 wbs_data_i[20] vssd1 vssd1 vccd1 vccd1 _5058_/A sky130_fd_sc_hd__buf_4
Xinput77 wbs_data_i[30] vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__buf_4
X_6250_ _6866_/B _6250_/B _6250_/C vssd1 vssd1 vccd1 vccd1 _6253_/C sky130_fd_sc_hd__and3_1
X_5201_ _5200_/X _5201_/B vssd1 vssd1 vccd1 vccd1 _5201_/X sky130_fd_sc_hd__and2b_1
X_6181_ _7802_/Q _7801_/Q _7800_/Q _7799_/Q vssd1 vssd1 vccd1 vccd1 _6197_/A sky130_fd_sc_hd__and4_1
X_5132_ _5132_/A vssd1 vssd1 vccd1 vccd1 _5132_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5063_ _5063_/A vssd1 vssd1 vccd1 vccd1 _5063_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4014_ _3932_/X _7625_/Q _4020_/S vssd1 vssd1 vccd1 vccd1 _4015_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__2815_ clkbuf_0__2815_/X vssd1 vssd1 vccd1 vccd1 _5920__315/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5965_ _4451_/A _5961_/X _5963_/X _5964_/X vssd1 vssd1 vccd1 vccd1 _5965_/X sky130_fd_sc_hd__o211a_1
XFILLER_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5896_ _7342_/Q _5069_/A _5902_/S vssd1 vssd1 vccd1 vccd1 _5897_/A sky130_fd_sc_hd__mux2_1
X_7704_ _7704_/CLK _7704_/D vssd1 vssd1 vccd1 vccd1 _7704_/Q sky130_fd_sc_hd__dfxtp_1
X_4916_ _4916_/A vssd1 vssd1 vccd1 vccd1 _7230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7635_ _7635_/CLK _7635_/D vssd1 vssd1 vccd1 vccd1 _7635_/Q sky130_fd_sc_hd__dfxtp_1
X_4847_ _4919_/A _4847_/B vssd1 vssd1 vccd1 vccd1 _4863_/S sky130_fd_sc_hd__or2_2
XFILLER_107_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7566_ _7566_/CLK _7566_/D vssd1 vssd1 vccd1 vccd1 _7566_/Q sky130_fd_sc_hd__dfxtp_1
X_4778_ _4778_/A vssd1 vssd1 vccd1 vccd1 _7288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3729_ _3703_/X _7743_/Q _3735_/S vssd1 vssd1 vccd1 vccd1 _3730_/A sky130_fd_sc_hd__mux2_1
X_7497_ _7497_/CLK _7497_/D vssd1 vssd1 vccd1 vccd1 _7497_/Q sky130_fd_sc_hd__dfxtp_1
X_6379_ _6379_/A vssd1 vssd1 vccd1 vccd1 _6379_/X sky130_fd_sc_hd__buf_1
XFILLER_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__3128_ _6451_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3128_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_28_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6518__83 _6519__84/A vssd1 vssd1 vccd1 vccd1 _7628_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5797__260 _5799__262/A vssd1 vssd1 vccd1 vccd1 _7277_/CLK sky130_fd_sc_hd__inv_2
X_6836__32 _6836__32/A vssd1 vssd1 vccd1 vccd1 _7774_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5681_ _7203_/Q _5735_/A _5679_/Y _5680_/Y vssd1 vssd1 vccd1 vccd1 _7203_/D sky130_fd_sc_hd__o211a_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _4414_/X _7318_/Q _4703_/S vssd1 vssd1 vccd1 vccd1 _4702_/A sky130_fd_sc_hd__mux2_1
X_7420_ _7420_/CLK _7420_/D vssd1 vssd1 vccd1 vccd1 _7420_/Q sky130_fd_sc_hd__dfxtp_1
X_4632_ _4632_/A _4632_/B vssd1 vssd1 vccd1 vccd1 _4648_/S sky130_fd_sc_hd__nand2_2
Xclkbuf_1_1_0__2393_ clkbuf_0__2393_/X vssd1 vssd1 vccd1 vccd1 _5358_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4563_ _4563_/A vssd1 vssd1 vccd1 vccd1 _7415_/D sky130_fd_sc_hd__clkbuf_1
X_7351_ _7351_/CLK _7351_/D vssd1 vssd1 vccd1 vccd1 _7351_/Q sky130_fd_sc_hd__dfxtp_1
X_3514_ _5388_/A _5457_/A vssd1 vssd1 vccd1 vccd1 _5462_/B sky130_fd_sc_hd__and2_1
X_6302_ _6342_/A vssd1 vssd1 vccd1 vccd1 _6302_/X sky130_fd_sc_hd__buf_1
X_4494_ _4494_/A vssd1 vssd1 vccd1 vccd1 _7446_/D sky130_fd_sc_hd__clkbuf_1
X_7282_ _7282_/CLK _7282_/D vssd1 vssd1 vccd1 vccd1 _7282_/Q sky130_fd_sc_hd__dfxtp_1
X_6233_ _7801_/Q _6933_/A _6930_/A _6233_/D vssd1 vssd1 vccd1 vccd1 _6871_/A sky130_fd_sc_hd__nand4_1
XFILLER_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5115_/A vssd1 vssd1 vccd1 vccd1 _5115_/X sky130_fd_sc_hd__clkbuf_1
X_6095_ _6095_/A _6095_/B vssd1 vssd1 vccd1 vccd1 _6095_/X sky130_fd_sc_hd__or2_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5046_ _5068_/A vssd1 vssd1 vccd1 vccd1 _5055_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6997_ _6997_/A vssd1 vssd1 vccd1 vccd1 _6997_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5948_ _5934_/X _5938_/X _5941_/X _5943_/X _5945_/X _5947_/X vssd1 vssd1 vccd1 vccd1
+ _5948_/X sky130_fd_sc_hd__mux4_2
XFILLER_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5879_ _5879_/A vssd1 vssd1 vccd1 vccd1 _7334_/D sky130_fd_sc_hd__clkbuf_1
X_7618_ _7618_/CLK _7618_/D vssd1 vssd1 vccd1 vccd1 _7618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7549_ _7549_/CLK _7549_/D vssd1 vssd1 vccd1 vccd1 _7549_/Q sky130_fd_sc_hd__dfxtp_1
X_6332__416 _6333__417/A vssd1 vssd1 vccd1 vccd1 _7479_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7864__238 vssd1 vssd1 vccd1 vccd1 partID[14] _7864__238/LO sky130_fd_sc_hd__conb_1
X_6265__381 _6266__382/A vssd1 vssd1 vccd1 vccd1 _7434_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6809__10 _6813__14/A vssd1 vssd1 vccd1 vccd1 _7752_/CLK sky130_fd_sc_hd__inv_2
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6920_ _6912_/X _6919_/X _6878_/B vssd1 vssd1 vccd1 vccd1 _6920_/X sky130_fd_sc_hd__a21bo_1
X_6851_ _6857_/A vssd1 vssd1 vccd1 vccd1 _6851_/X sky130_fd_sc_hd__buf_1
X_6428__491 _6428__491/A vssd1 vssd1 vccd1 vccd1 _7556_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5802_ _5814_/A vssd1 vssd1 vccd1 vccd1 _5802_/X sky130_fd_sc_hd__buf_1
X_3994_ _3994_/A vssd1 vssd1 vccd1 vccd1 _7634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5733_ _4998_/A _5457_/X _5679_/Y _5735_/B vssd1 vssd1 vccd1 vccd1 _7226_/D sky130_fd_sc_hd__o211a_1
X_5664_ _5667_/A _5664_/B vssd1 vssd1 vccd1 vccd1 _5665_/A sky130_fd_sc_hd__or2_1
X_7403_ _7403_/CLK _7403_/D vssd1 vssd1 vccd1 vccd1 _7403_/Q sky130_fd_sc_hd__dfxtp_1
X_4615_ _4630_/S vssd1 vssd1 vccd1 vccd1 _4624_/S sky130_fd_sc_hd__clkbuf_2
X_5595_ _5611_/S _5595_/B vssd1 vssd1 vccd1 vccd1 _5595_/X sky130_fd_sc_hd__and2_1
X_7334_ _7336_/CLK _7334_/D vssd1 vssd1 vccd1 vccd1 _7334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4546_ _4247_/X _7422_/Q _4552_/S vssd1 vssd1 vccd1 vccd1 _4547_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4477_ _4405_/X _7453_/Q _4479_/S vssd1 vssd1 vccd1 vccd1 _4478_/A sky130_fd_sc_hd__mux2_1
X_7265_ _7265_/CLK _7265_/D vssd1 vssd1 vccd1 vccd1 _7265_/Q sky130_fd_sc_hd__dfxtp_1
X_7196_ _7840_/CLK _7196_/D vssd1 vssd1 vccd1 vccd1 _7196_/Q sky130_fd_sc_hd__dfxtp_1
X_6216_ _7797_/Q _6918_/A _7795_/Q vssd1 vssd1 vccd1 vccd1 _6879_/A sky130_fd_sc_hd__nand3_2
X_6147_ _6147_/A vssd1 vssd1 vccd1 vccd1 _7406_/D sky130_fd_sc_hd__clkbuf_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_24 _5085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_13 _5555_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _7395_/Q _7379_/Q _7649_/Q _7641_/Q _5936_/A _5933_/A vssd1 vssd1 vccd1 vccd1
+ _6079_/B sky130_fd_sc_hd__mux4_2
XFILLER_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_35 _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_46 _5537_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5029_ _7030_/A _5033_/B vssd1 vssd1 vccd1 vccd1 _5030_/A sky130_fd_sc_hd__or2_1
XFILLER_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3144_ clkbuf_0__3144_/X vssd1 vssd1 vccd1 vccd1 _6537__99/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6759__145 _6760__146/A vssd1 vssd1 vccd1 vccd1 _7712_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6106__325 _6108__327/A vssd1 vssd1 vccd1 vccd1 _7374_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5748__221 _5749__222/A vssd1 vssd1 vccd1 vccd1 _7238_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4400_ _4399_/X _7484_/Q _4409_/S vssd1 vssd1 vccd1 vccd1 _4401_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4331_ _4164_/X _7513_/Q _4331_/S vssd1 vssd1 vccd1 vccd1 _4332_/A sky130_fd_sc_hd__mux2_1
X_7050_ _7074_/S vssd1 vssd1 vccd1 vccd1 _7067_/S sky130_fd_sc_hd__clkbuf_2
X_4262_ _7823_/Q vssd1 vssd1 vccd1 vccd1 _4262_/X sky130_fd_sc_hd__buf_2
XFILLER_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6001_ _7621_/Q _7613_/Q _7605_/Q _7597_/Q _5939_/X _5974_/X vssd1 vssd1 vccd1 vccd1
+ _6001_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4193_ _4193_/A vssd1 vssd1 vccd1 vccd1 _7555_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__2994_ clkbuf_0__2994_/X vssd1 vssd1 vccd1 vccd1 _6167_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6903_ _6943_/A _6939_/A _6897_/X _6904_/C _6916_/B vssd1 vssd1 vccd1 vccd1 _6905_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_50_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3977_ _7641_/Q _3657_/X _3983_/S vssd1 vssd1 vccd1 vccd1 _3978_/A sky130_fd_sc_hd__mux2_1
X_5716_ _5727_/A vssd1 vssd1 vccd1 vccd1 _5725_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_50_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6696_ _6711_/A _6696_/B _6696_/C _6711_/D vssd1 vssd1 vccd1 vccd1 _6696_/Y sky130_fd_sc_hd__nand4_1
X_7893__220 vssd1 vssd1 vccd1 vccd1 _7893__220/HI partID[3] sky130_fd_sc_hd__conb_1
X_5647_ _5647_/A vssd1 vssd1 vccd1 vccd1 _5667_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5578_ _5576_/X _5577_/X _5578_/S vssd1 vssd1 vccd1 vccd1 _5578_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4529_ _4250_/X _7429_/Q _4533_/S vssd1 vssd1 vccd1 vccd1 _4530_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7317_ _7317_/CLK _7317_/D vssd1 vssd1 vccd1 vccd1 _7317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7248_ _7248_/CLK _7248_/D vssd1 vssd1 vccd1 vccd1 _7248_/Q sky130_fd_sc_hd__dfxtp_1
X_6497__66 _6498__67/A vssd1 vssd1 vccd1 vccd1 _7611_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7179_ _7179_/CLK _7179_/D vssd1 vssd1 vccd1 vccd1 _7179_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3127_ clkbuf_0__3127_/X vssd1 vssd1 vccd1 vccd1 _6475_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6733__126 _6733__126/A vssd1 vssd1 vccd1 vccd1 _7692_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 caravel_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3900_ _3900_/A vssd1 vssd1 vccd1 vccd1 _7691_/D sky130_fd_sc_hd__clkbuf_1
X_4880_ _4880_/A vssd1 vssd1 vccd1 vccd1 _7246_/D sky130_fd_sc_hd__clkbuf_1
X_3831_ _7470_/Q vssd1 vssd1 vccd1 vccd1 _4411_/A sky130_fd_sc_hd__buf_2
X_3762_ _3721_/X _7729_/Q _3762_/S vssd1 vssd1 vccd1 vccd1 _3763_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5501_ _7095_/B _6326_/A _5457_/X _5459_/X vssd1 vssd1 vccd1 vccd1 _5501_/X sky130_fd_sc_hd__a31o_1
X_7877__204 vssd1 vssd1 vccd1 vccd1 _7877__204/HI core1Index[4] sky130_fd_sc_hd__conb_1
XFILLER_118_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3693_ _3693_/A vssd1 vssd1 vccd1 vccd1 _7755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6481_ _6481_/A vssd1 vssd1 vccd1 vccd1 _6481_/X sky130_fd_sc_hd__buf_1
X_6278__391 _6281__394/A vssd1 vssd1 vccd1 vccd1 _7444_/CLK sky130_fd_sc_hd__inv_2
X_5432_ _5430_/X _5431_/X _5432_/S vssd1 vssd1 vccd1 vccd1 _5432_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7102_ _7102_/A vssd1 vssd1 vccd1 vccd1 _7854_/D sky130_fd_sc_hd__clkbuf_1
X_4314_ _4314_/A _4314_/B vssd1 vssd1 vccd1 vccd1 _7520_/D sky130_fd_sc_hd__nor2_1
XFILLER_114_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5294_ _5287_/X _7333_/Q _5291_/X _5292_/X _7133_/Q vssd1 vssd1 vccd1 vccd1 _7133_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_99_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4245_ _4242_/X _7538_/Q _4257_/S vssd1 vssd1 vccd1 vccd1 _4246_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4176_ _4243_/A _4614_/D vssd1 vssd1 vccd1 vccd1 _4192_/S sky130_fd_sc_hd__or2_2
XFILLER_28_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6806__8 _6807__9/A vssd1 vssd1 vccd1 vccd1 _7750_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7797_ _7853_/CLK _7797_/D vssd1 vssd1 vccd1 vccd1 _7797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6679_ _6679_/A vssd1 vssd1 vccd1 vccd1 _6679_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6158__362 _6158__362/A vssd1 vssd1 vccd1 vccd1 _7414_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6119__335 _6123__339/A vssd1 vssd1 vccd1 vccd1 _7384_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4030_ _3926_/X _7618_/Q _4038_/S vssd1 vssd1 vccd1 vccd1 _4031_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5981_ _7409_/Q _7350_/Q _7417_/Q _7398_/Q _5979_/X _5980_/X vssd1 vssd1 vccd1 vccd1
+ _5981_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_1_1_0__2762_ clkbuf_0__2762_/X vssd1 vssd1 vccd1 vccd1 _5757__229/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7720_ _7720_/CLK _7720_/D vssd1 vssd1 vccd1 vccd1 _7720_/Q sky130_fd_sc_hd__dfxtp_1
X_4932_ _4932_/A vssd1 vssd1 vccd1 vccd1 _7178_/D sky130_fd_sc_hd__clkbuf_1
X_7651_ _7651_/CLK _7651_/D vssd1 vssd1 vccd1 vccd1 _7651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6602_ _6602_/A _6602_/B _6613_/B vssd1 vssd1 vccd1 vccd1 _6693_/B sky130_fd_sc_hd__nand3_1
XFILLER_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4863_ _4826_/X _7253_/Q _4863_/S vssd1 vssd1 vccd1 vccd1 _4864_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7582_ _7582_/CLK _7582_/D vssd1 vssd1 vccd1 vccd1 _7582_/Q sky130_fd_sc_hd__dfxtp_1
X_4794_ _4794_/A vssd1 vssd1 vccd1 vccd1 _7281_/D sky130_fd_sc_hd__clkbuf_1
X_3814_ _3814_/A vssd1 vssd1 vccd1 vccd1 _7720_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3314_ clkbuf_0__3314_/X vssd1 vssd1 vccd1 vccd1 _6844__39/A sky130_fd_sc_hd__clkbuf_4
X_3745_ _3745_/A vssd1 vssd1 vccd1 vccd1 _3991_/C sky130_fd_sc_hd__clkbuf_2
Xoutput110 _5139_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[25] sky130_fd_sc_hd__buf_2
X_3676_ _7761_/Q _3675_/X _3676_/S vssd1 vssd1 vccd1 vccd1 _3677_/A sky130_fd_sc_hd__mux2_1
X_5415_ _5521_/A vssd1 vssd1 vccd1 vccd1 _5416_/A sky130_fd_sc_hd__clkbuf_4
Xoutput143 _5078_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[29] sky130_fd_sc_hd__buf_2
Xoutput132 _5056_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[19] sky130_fd_sc_hd__buf_2
Xoutput121 _5002_/B vssd1 vssd1 vccd1 vccd1 caravel_wb_cyc_o sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_28_wb_clk_i _7474_/CLK vssd1 vssd1 vccd1 vccd1 _7855_/CLK sky130_fd_sc_hd__clkbuf_16
X_6395_ _6395_/A vssd1 vssd1 vccd1 vccd1 _7529_/D sky130_fd_sc_hd__clkbuf_1
Xoutput154 _5001_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[0] sky130_fd_sc_hd__buf_2
XFILLER_99_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5346_ _7369_/Q _7370_/Q _7371_/Q _7372_/Q _6718_/A _7686_/Q vssd1 vssd1 vccd1 vccd1
+ _5346_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput176 _5219_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[23] sky130_fd_sc_hd__buf_2
XFILLER_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput165 _5186_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[13] sky130_fd_sc_hd__buf_2
Xclkbuf_0__3144_ _6532_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3144_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_102_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5277_ _5270_/X hold1/X _5274_/X _5275_/X _7123_/Q vssd1 vssd1 vccd1 vccd1 _7123_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput187 _5162_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[4] sky130_fd_sc_hd__buf_2
XFILLER_102_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7016_ _7016_/A _7024_/B vssd1 vssd1 vccd1 vccd1 _7017_/A sky130_fd_sc_hd__and2_1
X_4228_ _7543_/Q _4227_/X _4231_/S vssd1 vssd1 vccd1 vccd1 _4229_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4159_ _4158_/X _7568_/Q _4165_/S vssd1 vssd1 vccd1 vccd1 _4160_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7849_ _7853_/CLK _7849_/D vssd1 vssd1 vccd1 vccd1 _7849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6381__456 _6381__456/A vssd1 vssd1 vccd1 vccd1 _7519_/CLK sky130_fd_sc_hd__inv_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6422__486 _6422__486/A vssd1 vssd1 vccd1 vccd1 _7551_/CLK sky130_fd_sc_hd__inv_2
Xinput12 caravel_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 _5201_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput34 caravel_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_2
Xinput23 caravel_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 _5228_/B sky130_fd_sc_hd__clkbuf_1
X_3530_ _7457_/Q _3585_/A vssd1 vssd1 vccd1 vccd1 _4447_/B sky130_fd_sc_hd__and2b_1
Xinput45 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__buf_8
Xclkbuf_1_1__f__3108_ clkbuf_0__3108_/X vssd1 vssd1 vccd1 vccd1 _6379_/A sky130_fd_sc_hd__clkbuf_16
Xinput89 wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 _5892_/A sky130_fd_sc_hd__buf_6
Xinput56 wbs_data_i[11] vssd1 vssd1 vccd1 vccd1 _5038_/A sky130_fd_sc_hd__buf_6
Xinput67 wbs_data_i[21] vssd1 vssd1 vccd1 vccd1 _5060_/A sky130_fd_sc_hd__buf_4
Xinput78 wbs_data_i[31] vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__buf_4
XFILLER_6_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5200_ _5200_/A vssd1 vssd1 vccd1 vccd1 _5200_/X sky130_fd_sc_hd__clkbuf_2
X_6180_ _7798_/Q _7797_/Q _7796_/Q _7795_/Q vssd1 vssd1 vccd1 vccd1 _6228_/B sky130_fd_sc_hd__and4_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5131_ _7339_/Q _5131_/B vssd1 vssd1 vccd1 vccd1 _5132_/A sky130_fd_sc_hd__and2_1
XFILLER_96_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5062_ _5062_/A _5066_/B vssd1 vssd1 vccd1 vccd1 _5063_/A sky130_fd_sc_hd__or2_1
XFILLER_111_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4013_ _4013_/A vssd1 vssd1 vccd1 vccd1 _7626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__2814_ clkbuf_0__2814_/X vssd1 vssd1 vccd1 vccd1 _5916__312/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5964_ _5964_/A vssd1 vssd1 vccd1 vccd1 _5964_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7703_ _7703_/CLK _7703_/D vssd1 vssd1 vccd1 vccd1 _7703_/Q sky130_fd_sc_hd__dfxtp_1
X_5895_ _5895_/A vssd1 vssd1 vccd1 vccd1 _7341_/D sky130_fd_sc_hd__clkbuf_1
X_4915_ _4823_/X _7230_/Q _4917_/S vssd1 vssd1 vccd1 vccd1 _4916_/A sky130_fd_sc_hd__mux2_1
X_7634_ _7634_/CLK _7634_/D vssd1 vssd1 vccd1 vccd1 _7634_/Q sky130_fd_sc_hd__dfxtp_1
X_4846_ _4846_/A vssd1 vssd1 vccd1 vccd1 _7261_/D sky130_fd_sc_hd__clkbuf_1
X_7565_ _7565_/CLK _7565_/D vssd1 vssd1 vccd1 vccd1 _7565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4777_ _4719_/X _7288_/Q _4777_/S vssd1 vssd1 vccd1 vccd1 _4778_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3728_ _3728_/A vssd1 vssd1 vccd1 vccd1 _7744_/D sky130_fd_sc_hd__clkbuf_1
X_5742__216 _5743__217/A vssd1 vssd1 vccd1 vccd1 _7233_/CLK sky130_fd_sc_hd__inv_2
X_7496_ _7496_/CLK _7496_/D vssd1 vssd1 vccd1 vccd1 _7496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3659_ _3659_/A vssd1 vssd1 vccd1 vccd1 _7767_/D sky130_fd_sc_hd__clkbuf_1
X_5329_ _5329_/A vssd1 vssd1 vccd1 vccd1 _7153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__3127_ _6450_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3127_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_102_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5680_ _5680_/A _5682_/A vssd1 vssd1 vccd1 vccd1 _5680_/Y sky130_fd_sc_hd__nor2_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4700_ _4700_/A vssd1 vssd1 vccd1 vccd1 _7319_/D sky130_fd_sc_hd__clkbuf_1
X_4631_ _4631_/A vssd1 vssd1 vccd1 vccd1 _7381_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__2392_ clkbuf_0__2392_/X vssd1 vssd1 vccd1 vccd1 _5252__182/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4562_ _4242_/X _7415_/Q _4570_/S vssd1 vssd1 vccd1 vccd1 _4563_/A sky130_fd_sc_hd__mux2_1
X_7350_ _7350_/CLK _7350_/D vssd1 vssd1 vccd1 vccd1 _7350_/Q sky130_fd_sc_hd__dfxtp_1
X_3513_ _7227_/Q _5679_/B vssd1 vssd1 vccd1 vccd1 _5457_/A sky130_fd_sc_hd__or2_2
X_6301_ _6385_/A vssd1 vssd1 vccd1 vccd1 _6301_/X sky130_fd_sc_hd__buf_1
X_4493_ _4402_/X _7446_/Q _4497_/S vssd1 vssd1 vccd1 vccd1 _4494_/A sky130_fd_sc_hd__mux2_1
X_7281_ _7281_/CLK _7281_/D vssd1 vssd1 vccd1 vccd1 _7281_/Q sky130_fd_sc_hd__dfxtp_1
X_5806__268 _5807__269/A vssd1 vssd1 vccd1 vccd1 _7285_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6232_ _6232_/A vssd1 vssd1 vccd1 vccd1 _6873_/B sky130_fd_sc_hd__clkbuf_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5114_/A _5120_/B vssd1 vssd1 vccd1 vccd1 _5115_/A sky130_fd_sc_hd__and2_1
X_6094_ _7396_/Q _7380_/Q _7650_/Q _7642_/Q _5936_/A _5933_/A vssd1 vssd1 vccd1 vccd1
+ _6095_/B sky130_fd_sc_hd__mux4_2
XFILLER_85_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5045_/A vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__clkbuf_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6996_ _6996_/A vssd1 vssd1 vccd1 vccd1 _6996_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5947_ _5959_/A vssd1 vssd1 vccd1 vccd1 _5947_/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_0_0__3091_ clkbuf_0__3091_/X vssd1 vssd1 vccd1 vccd1 _6306__413/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5878_ _5051_/A _7334_/Q _5884_/S vssd1 vssd1 vccd1 vccd1 _5879_/A sky130_fd_sc_hd__mux2_1
X_7617_ _7617_/CLK _7617_/D vssd1 vssd1 vccd1 vccd1 _7617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4829_ _4937_/A _4829_/B vssd1 vssd1 vccd1 vccd1 _4845_/S sky130_fd_sc_hd__nand2_2
XFILLER_119_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7548_ _7548_/CLK _7548_/D vssd1 vssd1 vccd1 vccd1 _7548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7479_ _7479_/CLK _7479_/D vssd1 vssd1 vccd1 vccd1 _7479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6272__386 _6273__387/A vssd1 vssd1 vccd1 vccd1 _7439_/CLK sky130_fd_sc_hd__inv_2
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_67_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5732_ _5269_/A _5682_/A _5682_/B _5682_/C vssd1 vssd1 vccd1 vccd1 _5735_/B sky130_fd_sc_hd__a2bb2o_1
X_3993_ _3926_/X _7634_/Q _4001_/S vssd1 vssd1 vccd1 vccd1 _3994_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5663_ _5661_/X _5649_/X _5638_/A _7198_/Q _7105_/B vssd1 vssd1 vccd1 vccd1 _5664_/B
+ sky130_fd_sc_hd__a32o_1
X_7402_ _7402_/CLK _7402_/D vssd1 vssd1 vccd1 vccd1 _7402_/Q sky130_fd_sc_hd__dfxtp_1
X_4614_ _4614_/A _4614_/B _4614_/C _4614_/D vssd1 vssd1 vccd1 vccd1 _4630_/S sky130_fd_sc_hd__or4_4
X_5594_ _7243_/Q _7174_/Q _7484_/Q _7251_/Q _4296_/A _4300_/A vssd1 vssd1 vccd1 vccd1
+ _5595_/B sky130_fd_sc_hd__mux4_1
X_7333_ _7333_/CLK _7333_/D vssd1 vssd1 vccd1 vccd1 _7333_/Q sky130_fd_sc_hd__dfxtp_1
X_4545_ _4545_/A vssd1 vssd1 vccd1 vccd1 _7423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4476_ _4476_/A vssd1 vssd1 vccd1 vccd1 _7454_/D sky130_fd_sc_hd__clkbuf_1
X_7264_ _7264_/CLK _7264_/D vssd1 vssd1 vccd1 vccd1 _7264_/Q sky130_fd_sc_hd__dfxtp_1
X_7195_ _7838_/CLK _7195_/D vssd1 vssd1 vccd1 vccd1 _7195_/Q sky130_fd_sc_hd__dfxtp_1
X_6215_ _7796_/Q vssd1 vssd1 vccd1 vccd1 _6918_/A sky130_fd_sc_hd__clkbuf_2
X_6512__79 _6512__79/A vssd1 vssd1 vccd1 vccd1 _7624_/CLK sky130_fd_sc_hd__inv_2
X_6146_ _7406_/Q _5856_/A _6148_/S vssd1 vssd1 vccd1 vccd1 _6147_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5854__306 _5855__307/A vssd1 vssd1 vccd1 vccd1 _7323_/CLK sky130_fd_sc_hd__inv_2
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_25 _5085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_14 _5577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_47 _5036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6077_ _7414_/Q _7355_/Q _7422_/Q _7403_/Q _5956_/X _5942_/X vssd1 vssd1 vccd1 vccd1
+ _6077_/X sky130_fd_sc_hd__mux4_1
XINSDIODE2_36 _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5028_ _5028_/A vssd1 vssd1 vccd1 vccd1 _5028_/X sky130_fd_sc_hd__clkbuf_1
X_6830__28 _6831__29/A vssd1 vssd1 vccd1 vccd1 _7770_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3143_ clkbuf_0__3143_/X vssd1 vssd1 vccd1 vccd1 _6529__92/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6979_ _7812_/Q _7811_/Q vssd1 vssd1 vccd1 vccd1 _6979_/X sky130_fd_sc_hd__or2_1
XFILLER_41_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__2452_ clkbuf_0__2452_/X vssd1 vssd1 vccd1 vccd1 _5385__211/A sky130_fd_sc_hd__clkbuf_16
XFILLER_74_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4330_ _4330_/A vssd1 vssd1 vccd1 vccd1 _7514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4261_ _4261_/A vssd1 vssd1 vccd1 vccd1 _7533_/D sky130_fd_sc_hd__clkbuf_1
X_5918__314 _5918__314/A vssd1 vssd1 vccd1 vccd1 _7355_/CLK sky130_fd_sc_hd__inv_2
X_6000_ _7755_/Q _7747_/Q _7739_/Q _7653_/Q _4465_/A _5937_/X vssd1 vssd1 vccd1 vccd1
+ _6000_/X sky130_fd_sc_hd__mux4_1
X_4192_ _4069_/X _7555_/Q _4192_/S vssd1 vssd1 vccd1 vccd1 _4193_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6902_ _6899_/X _6900_/Y _6902_/S vssd1 vssd1 vccd1 vccd1 _6904_/C sky130_fd_sc_hd__mux2_1
X_6833_ _6845_/A vssd1 vssd1 vccd1 vccd1 _6833_/X sky130_fd_sc_hd__buf_1
XFILLER_63_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3976_ _3976_/A vssd1 vssd1 vccd1 vccd1 _7642_/D sky130_fd_sc_hd__clkbuf_1
X_6764_ _6764_/A vssd1 vssd1 vccd1 vccd1 _6764_/X sky130_fd_sc_hd__buf_1
X_5715_ _5715_/A vssd1 vssd1 vccd1 vccd1 _7218_/D sky130_fd_sc_hd__clkbuf_1
X_6695_ _6679_/X _6684_/X _7678_/Q vssd1 vssd1 vccd1 vccd1 _6695_/X sky130_fd_sc_hd__a21bo_1
XFILLER_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6476__530 _6478__532/A vssd1 vssd1 vccd1 vccd1 _7595_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5646_ _5646_/A vssd1 vssd1 vccd1 vccd1 _7194_/D sky130_fd_sc_hd__clkbuf_1
X_5577_ _7515_/Q _7507_/Q _7446_/Q _7438_/Q _5520_/X _5513_/X vssd1 vssd1 vccd1 vccd1
+ _5577_/X sky130_fd_sc_hd__mux4_2
X_4528_ _4528_/A vssd1 vssd1 vccd1 vccd1 _7430_/D sky130_fd_sc_hd__clkbuf_1
X_7316_ _7316_/CLK _7316_/D vssd1 vssd1 vccd1 vccd1 _7316_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_104_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4459_ _4459_/A _4459_/B vssd1 vssd1 vccd1 vccd1 _7459_/D sky130_fd_sc_hd__nor2_1
X_7247_ _7247_/CLK _7247_/D vssd1 vssd1 vccd1 vccd1 _7247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6765__150 _6768__153/A vssd1 vssd1 vccd1 vccd1 _7717_/CLK sky130_fd_sc_hd__inv_2
X_7178_ _7178_/CLK _7178_/D vssd1 vssd1 vccd1 vccd1 _7178_/Q sky130_fd_sc_hd__dfxtp_1
X_6112__330 _6113__331/A vssd1 vssd1 vccd1 vccd1 _7379_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3126_ clkbuf_0__3126_/X vssd1 vssd1 vccd1 vccd1 _6449__509/A sky130_fd_sc_hd__clkbuf_4
XFILLER_14_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5360__191 _5362__193/A vssd1 vssd1 vccd1 vccd1 _7163_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6345__427 _6347__429/A vssd1 vssd1 vccd1 vccd1 _7490_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3830_ _3830_/A vssd1 vssd1 vccd1 vccd1 _7716_/D sky130_fd_sc_hd__clkbuf_1
X_3761_ _3761_/A vssd1 vssd1 vccd1 vccd1 _7730_/D sky130_fd_sc_hd__clkbuf_1
X_5500_ _7853_/Q vssd1 vssd1 vccd1 vccd1 _7095_/B sky130_fd_sc_hd__buf_2
XFILLER_118_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3692_ _3570_/X _7755_/Q _3696_/S vssd1 vssd1 vccd1 vccd1 _3693_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5431_ _7688_/Q _7277_/Q _7160_/Q _7269_/Q _5426_/X _5427_/X vssd1 vssd1 vccd1 vccd1
+ _5431_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7101_ _7106_/A _7101_/B _7101_/C vssd1 vssd1 vccd1 vccd1 _7102_/A sky130_fd_sc_hd__or3_1
X_4313_ _5613_/A _4316_/A _6308_/B vssd1 vssd1 vccd1 vccd1 _4314_/B sky130_fd_sc_hd__o21ai_1
XFILLER_113_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5293_ _5287_/X _7332_/Q _5291_/X _5292_/X _7132_/Q vssd1 vssd1 vccd1 vccd1 _7132_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_59_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4244_ _4266_/S vssd1 vssd1 vccd1 vccd1 _4257_/S sky130_fd_sc_hd__buf_2
XFILLER_68_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3091_ _6302_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3091_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_101_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4175_ _4175_/A vssd1 vssd1 vccd1 vccd1 _7563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7796_ _7799_/CLK _7796_/D vssd1 vssd1 vccd1 vccd1 _7796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3959_ _3959_/A vssd1 vssd1 vccd1 vccd1 _7649_/D sky130_fd_sc_hd__clkbuf_1
X_6678_ _6675_/X _6677_/X _6665_/X vssd1 vssd1 vccd1 vccd1 _7673_/D sky130_fd_sc_hd__a21oi_1
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5629_ _7191_/Q _7092_/B _5680_/A vssd1 vssd1 vccd1 vccd1 _5629_/X sky130_fd_sc_hd__a21o_1
XFILLER_117_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5791__256 _5792__257/A vssd1 vssd1 vccd1 vccd1 _7273_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3109_ clkbuf_0__3109_/X vssd1 vssd1 vccd1 vccd1 _6359__438/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5980_ _6011_/A vssd1 vssd1 vccd1 vccd1 _5980_/X sky130_fd_sc_hd__buf_2
XFILLER_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2761_ clkbuf_0__2761_/X vssd1 vssd1 vccd1 vccd1 _5749__222/A sky130_fd_sc_hd__clkbuf_4
X_4931_ _4233_/X _7178_/Q _4935_/S vssd1 vssd1 vccd1 vccd1 _4932_/A sky130_fd_sc_hd__mux2_1
X_7650_ _7650_/CLK _7650_/D vssd1 vssd1 vccd1 vccd1 _7650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4862_ _4862_/A vssd1 vssd1 vccd1 vccd1 _7254_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6601_ _5584_/X _6686_/B _6682_/B _5565_/X _6600_/X vssd1 vssd1 vccd1 vccd1 _6601_/Y
+ sky130_fd_sc_hd__a221oi_4
X_3813_ _3784_/X _7720_/Q _3829_/S vssd1 vssd1 vccd1 vccd1 _3814_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3313_ clkbuf_0__3313_/X vssd1 vssd1 vccd1 vccd1 _6836__32/A sky130_fd_sc_hd__clkbuf_4
X_4793_ _4716_/X _7281_/Q _4795_/S vssd1 vssd1 vccd1 vccd1 _4794_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7581_ _7581_/CLK _7581_/D vssd1 vssd1 vccd1 vccd1 _7581_/Q sky130_fd_sc_hd__dfxtp_1
X_6532_ _6538_/A vssd1 vssd1 vccd1 vccd1 _6532_/X sky130_fd_sc_hd__buf_1
X_3744_ _4009_/B vssd1 vssd1 vccd1 vccd1 _4424_/A sky130_fd_sc_hd__clkbuf_2
X_3675_ _7822_/Q vssd1 vssd1 vccd1 vccd1 _3675_/X sky130_fd_sc_hd__clkbuf_4
X_6463_ _6475_/A vssd1 vssd1 vccd1 vccd1 _6463_/X sky130_fd_sc_hd__buf_1
Xoutput100 _5119_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[16] sky130_fd_sc_hd__buf_2
XFILLER_118_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5414_ _7519_/Q vssd1 vssd1 vccd1 vccd1 _5521_/A sky130_fd_sc_hd__clkbuf_4
Xoutput111 _5141_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[26] sky130_fd_sc_hd__buf_2
Xoutput133 _5017_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[1] sky130_fd_sc_hd__buf_2
Xoutput122 _5014_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[0] sky130_fd_sc_hd__buf_2
X_6394_ _6394_/A _7432_/Q _6394_/C vssd1 vssd1 vccd1 vccd1 _6395_/A sky130_fd_sc_hd__and3_1
Xoutput144 _5019_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[2] sky130_fd_sc_hd__buf_2
Xoutput155 _5003_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[1] sky130_fd_sc_hd__buf_2
X_5345_ _7685_/Q vssd1 vssd1 vccd1 vccd1 _6718_/A sky130_fd_sc_hd__clkbuf_2
Xoutput177 _5221_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[24] sky130_fd_sc_hd__buf_2
Xoutput166 _5190_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[14] sky130_fd_sc_hd__buf_2
X_5367__197 _5368__198/A vssd1 vssd1 vccd1 vccd1 _7169_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3143_ _6526_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3143_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5276_ _5270_/X _7154_/Q _5274_/X _5275_/X _7122_/Q vssd1 vssd1 vccd1 vccd1 _7122_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_87_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput188 _5166_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_101_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7015_ _7030_/B vssd1 vssd1 vccd1 vccd1 _7024_/B sky130_fd_sc_hd__clkbuf_2
X_4227_ _7472_/Q vssd1 vssd1 vccd1 vccd1 _4227_/X sky130_fd_sc_hd__buf_4
XFILLER_56_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4158_ _4402_/A vssd1 vssd1 vccd1 vccd1 _4158_/X sky130_fd_sc_hd__buf_2
X_4089_ _4089_/A vssd1 vssd1 vccd1 vccd1 _7595_/D sky130_fd_sc_hd__clkbuf_1
X_7034__53 _7035__54/A vssd1 vssd1 vccd1 vccd1 _7832_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7848_ _7854_/CLK _7848_/D vssd1 vssd1 vccd1 vccd1 _7848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7779_ _7779_/CLK _7779_/D vssd1 vssd1 vccd1 vccd1 _7779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6848__42 _6848__42/A vssd1 vssd1 vccd1 vccd1 _7784_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6778__160 _6779__161/A vssd1 vssd1 vccd1 vccd1 _7727_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6125__340 _6127__342/A vssd1 vssd1 vccd1 vccd1 _7389_/CLK sky130_fd_sc_hd__inv_2
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 caravel_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 _5207_/B sky130_fd_sc_hd__clkbuf_1
Xinput24 caravel_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 _5230_/B sky130_fd_sc_hd__clkbuf_1
Xinput35 caravel_wb_error_i vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
Xinput46 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__buf_8
XFILLER_6_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput79 wbs_data_i[3] vssd1 vssd1 vccd1 vccd1 _3587_/A sky130_fd_sc_hd__clkbuf_4
Xinput57 wbs_data_i[12] vssd1 vssd1 vccd1 vccd1 _5040_/A sky130_fd_sc_hd__buf_6
Xinput68 wbs_data_i[22] vssd1 vssd1 vccd1 vccd1 _5062_/A sky130_fd_sc_hd__buf_4
X_5130_ _5130_/A vssd1 vssd1 vccd1 vccd1 _5130_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5061_ _5061_/A vssd1 vssd1 vccd1 vccd1 _5061_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4012_ _3926_/X _7626_/Q _4020_/S vssd1 vssd1 vccd1 vccd1 _4013_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__2813_ clkbuf_0__2813_/X vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5963_ _6016_/A _5963_/B vssd1 vssd1 vccd1 vccd1 _5963_/X sky130_fd_sc_hd__or2_1
XFILLER_65_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7702_ _7702_/CLK _7702_/D vssd1 vssd1 vccd1 vccd1 _7702_/Q sky130_fd_sc_hd__dfxtp_1
X_4914_ _4914_/A vssd1 vssd1 vccd1 vccd1 _7231_/D sky130_fd_sc_hd__clkbuf_1
X_5894_ _7341_/Q _5066_/A _5902_/S vssd1 vssd1 vccd1 vccd1 _5895_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7633_ _7633_/CLK _7633_/D vssd1 vssd1 vccd1 vccd1 _7633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4845_ _4826_/X _7261_/Q _4845_/S vssd1 vssd1 vccd1 vccd1 _4846_/A sky130_fd_sc_hd__mux2_1
X_4776_ _4776_/A vssd1 vssd1 vccd1 vccd1 _7289_/D sky130_fd_sc_hd__clkbuf_1
X_7564_ _7564_/CLK _7564_/D vssd1 vssd1 vccd1 vccd1 _7564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3727_ _3698_/X _7744_/Q _3735_/S vssd1 vssd1 vccd1 vccd1 _3728_/A sky130_fd_sc_hd__mux2_1
X_6358__437 _6359__438/A vssd1 vssd1 vccd1 vccd1 _7500_/CLK sky130_fd_sc_hd__inv_2
X_7495_ _7495_/CLK _7495_/D vssd1 vssd1 vccd1 vccd1 _7495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3658_ _7767_/Q _3657_/X _3667_/S vssd1 vssd1 vccd1 vccd1 _3659_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3589_ _3589_/A vssd1 vssd1 vccd1 vccd1 _5239_/A sky130_fd_sc_hd__clkbuf_2
X_5328_ _7024_/A _7153_/Q _5328_/S vssd1 vssd1 vccd1 vccd1 _5329_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3089_ clkbuf_0__3089_/X vssd1 vssd1 vccd1 vccd1 _6385_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3126_ _6444_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3126_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_28_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4630_ _3675_/X _7381_/Q _4630_/S vssd1 vssd1 vccd1 vccd1 _4631_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__2391_ clkbuf_0__2391_/X vssd1 vssd1 vccd1 vccd1 _5249_/A sky130_fd_sc_hd__clkbuf_4
X_5253__183 _5254__184/A vssd1 vssd1 vccd1 vccd1 _7112_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4561_ _4576_/S vssd1 vssd1 vccd1 vccd1 _4570_/S sky130_fd_sc_hd__buf_2
X_6300_ _6300_/A vssd1 vssd1 vccd1 vccd1 _6300_/X sky130_fd_sc_hd__buf_1
X_3512_ _7226_/Q vssd1 vssd1 vccd1 vccd1 _5679_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6470__525 _6471__526/A vssd1 vssd1 vccd1 vccd1 _7590_/CLK sky130_fd_sc_hd__inv_2
X_7280_ _7280_/CLK _7280_/D vssd1 vssd1 vccd1 vccd1 _7280_/Q sky130_fd_sc_hd__dfxtp_1
X_4492_ _4492_/A vssd1 vssd1 vccd1 vccd1 _7447_/D sky130_fd_sc_hd__clkbuf_1
X_6231_ _6231_/A _6231_/B vssd1 vssd1 vccd1 vccd1 _6232_/A sky130_fd_sc_hd__nand2_1
X_6524__88 _6524__88/A vssd1 vssd1 vccd1 vccd1 _7633_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5113_/A vssd1 vssd1 vccd1 vccd1 _5113_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6093_ _7415_/Q _7356_/Q _7423_/Q _7404_/Q _5956_/X _5942_/X vssd1 vssd1 vccd1 vccd1
+ _6093_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5044_/A _5044_/B vssd1 vssd1 vccd1 vccd1 _5045_/A sky130_fd_sc_hd__or2_1
XFILLER_84_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6842__37 _6842__37/A vssd1 vssd1 vccd1 vccd1 _7779_/CLK sky130_fd_sc_hd__inv_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6995_ _7013_/S vssd1 vssd1 vccd1 vccd1 _6995_/X sky130_fd_sc_hd__clkbuf_2
X_5946_ _7461_/Q vssd1 vssd1 vccd1 vccd1 _5959_/A sky130_fd_sc_hd__clkinv_2
Xclkbuf_1_0_0__3090_ clkbuf_0__3090_/X vssd1 vssd1 vccd1 vccd1 _6348_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5877_ _5877_/A vssd1 vssd1 vccd1 vccd1 _7333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7616_ _7616_/CLK _7616_/D vssd1 vssd1 vccd1 vccd1 _7616_/Q sky130_fd_sc_hd__dfxtp_1
X_4828_ _4828_/A vssd1 vssd1 vccd1 vccd1 _7269_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4759_ _4719_/X _7296_/Q _4759_/S vssd1 vssd1 vccd1 vccd1 _4760_/A sky130_fd_sc_hd__mux2_1
X_7547_ _7547_/CLK _7547_/D vssd1 vssd1 vccd1 vccd1 _7547_/Q sky130_fd_sc_hd__dfxtp_1
X_7478_ _7478_/CLK _7478_/D vssd1 vssd1 vccd1 vccd1 _7478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_12_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7331_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3109_ _6355_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3109_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3992_ _4007_/S vssd1 vssd1 vccd1 vccd1 _4001_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5731_ _5731_/A vssd1 vssd1 vccd1 vccd1 _7225_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5812__273 _5812__273/A vssd1 vssd1 vccd1 vccd1 _7290_/CLK sky130_fd_sc_hd__inv_2
X_5662_ _5662_/A vssd1 vssd1 vccd1 vccd1 _7105_/B sky130_fd_sc_hd__clkbuf_2
X_7401_ _7401_/CLK _7401_/D vssd1 vssd1 vccd1 vccd1 _7401_/Q sky130_fd_sc_hd__dfxtp_1
X_4613_ _4613_/A vssd1 vssd1 vccd1 vccd1 _7389_/D sky130_fd_sc_hd__clkbuf_1
X_5593_ _5586_/X _5588_/X _5590_/X _5592_/X vssd1 vssd1 vccd1 vccd1 _5593_/X sky130_fd_sc_hd__o22a_1
X_4544_ _4242_/X _7423_/Q _4552_/S vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__mux2_1
X_7332_ _7336_/CLK _7332_/D vssd1 vssd1 vccd1 vccd1 _7332_/Q sky130_fd_sc_hd__dfxtp_1
X_7263_ _7263_/CLK _7263_/D vssd1 vssd1 vccd1 vccd1 _7263_/Q sky130_fd_sc_hd__dfxtp_1
X_6214_ _7850_/Q _6884_/A _6884_/B vssd1 vssd1 vccd1 vccd1 _6214_/X sky130_fd_sc_hd__and3_1
X_6435__497 _6435__497/A vssd1 vssd1 vccd1 vccd1 _7562_/CLK sky130_fd_sc_hd__inv_2
X_4475_ _4402_/X _7454_/Q _4479_/S vssd1 vssd1 vccd1 vccd1 _4476_/A sky130_fd_sc_hd__mux2_1
X_7194_ _7329_/CLK _7194_/D vssd1 vssd1 vccd1 vccd1 _7194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6145_ _6145_/A vssd1 vssd1 vccd1 vccd1 _7405_/D sky130_fd_sc_hd__clkbuf_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6815__15 _6818__18/A vssd1 vssd1 vccd1 vccd1 _7757_/CLK sky130_fd_sc_hd__inv_2
X_6076_ _6072_/X _6073_/X _6074_/X _6075_/X _5953_/X _4436_/X vssd1 vssd1 vccd1 vccd1
+ _6076_/X sky130_fd_sc_hd__mux4_2
XINSDIODE2_15 _5190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _7028_/A _5033_/B vssd1 vssd1 vccd1 vccd1 _5028_/A sky130_fd_sc_hd__or2_1
XINSDIODE2_48 _7340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_37 _7030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_26 _5085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3142_ clkbuf_0__3142_/X vssd1 vssd1 vccd1 vccd1 _6524__88/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6978_ _6978_/A vssd1 vssd1 vccd1 vccd1 _6996_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6152__358 _6152__358/A vssd1 vssd1 vccd1 vccd1 _7410_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5755__227 _5755__227/A vssd1 vssd1 vccd1 vccd1 _7244_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7868__195 vssd1 vssd1 vccd1 vccd1 _7868__195/HI core0Index[2] sky130_fd_sc_hd__conb_1
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4260_ _4259_/X _7533_/Q _4266_/S vssd1 vssd1 vccd1 vccd1 _4261_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4191_ _4191_/A vssd1 vssd1 vccd1 vccd1 _7556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6901_ _6901_/A input1/X vssd1 vssd1 vccd1 vccd1 _6902_/S sky130_fd_sc_hd__nor2_1
X_6832_ _6832_/A vssd1 vssd1 vccd1 vccd1 _6832_/X sky130_fd_sc_hd__buf_1
XFILLER_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3975_ _7642_/Q _3649_/X _3983_/S vssd1 vssd1 vccd1 vccd1 _3976_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5714_ _7218_/Q _7333_/Q _5714_/S vssd1 vssd1 vccd1 vccd1 _5715_/A sky130_fd_sc_hd__mux2_1
X_6694_ _6692_/Y _6693_/X _5970_/X vssd1 vssd1 vccd1 vccd1 _7677_/D sky130_fd_sc_hd__o21a_1
XFILLER_50_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5645_ _5645_/A _5645_/B vssd1 vssd1 vccd1 vccd1 _5646_/A sky130_fd_sc_hd__or2_1
XFILLER_31_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5576_ _7242_/Q _7173_/Q _7483_/Q _7250_/Q _5479_/X _5518_/X vssd1 vssd1 vccd1 vccd1
+ _5576_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4527_ _4247_/X _7430_/Q _4533_/S vssd1 vssd1 vccd1 vccd1 _4528_/A sky130_fd_sc_hd__mux2_1
X_7315_ _7315_/CLK _7315_/D vssd1 vssd1 vccd1 vccd1 _7315_/Q sky130_fd_sc_hd__dfxtp_2
X_4458_ _4451_/A _4461_/A _4421_/X vssd1 vssd1 vccd1 vccd1 _4459_/B sky130_fd_sc_hd__o21ai_1
XFILLER_49_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7246_ _7246_/CLK _7246_/D vssd1 vssd1 vccd1 vccd1 _7246_/Q sky130_fd_sc_hd__dfxtp_1
X_7177_ _7177_/CLK _7177_/D vssd1 vssd1 vccd1 vccd1 _7177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4389_ _7487_/Q _3947_/A _4391_/S vssd1 vssd1 vccd1 vccd1 _4390_/A sky130_fd_sc_hd__mux2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _7576_/Q _7386_/Q _7734_/Q _7632_/Q _6002_/X _4465_/X vssd1 vssd1 vccd1 vccd1
+ _6059_/X sky130_fd_sc_hd__mux4_1
X_5819__279 _5819__279/A vssd1 vssd1 vccd1 vccd1 _7296_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3125_ clkbuf_0__3125_/X vssd1 vssd1 vccd1 vccd1 _6442__503/A sky130_fd_sc_hd__clkbuf_4
X_7902__229 vssd1 vssd1 vccd1 vccd1 _7902__229/HI versionID[3] sky130_fd_sc_hd__conb_1
XFILLER_14_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7038__3 _7039__4/A vssd1 vssd1 vccd1 vccd1 _7836_/CLK sky130_fd_sc_hd__inv_2
X_6772__155 _6773__156/A vssd1 vssd1 vccd1 vccd1 _7722_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3760_ _3718_/X _7730_/Q _3762_/S vssd1 vssd1 vccd1 vccd1 _3761_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3691_ _3691_/A vssd1 vssd1 vccd1 vccd1 _7756_/D sky130_fd_sc_hd__clkbuf_1
X_5430_ _7293_/Q _7285_/Q _7261_/Q _7109_/Q _5413_/X _5416_/X vssd1 vssd1 vccd1 vccd1
+ _5430_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5292_ _5308_/A vssd1 vssd1 vccd1 vccd1 _5292_/X sky130_fd_sc_hd__clkbuf_2
X_7100_ _7100_/A _7105_/B _7100_/C vssd1 vssd1 vccd1 vccd1 _7101_/C sky130_fd_sc_hd__and3_1
X_4312_ _4312_/A _4312_/B vssd1 vssd1 vccd1 vccd1 _4316_/A sky130_fd_sc_hd__and2_1
X_7031_ _7031_/A vssd1 vssd1 vccd1 vccd1 _7829_/D sky130_fd_sc_hd__clkbuf_1
X_4243_ _4243_/A _4243_/B vssd1 vssd1 vccd1 vccd1 _4266_/S sky130_fd_sc_hd__or2_2
XFILLER_101_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3090_ _6301_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3090_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_67_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4174_ _4173_/X _7563_/Q _4174_/S vssd1 vssd1 vccd1 vccd1 _4175_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6285__397 _6287__399/A vssd1 vssd1 vccd1 vccd1 _7450_/CLK sky130_fd_sc_hd__inv_2
X_7795_ _7799_/CLK _7795_/D vssd1 vssd1 vccd1 vccd1 _7795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6746_ _6746_/A vssd1 vssd1 vccd1 vccd1 _6746_/X sky130_fd_sc_hd__buf_1
X_3958_ _3932_/X _7649_/Q _3964_/S vssd1 vssd1 vccd1 vccd1 _3959_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6677_ _6677_/A _6677_/B _6702_/C vssd1 vssd1 vccd1 vccd1 _6677_/X sky130_fd_sc_hd__or3_1
X_3889_ _4919_/B _4955_/B vssd1 vssd1 vccd1 vccd1 _3905_/S sky130_fd_sc_hd__or2_2
X_5628_ _6872_/A _5394_/Y _5448_/X _5627_/X vssd1 vssd1 vccd1 vccd1 _5628_/X sky130_fd_sc_hd__a22o_1
X_5559_ _5557_/X _5558_/X _5578_/S vssd1 vssd1 vccd1 vccd1 _5559_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7229_ _7229_/CLK _7229_/D vssd1 vssd1 vccd1 vccd1 _7229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6305__412 _6307__414/A vssd1 vssd1 vccd1 vccd1 _7465_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6351__432 _6353__434/A vssd1 vssd1 vccd1 vccd1 _7495_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2760_ clkbuf_0__2760_/X vssd1 vssd1 vccd1 vccd1 _5745__219/A sky130_fd_sc_hd__clkbuf_4
X_7883__210 vssd1 vssd1 vccd1 vccd1 _7883__210/HI manufacturerID[2] sky130_fd_sc_hd__conb_1
X_4930_ _4930_/A vssd1 vssd1 vccd1 vccd1 _7179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6165__368 _6166__369/A vssd1 vssd1 vccd1 vccd1 _7420_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4861_ _4823_/X _7254_/Q _4863_/S vssd1 vssd1 vccd1 vccd1 _4862_/A sky130_fd_sc_hd__mux2_1
X_6600_ _7852_/Q _6600_/B vssd1 vssd1 vccd1 vccd1 _6600_/X sky130_fd_sc_hd__xor2_1
XFILLER_60_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3812_ _3841_/S vssd1 vssd1 vccd1 vccd1 _3829_/S sky130_fd_sc_hd__buf_2
X_5768__237 _5769__238/A vssd1 vssd1 vccd1 vccd1 _7254_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3312_ clkbuf_0__3312_/X vssd1 vssd1 vccd1 vccd1 _6845_/A sky130_fd_sc_hd__clkbuf_4
X_4792_ _4792_/A vssd1 vssd1 vccd1 vccd1 _7282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7580_ _7580_/CLK _7580_/D vssd1 vssd1 vccd1 vccd1 _7580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3743_ _4009_/A vssd1 vssd1 vccd1 vccd1 _4131_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3674_ _3674_/A vssd1 vssd1 vccd1 vccd1 _7762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput101 _5121_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[17] sky130_fd_sc_hd__buf_2
XFILLER_118_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5413_ _5427_/A vssd1 vssd1 vccd1 vccd1 _5413_/X sky130_fd_sc_hd__buf_4
Xoutput112 _5143_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[27] sky130_fd_sc_hd__buf_2
Xoutput134 _5059_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[20] sky130_fd_sc_hd__buf_2
Xoutput123 _5037_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[10] sky130_fd_sc_hd__buf_2
X_5344_ _7660_/Q vssd1 vssd1 vccd1 vccd1 _6725_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput145 _5080_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[30] sky130_fd_sc_hd__buf_2
Xoutput156 _5007_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[2] sky130_fd_sc_hd__buf_2
XFILLER_114_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput167 _5193_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[15] sky130_fd_sc_hd__buf_2
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5275_ _5284_/A vssd1 vssd1 vccd1 vccd1 _5275_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3142_ _6520_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3142_/X sky130_fd_sc_hd__clkbuf_16
Xoutput189 _5168_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[6] sky130_fd_sc_hd__buf_2
Xoutput178 _5223_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[25] sky130_fd_sc_hd__buf_2
XFILLER_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4226_ _4226_/A vssd1 vssd1 vccd1 vccd1 _7544_/D sky130_fd_sc_hd__clkbuf_1
X_7014_ _7014_/A _7014_/B vssd1 vssd1 vccd1 vccd1 _7821_/D sky130_fd_sc_hd__nor2_1
X_4157_ _4157_/A vssd1 vssd1 vccd1 vccd1 _7569_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4088_ _4069_/X _7595_/Q _4088_/S vssd1 vssd1 vccd1 vccd1 _4089_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_37_wb_clk_i clkbuf_opt_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7473_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7847_ _7855_/CLK _7847_/D vssd1 vssd1 vccd1 vccd1 _7847_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7778_ _7778_/CLK _7778_/D vssd1 vssd1 vccd1 vccd1 _7778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput25 caravel_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_2
Xinput14 caravel_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_4
Xinput36 wb_rst_i vssd1 vssd1 vccd1 vccd1 _3589_/A sky130_fd_sc_hd__buf_4
XFILLER_116_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput47 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _5092_/A sky130_fd_sc_hd__buf_6
Xinput69 wbs_data_i[23] vssd1 vssd1 vccd1 vccd1 _5064_/A sky130_fd_sc_hd__buf_4
Xinput58 wbs_data_i[13] vssd1 vssd1 vccd1 vccd1 _5042_/A sky130_fd_sc_hd__buf_6
XFILLER_6_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5060_ _5060_/A _5066_/B vssd1 vssd1 vccd1 vccd1 _5061_/A sky130_fd_sc_hd__or2_1
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4011_ _4026_/S vssd1 vssd1 vccd1 vccd1 _4020_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_65_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6642__114 _6642__114/A vssd1 vssd1 vccd1 vccd1 _7661_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5962_ _7389_/Q _7373_/Q _7643_/Q _7635_/Q _6002_/A _5956_/X vssd1 vssd1 vccd1 vccd1
+ _5963_/B sky130_fd_sc_hd__mux4_1
XFILLER_65_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7701_ _7701_/CLK _7701_/D vssd1 vssd1 vccd1 vccd1 _7701_/Q sky130_fd_sc_hd__dfxtp_1
X_4913_ _4820_/X _7231_/Q _4917_/S vssd1 vssd1 vccd1 vccd1 _4914_/A sky130_fd_sc_hd__mux2_1
X_5893_ _5908_/S vssd1 vssd1 vccd1 vccd1 _5902_/S sky130_fd_sc_hd__clkbuf_2
X_7632_ _7632_/CLK _7632_/D vssd1 vssd1 vccd1 vccd1 _7632_/Q sky130_fd_sc_hd__dfxtp_1
X_4844_ _4844_/A vssd1 vssd1 vccd1 vccd1 _7262_/D sky130_fd_sc_hd__clkbuf_1
X_4775_ _4716_/X _7289_/Q _4777_/S vssd1 vssd1 vccd1 vccd1 _4776_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7563_ _7563_/CLK _7563_/D vssd1 vssd1 vccd1 vccd1 _7563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3726_ _3741_/S vssd1 vssd1 vccd1 vccd1 _3735_/S sky130_fd_sc_hd__buf_2
X_6514_ _6520_/A vssd1 vssd1 vccd1 vccd1 _6514_/X sky130_fd_sc_hd__buf_1
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7494_ _7494_/CLK _7494_/D vssd1 vssd1 vccd1 vccd1 _7494_/Q sky130_fd_sc_hd__dfxtp_1
X_3657_ _7828_/Q vssd1 vssd1 vccd1 vccd1 _3657_/X sky130_fd_sc_hd__buf_4
X_3588_ _3588_/A vssd1 vssd1 vccd1 vccd1 _3588_/X sky130_fd_sc_hd__clkbuf_4
X_5327_ _5327_/A vssd1 vssd1 vccd1 vccd1 _7152_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3088_ clkbuf_0__3088_/X vssd1 vssd1 vccd1 vccd1 _6299__409/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3125_ _6438_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3125_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5189_ _7198_/Q _5189_/B _5198_/A vssd1 vssd1 vccd1 vccd1 _5189_/X sky130_fd_sc_hd__and3_1
X_4209_ _4170_/X _7548_/Q _4211_/S vssd1 vssd1 vccd1 vccd1 _4210_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5838__293 _5838__293/A vssd1 vssd1 vccd1 vccd1 _7310_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__2390_ clkbuf_0__2390_/X vssd1 vssd1 vccd1 vccd1 _5795_/A sky130_fd_sc_hd__clkbuf_4
X_4560_ _4596_/A _4668_/B vssd1 vssd1 vccd1 vccd1 _4576_/S sky130_fd_sc_hd__nand2_2
XFILLER_8_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3511_ _7206_/Q _7207_/Q _5435_/B vssd1 vssd1 vccd1 vccd1 _5388_/A sky130_fd_sc_hd__or3_1
X_4491_ _4399_/X _7447_/Q _4497_/S vssd1 vssd1 vccd1 vccd1 _4492_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6230_ _6213_/Y _6214_/X _6225_/X _6991_/C _6229_/X vssd1 vssd1 vccd1 vccd1 _6238_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_6_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6161_ _6167_/A vssd1 vssd1 vccd1 vccd1 _6161_/X sky130_fd_sc_hd__buf_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5112_/A _5120_/B vssd1 vssd1 vccd1 vccd1 _5113_/A sky130_fd_sc_hd__and2_1
XFILLER_69_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6092_ _6088_/X _6089_/X _6090_/X _6091_/X _5953_/X _5947_/X vssd1 vssd1 vccd1 vccd1
+ _6092_/X sky130_fd_sc_hd__mux4_2
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5043_/A vssd1 vssd1 vccd1 vccd1 _5043_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6364__442 _6366__444/A vssd1 vssd1 vccd1 vccd1 _7505_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6994_ _6996_/A _6994_/B vssd1 vssd1 vccd1 vccd1 _7013_/S sky130_fd_sc_hd__nand2_1
X_5945_ _6095_/A vssd1 vssd1 vccd1 vccd1 _5945_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_40_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5876_ _5049_/A _7333_/Q _5884_/S vssd1 vssd1 vccd1 vccd1 _5877_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7615_ _7615_/CLK _7615_/D vssd1 vssd1 vccd1 vccd1 _7615_/Q sky130_fd_sc_hd__dfxtp_1
X_4827_ _4826_/X _7269_/Q _4827_/S vssd1 vssd1 vccd1 vccd1 _4828_/A sky130_fd_sc_hd__mux2_1
X_4758_ _4758_/A vssd1 vssd1 vccd1 vccd1 _7297_/D sky130_fd_sc_hd__clkbuf_1
X_7546_ _7546_/CLK _7546_/D vssd1 vssd1 vccd1 vccd1 _7546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3709_ _3938_/A vssd1 vssd1 vccd1 vccd1 _3709_/X sky130_fd_sc_hd__clkbuf_2
X_7477_ _7477_/CLK _7477_/D vssd1 vssd1 vccd1 vccd1 _7477_/Q sky130_fd_sc_hd__dfxtp_1
X_4689_ _4393_/X _7324_/Q _4697_/S vssd1 vssd1 vccd1 vccd1 _4690_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3108_ _6354_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3108_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3991_ _4131_/A _4424_/A _3991_/C _4243_/B vssd1 vssd1 vccd1 vccd1 _4007_/S sky130_fd_sc_hd__or4_4
X_5730_ _7225_/Q _7340_/Q _6148_/S vssd1 vssd1 vccd1 vccd1 _5731_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7400_ _7400_/CLK _7400_/D vssd1 vssd1 vccd1 vccd1 _7400_/Q sky130_fd_sc_hd__dfxtp_1
X_5661_ _7841_/Q vssd1 vssd1 vccd1 vccd1 _5661_/X sky130_fd_sc_hd__buf_2
X_4612_ _4265_/X _7389_/Q _4612_/S vssd1 vssd1 vccd1 vccd1 _4613_/A sky130_fd_sc_hd__mux2_1
X_5592_ _5432_/S _5591_/X _5404_/X vssd1 vssd1 vccd1 vccd1 _5592_/X sky130_fd_sc_hd__a21o_1
XFILLER_116_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4543_ _4558_/S vssd1 vssd1 vccd1 vccd1 _4552_/S sky130_fd_sc_hd__buf_2
X_7331_ _7331_/CLK _7331_/D vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XFILLER_116_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7262_ _7262_/CLK _7262_/D vssd1 vssd1 vccd1 vccd1 _7262_/Q sky130_fd_sc_hd__dfxtp_1
X_6213_ _6884_/A _6884_/B _5565_/X vssd1 vssd1 vccd1 vccd1 _6213_/Y sky130_fd_sc_hd__a21oi_2
X_4474_ _4474_/A vssd1 vssd1 vccd1 vccd1 _7455_/D sky130_fd_sc_hd__clkbuf_1
X_6138__351 _6138__351/A vssd1 vssd1 vccd1 vccd1 _7400_/CLK sky130_fd_sc_hd__inv_2
X_7193_ _7329_/CLK _7193_/D vssd1 vssd1 vccd1 vccd1 _7193_/Q sky130_fd_sc_hd__dfxtp_1
X_6144_ _6326_/A _5318_/A _6148_/S vssd1 vssd1 vccd1 vccd1 _6145_/A sky130_fd_sc_hd__mux2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6075_ _7759_/Q _7751_/Q _7743_/Q _7657_/Q _5939_/X _5940_/X vssd1 vssd1 vccd1 vccd1
+ _6075_/X sky130_fd_sc_hd__mux4_1
XINSDIODE2_16 _5210_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_49 _7100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5026_ _5026_/A vssd1 vssd1 vccd1 vccd1 _5026_/X sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_38 _5031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_27 _5085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3141_ clkbuf_0__3141_/X vssd1 vssd1 vccd1 vccd1 _6516__81/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6977_ _7811_/Q _6974_/Y _6976_/X _6909_/X vssd1 vssd1 vccd1 vccd1 _7811_/D sky130_fd_sc_hd__o211a_1
XFILLER_41_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5859_ _5859_/A vssd1 vssd1 vccd1 vccd1 _7325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7529_ _7799_/CLK _7529_/D vssd1 vssd1 vccd1 vccd1 _7529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4190_ _4066_/X _7556_/Q _4192_/S vssd1 vssd1 vccd1 vccd1 _4191_/A sky130_fd_sc_hd__mux2_1
X_6502__70 _6504__72/A vssd1 vssd1 vccd1 vccd1 _7615_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6900_ _6916_/A _6900_/B vssd1 vssd1 vccd1 vccd1 _6900_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5372__201 _5374__203/A vssd1 vssd1 vccd1 vccd1 _7173_/CLK sky130_fd_sc_hd__inv_2
X_3974_ _3989_/S vssd1 vssd1 vccd1 vccd1 _3983_/S sky130_fd_sc_hd__buf_2
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5713_ _5713_/A vssd1 vssd1 vccd1 vccd1 _7217_/D sky130_fd_sc_hd__clkbuf_1
X_6693_ _6711_/A _6693_/B _6693_/C _6711_/D vssd1 vssd1 vccd1 vccd1 _6693_/X sky130_fd_sc_hd__and4_1
XFILLER_31_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5644_ _6249_/A _5672_/D _5638_/X _7194_/Q _5639_/X vssd1 vssd1 vccd1 vccd1 _5645_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_117_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7314_ _7314_/CLK _7314_/D vssd1 vssd1 vccd1 vccd1 _7314_/Q sky130_fd_sc_hd__dfxtp_2
X_5575_ _5573_/X _5574_/X _5575_/S vssd1 vssd1 vccd1 vccd1 _5575_/X sky130_fd_sc_hd__mux2_1
X_4526_ _4526_/A vssd1 vssd1 vccd1 vccd1 _7431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4457_ _4457_/A _4457_/B vssd1 vssd1 vccd1 vccd1 _4461_/A sky130_fd_sc_hd__and2_1
XFILLER_49_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7245_ _7245_/CLK _7245_/D vssd1 vssd1 vccd1 vccd1 _7245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7176_ _7176_/CLK _7176_/D vssd1 vssd1 vccd1 vccd1 _7176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4388_ _4388_/A vssd1 vssd1 vccd1 vccd1 _7488_/D sky130_fd_sc_hd__clkbuf_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6058_ _7624_/Q _7616_/Q _7608_/Q _7600_/Q _5935_/X _5974_/X vssd1 vssd1 vccd1 vccd1
+ _6058_/X sky130_fd_sc_hd__mux4_2
XFILLER_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5009_ _5009_/A vssd1 vssd1 vccd1 vccd1 _5009_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3124_ clkbuf_0__3124_/X vssd1 vssd1 vccd1 vccd1 _6437__499/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5761__232 _5762__233/A vssd1 vssd1 vccd1 vccd1 _7249_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3690_ _3566_/X _7756_/Q _3690_/S vssd1 vssd1 vccd1 vccd1 _3691_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5291_ _5307_/A vssd1 vssd1 vccd1 vccd1 _5291_/X sky130_fd_sc_hd__clkbuf_2
X_4311_ _5433_/S _4314_/A _4310_/Y vssd1 vssd1 vccd1 vccd1 _7521_/D sky130_fd_sc_hd__o21a_1
X_4242_ _7829_/Q vssd1 vssd1 vccd1 vccd1 _4242_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_87_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7030_ _7030_/A _7030_/B vssd1 vssd1 vccd1 vccd1 _7031_/A sky130_fd_sc_hd__and2_1
XFILLER_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4173_ _4417_/A vssd1 vssd1 vccd1 vccd1 _4173_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6814_ _6814_/A vssd1 vssd1 vccd1 vccd1 _6814_/X sky130_fd_sc_hd__buf_1
XFILLER_23_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7794_ _7821_/CLK _7794_/D vssd1 vssd1 vccd1 vccd1 _7794_/Q sky130_fd_sc_hd__dfxtp_1
X_3957_ _3957_/A vssd1 vssd1 vccd1 vccd1 _7650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6676_ _6676_/A vssd1 vssd1 vccd1 vccd1 _6702_/C sky130_fd_sc_hd__clkbuf_2
X_3888_ _7527_/Q _4111_/A _4394_/B vssd1 vssd1 vccd1 vccd1 _4955_/B sky130_fd_sc_hd__or3b_1
X_5627_ _6396_/B _5627_/B vssd1 vssd1 vccd1 vccd1 _5627_/X sky130_fd_sc_hd__or2_1
XFILLER_117_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5558_ _7180_/Q _7361_/Q _7717_/Q _7257_/Q _5520_/X _5521_/X vssd1 vssd1 vccd1 vccd1
+ _5558_/X sky130_fd_sc_hd__mux4_1
X_5825__284 _5825__284/A vssd1 vssd1 vccd1 vccd1 _7301_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4509_ _7439_/Q _4221_/X _4515_/S vssd1 vssd1 vccd1 vccd1 _4510_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7228_ _7331_/CLK _7228_/D vssd1 vssd1 vccd1 vccd1 _7228_/Q sky130_fd_sc_hd__dfxtp_1
X_5489_ _4291_/A _5483_/X _5485_/X _5488_/X _5421_/Y vssd1 vssd1 vccd1 vccd1 _5489_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7159_ _7684_/CLK _7159_/D vssd1 vssd1 vccd1 vccd1 _7159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5379__207 _5381__209/A vssd1 vssd1 vccd1 vccd1 _7179_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5832__288 _5833__289/A vssd1 vssd1 vccd1 vccd1 _7305_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3107_ clkbuf_0__3107_/X vssd1 vssd1 vccd1 vccd1 _6353__434/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7224_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_111_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4860_ _4860_/A vssd1 vssd1 vccd1 vccd1 _7255_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3811_ _4901_/D _4919_/A vssd1 vssd1 vccd1 vccd1 _3841_/S sky130_fd_sc_hd__or2_4
XFILLER_119_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3311_ clkbuf_0__3311_/X vssd1 vssd1 vccd1 vccd1 _6828__26/A sky130_fd_sc_hd__clkbuf_4
X_4791_ _4713_/X _7282_/Q _4795_/S vssd1 vssd1 vccd1 vccd1 _4792_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3742_ _3742_/A vssd1 vssd1 vccd1 vccd1 _7737_/D sky130_fd_sc_hd__clkbuf_1
X_3673_ _7762_/Q _3672_/X _3676_/S vssd1 vssd1 vccd1 vccd1 _3674_/A sky130_fd_sc_hd__mux2_1
X_6392_ _6392_/A vssd1 vssd1 vccd1 vccd1 _6392_/X sky130_fd_sc_hd__buf_1
X_5412_ _5520_/A vssd1 vssd1 vccd1 vccd1 _5427_/A sky130_fd_sc_hd__clkbuf_4
Xoutput102 _5124_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[18] sky130_fd_sc_hd__buf_2
Xoutput113 _5088_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[2] sky130_fd_sc_hd__buf_2
Xoutput124 _5039_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[11] sky130_fd_sc_hd__buf_2
XFILLER_114_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5343_ _5343_/A _5343_/B vssd1 vssd1 vccd1 vccd1 _7158_/D sky130_fd_sc_hd__nor2_1
XFILLER_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput146 _5082_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[31] sky130_fd_sc_hd__buf_2
Xoutput135 _5061_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[21] sky130_fd_sc_hd__buf_2
Xoutput157 _5009_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[3] sky130_fd_sc_hd__buf_2
XFILLER_99_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput168 _5195_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[16] sky130_fd_sc_hd__buf_2
XFILLER_114_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5274_ _5274_/A vssd1 vssd1 vccd1 vccd1 _5274_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3141_ _6514_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3141_/X sky130_fd_sc_hd__clkbuf_16
Xoutput179 _5225_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[26] sky130_fd_sc_hd__buf_2
XFILLER_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4225_ _7544_/Q _4224_/X _4231_/S vssd1 vssd1 vccd1 vccd1 _4226_/A sky130_fd_sc_hd__mux2_1
X_7013_ _6902_/S _6324_/A _7013_/S vssd1 vssd1 vccd1 vccd1 _7014_/B sky130_fd_sc_hd__mux2_1
XFILLER_101_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4156_ _4155_/X _7569_/Q _4165_/S vssd1 vssd1 vccd1 vccd1 _4157_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4087_ _4087_/A vssd1 vssd1 vccd1 vccd1 _7596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7846_ _7855_/CLK _7846_/D vssd1 vssd1 vccd1 vccd1 _7846_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_24_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4989_ _7348_/Q _7347_/Q _7346_/Q _7345_/Q vssd1 vssd1 vccd1 vccd1 _5138_/C sky130_fd_sc_hd__and4bb_2
X_7777_ _7777_/CLK _7777_/D vssd1 vssd1 vccd1 vccd1 _7777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6659_ _6583_/B _6677_/A _6656_/X _6658_/X vssd1 vssd1 vccd1 vccd1 _6659_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_109_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5385__211 _5385__211/A vssd1 vssd1 vccd1 vccd1 _7183_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput26 caravel_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 _5232_/B sky130_fd_sc_hd__clkbuf_1
Xinput15 caravel_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 _5209_/B sky130_fd_sc_hd__clkbuf_1
Xinput37 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__buf_4
XFILLER_116_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6536__98 _6537__99/A vssd1 vssd1 vccd1 vccd1 _7643_/CLK sky130_fd_sc_hd__inv_2
Xinput48 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _5094_/A sky130_fd_sc_hd__buf_6
Xinput59 wbs_data_i[14] vssd1 vssd1 vccd1 vccd1 _5044_/A sky130_fd_sc_hd__buf_6
XFILLER_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6785__166 _6787__168/A vssd1 vssd1 vccd1 vccd1 _7733_/CLK sky130_fd_sc_hd__inv_2
X_6854__47 _6855__48/A vssd1 vssd1 vccd1 vccd1 _7789_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6132__346 _6133__347/A vssd1 vssd1 vccd1 vccd1 _7395_/CLK sky130_fd_sc_hd__inv_2
X_6171__373 _6172__374/A vssd1 vssd1 vccd1 vccd1 _7425_/CLK sky130_fd_sc_hd__inv_2
X_4010_ _4131_/D _4072_/B vssd1 vssd1 vccd1 vccd1 _4026_/S sky130_fd_sc_hd__or2_2
XFILLER_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5774__242 _5775__243/A vssd1 vssd1 vccd1 vccd1 _7259_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5961_ _7408_/Q _7349_/Q _7416_/Q _7397_/Q _4446_/A _5954_/X vssd1 vssd1 vccd1 vccd1
+ _5961_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6440__501 _6442__503/A vssd1 vssd1 vccd1 vccd1 _7566_/CLK sky130_fd_sc_hd__inv_2
X_4912_ _4912_/A vssd1 vssd1 vccd1 vccd1 _7232_/D sky130_fd_sc_hd__clkbuf_1
X_7700_ _7700_/CLK _7700_/D vssd1 vssd1 vccd1 vccd1 _7700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5892_ _5892_/A _5892_/B vssd1 vssd1 vccd1 vccd1 _5908_/S sky130_fd_sc_hd__and2_2
X_7631_ _7631_/CLK _7631_/D vssd1 vssd1 vccd1 vccd1 _7631_/Q sky130_fd_sc_hd__dfxtp_1
X_4843_ _4823_/X _7262_/Q _4845_/S vssd1 vssd1 vccd1 vccd1 _4844_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7562_ _7562_/CLK _7562_/D vssd1 vssd1 vccd1 vccd1 _7562_/Q sky130_fd_sc_hd__dfxtp_1
X_4774_ _4774_/A vssd1 vssd1 vccd1 vccd1 _7290_/D sky130_fd_sc_hd__clkbuf_1
X_7493_ _7493_/CLK _7493_/D vssd1 vssd1 vccd1 vccd1 _7493_/Q sky130_fd_sc_hd__dfxtp_1
X_6397__466 _6400__469/A vssd1 vssd1 vccd1 vccd1 _7531_/CLK sky130_fd_sc_hd__inv_2
X_3725_ _4614_/D _3928_/B vssd1 vssd1 vccd1 vccd1 _3741_/S sky130_fd_sc_hd__or2_2
X_6513_ _6770_/A vssd1 vssd1 vccd1 vccd1 _6513_/X sky130_fd_sc_hd__buf_1
XFILLER_9_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6444_ _6444_/A vssd1 vssd1 vccd1 vccd1 _6444_/X sky130_fd_sc_hd__buf_1
X_3656_ _3656_/A vssd1 vssd1 vccd1 vccd1 _7768_/D sky130_fd_sc_hd__clkbuf_1
X_3587_ _3587_/A vssd1 vssd1 vccd1 vccd1 _7092_/A sky130_fd_sc_hd__buf_6
X_5326_ _7092_/A _7152_/Q _5328_/S vssd1 vssd1 vccd1 vccd1 _5327_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3087_ clkbuf_0__3087_/X vssd1 vssd1 vccd1 vccd1 _6293__404/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3124_ _6432_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3124_/X sky130_fd_sc_hd__clkbuf_16
X_4208_ _4208_/A vssd1 vssd1 vccd1 vccd1 _7549_/D sky130_fd_sc_hd__clkbuf_1
X_5188_ _5236_/B vssd1 vssd1 vccd1 vccd1 _5198_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4139_ _4057_/X _7575_/Q _4141_/S vssd1 vssd1 vccd1 vccd1 _4140_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7829_ _7829_/CLK _7829_/D vssd1 vssd1 vccd1 vccd1 _7829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3510_ _7208_/Q _7209_/Q _7210_/Q _7211_/Q vssd1 vssd1 vccd1 vccd1 _5435_/B sky130_fd_sc_hd__or4_1
X_6509__76 _6510__77/A vssd1 vssd1 vccd1 vccd1 _7621_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4490_ _4490_/A vssd1 vssd1 vccd1 vccd1 _7448_/D sky130_fd_sc_hd__clkbuf_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5122_/A vssd1 vssd1 vccd1 vccd1 _5120_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6827__25 _6828__26/A vssd1 vssd1 vccd1 vccd1 _7767_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6091_ _7578_/Q _7388_/Q _7736_/Q _7634_/Q _6002_/X _4450_/A vssd1 vssd1 vccd1 vccd1
+ _6091_/X sky130_fd_sc_hd__mux4_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5042_/A _5044_/B vssd1 vssd1 vccd1 vccd1 _5043_/A sky130_fd_sc_hd__or2_1
XFILLER_85_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6993_ _6993_/A _6993_/B _6993_/C _6993_/D vssd1 vssd1 vccd1 vccd1 _6994_/B sky130_fd_sc_hd__and4_1
XFILLER_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5944_ _7459_/Q vssd1 vssd1 vccd1 vccd1 _6095_/A sky130_fd_sc_hd__clkinv_2
XFILLER_18_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5875_ _5890_/S vssd1 vssd1 vccd1 vccd1 _5884_/S sky130_fd_sc_hd__clkbuf_2
X_6405__473 _6406__474/A vssd1 vssd1 vccd1 vccd1 _7538_/CLK sky130_fd_sc_hd__inv_2
X_7614_ _7614_/CLK _7614_/D vssd1 vssd1 vccd1 vccd1 _7614_/Q sky130_fd_sc_hd__dfxtp_1
X_4826_ _7468_/Q vssd1 vssd1 vccd1 vccd1 _4826_/X sky130_fd_sc_hd__buf_2
X_7545_ _7545_/CLK _7545_/D vssd1 vssd1 vccd1 vccd1 _7545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4757_ _4716_/X _7297_/Q _4759_/S vssd1 vssd1 vccd1 vccd1 _4758_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3708_ _3708_/A vssd1 vssd1 vccd1 vccd1 _7750_/D sky130_fd_sc_hd__clkbuf_1
X_7476_ _7477_/CLK _7476_/D vssd1 vssd1 vccd1 vccd1 _7476_/Q sky130_fd_sc_hd__dfxtp_1
X_4688_ _4703_/S vssd1 vssd1 vccd1 vccd1 _4697_/S sky130_fd_sc_hd__buf_2
X_3639_ _3562_/X _7773_/Q _3641_/S vssd1 vssd1 vccd1 vccd1 _3640_/A sky130_fd_sc_hd__mux2_1
X_6178__379 _6178__379/A vssd1 vssd1 vccd1 vccd1 _7431_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3139_ clkbuf_0__3139_/X vssd1 vssd1 vccd1 vccd1 _6510__77/A sky130_fd_sc_hd__clkbuf_4
X_5309_ _5303_/X _7342_/Q _5307_/X _5308_/X _7142_/Q vssd1 vssd1 vccd1 vccd1 _7142_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_103_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6729__123 _6730__124/A vssd1 vssd1 vccd1 vccd1 _7689_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6447__507 _6448__508/A vssd1 vssd1 vccd1 vccd1 _7572_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3107_ _6348_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3107_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7679_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_17_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3990_ _3990_/A vssd1 vssd1 vccd1 vccd1 _7635_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5660_ _5660_/A vssd1 vssd1 vccd1 vccd1 _7197_/D sky130_fd_sc_hd__clkbuf_1
X_4611_ _4611_/A vssd1 vssd1 vccd1 vccd1 _7390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5591_ _7694_/Q _7283_/Q _7166_/Q _7275_/Q _5467_/X _5413_/X vssd1 vssd1 vccd1 vccd1
+ _5591_/X sky130_fd_sc_hd__mux4_1
X_7330_ _7372_/CLK _7330_/D vssd1 vssd1 vccd1 vccd1 _7330_/Q sky130_fd_sc_hd__dfxtp_1
X_4542_ _4632_/A _4668_/B vssd1 vssd1 vccd1 vccd1 _4558_/S sky130_fd_sc_hd__nand2_2
XFILLER_116_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6290__401 _6292__403/A vssd1 vssd1 vccd1 vccd1 _7454_/CLK sky130_fd_sc_hd__inv_2
X_4473_ _4399_/X _7455_/Q _4479_/S vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__mux2_1
X_7261_ _7261_/CLK _7261_/D vssd1 vssd1 vccd1 vccd1 _7261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6212_ _6930_/A _6233_/D _6933_/A vssd1 vssd1 vccd1 vccd1 _6884_/B sky130_fd_sc_hd__a21o_1
X_7192_ _7226_/CLK _7192_/D vssd1 vssd1 vccd1 vccd1 _7192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6074_ _7727_/Q _7711_/Q _7430_/Q _7492_/Q _5935_/X _5937_/X vssd1 vssd1 vccd1 vccd1
+ _6074_/X sky130_fd_sc_hd__mux4_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _7026_/A _5033_/B vssd1 vssd1 vccd1 vccd1 _5026_/A sky130_fd_sc_hd__or2_1
XINSDIODE2_39 _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_17 _5214_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_28 _5085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3140_ clkbuf_0__3140_/X vssd1 vssd1 vccd1 vccd1 _6520_/A sky130_fd_sc_hd__clkbuf_4
X_6976_ _6975_/Y _6916_/A _6983_/A _6974_/B vssd1 vssd1 vccd1 vccd1 _6976_/X sky130_fd_sc_hd__a211o_1
XFILLER_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5858_ _5031_/A _7325_/Q _5866_/S vssd1 vssd1 vccd1 vccd1 _5859_/A sky130_fd_sc_hd__mux2_1
X_4809_ _4808_/X _7275_/Q _4818_/S vssd1 vssd1 vccd1 vccd1 _4810_/A sky130_fd_sc_hd__mux2_1
X_5789_ _5789_/A vssd1 vssd1 vccd1 vccd1 _5789_/X sky130_fd_sc_hd__buf_1
XFILLER_107_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7528_ _7528_/CLK _7528_/D vssd1 vssd1 vccd1 vccd1 _7528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7459_ _7459_/CLK _7459_/D vssd1 vssd1 vccd1 vccd1 _7459_/Q sky130_fd_sc_hd__dfxtp_1
X_6453__511 _6455__513/A vssd1 vssd1 vccd1 vccd1 _7576_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6742__131 _6743__132/A vssd1 vssd1 vccd1 vccd1 _7698_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2990_ clkbuf_0__2990_/X vssd1 vssd1 vccd1 vccd1 _6152__358/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5712_ _7217_/Q _7332_/Q _5714_/S vssd1 vssd1 vccd1 vccd1 _5713_/A sky130_fd_sc_hd__mux2_1
X_3973_ _4243_/B _3973_/B vssd1 vssd1 vccd1 vccd1 _3989_/S sky130_fd_sc_hd__nor2_4
X_6692_ _6656_/X _6658_/X _6602_/A vssd1 vssd1 vccd1 vccd1 _6692_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5643_ _7845_/Q vssd1 vssd1 vccd1 vccd1 _6249_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_117_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5574_ _7181_/Q _7362_/Q _7718_/Q _7258_/Q _5481_/X _5506_/X vssd1 vssd1 vccd1 vccd1
+ _5574_/X sky130_fd_sc_hd__mux4_1
X_4525_ _4242_/X _7431_/Q _4533_/S vssd1 vssd1 vccd1 vccd1 _4526_/A sky130_fd_sc_hd__mux2_1
X_7313_ _7313_/CLK _7313_/D vssd1 vssd1 vccd1 vccd1 _7313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4456_ _4452_/A _4459_/A _4455_/Y vssd1 vssd1 vccd1 vccd1 _7460_/D sky130_fd_sc_hd__o21a_1
X_7244_ _7244_/CLK _7244_/D vssd1 vssd1 vccd1 vccd1 _7244_/Q sky130_fd_sc_hd__dfxtp_1
X_4387_ _7488_/Q _3944_/A _4391_/S vssd1 vssd1 vccd1 vccd1 _4388_/A sky130_fd_sc_hd__mux2_1
X_7175_ _7175_/CLK _7175_/D vssd1 vssd1 vccd1 vccd1 _7175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _7758_/Q _7750_/Q _7742_/Q _7656_/Q _4465_/A _5954_/X vssd1 vssd1 vccd1 vccd1
+ _6057_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5008_ _5892_/A _5087_/B vssd1 vssd1 vccd1 vccd1 _5009_/A sky130_fd_sc_hd__and2_1
XFILLER_85_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3123_ clkbuf_0__3123_/X vssd1 vssd1 vccd1 vccd1 _6431__494/A sky130_fd_sc_hd__clkbuf_4
X_6959_ _6957_/Y _6958_/X _6954_/X vssd1 vssd1 vccd1 vccd1 _7806_/D sky130_fd_sc_hd__a21oi_1
XFILLER_41_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6297__407 _6298__408/A vssd1 vssd1 vccd1 vccd1 _7460_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6377__453 _6378__454/A vssd1 vssd1 vccd1 vccd1 _7516_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6488__59 _6488__59/A vssd1 vssd1 vccd1 vccd1 _7604_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2769_ clkbuf_0__2769_/X vssd1 vssd1 vccd1 vccd1 _5792__257/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5290_ _5287_/X hold3/X _5283_/X _5284_/X _7131_/Q vssd1 vssd1 vccd1 vccd1 _7131_/D
+ sky130_fd_sc_hd__o32a_1
X_4310_ _6396_/A _4310_/B vssd1 vssd1 vccd1 vccd1 _4310_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6749__137 _6749__137/A vssd1 vssd1 vccd1 vccd1 _7704_/CLK sky130_fd_sc_hd__inv_2
X_4241_ _4241_/A vssd1 vssd1 vccd1 vccd1 _7539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5738__213 _5739__214/A vssd1 vssd1 vccd1 vccd1 _7230_/CLK sky130_fd_sc_hd__inv_2
X_4172_ _4172_/A vssd1 vssd1 vccd1 vccd1 _7564_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7793_ _7799_/CLK _7793_/D vssd1 vssd1 vccd1 vccd1 _7793_/Q sky130_fd_sc_hd__dfxtp_1
X_3956_ _3926_/X _7650_/Q _3964_/S vssd1 vssd1 vccd1 vccd1 _3957_/A sky130_fd_sc_hd__mux2_1
X_7860__234 vssd1 vssd1 vccd1 vccd1 partID[6] _7860__234/LO sky130_fd_sc_hd__conb_1
XFILLER_51_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6675_ _6640_/C _6661_/X _6595_/B vssd1 vssd1 vccd1 vccd1 _6675_/X sky130_fd_sc_hd__a21bo_1
XFILLER_50_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3887_ _3907_/B vssd1 vssd1 vccd1 vccd1 _4394_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5626_ _5434_/A _5616_/X _5625_/Y _5492_/A vssd1 vssd1 vccd1 vccd1 _5627_/B sky130_fd_sc_hd__a211oi_1
XFILLER_117_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5557_ _7583_/Q _7567_/Q _7551_/Q _7543_/Q _5520_/X _5521_/X vssd1 vssd1 vccd1 vccd1
+ _5557_/X sky130_fd_sc_hd__mux4_1
X_4508_ _4508_/A vssd1 vssd1 vccd1 vccd1 _7440_/D sky130_fd_sc_hd__clkbuf_1
X_5488_ _5572_/S _5487_/X _5404_/A vssd1 vssd1 vccd1 vccd1 _5488_/X sky130_fd_sc_hd__a21o_1
XFILLER_105_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4439_ _6051_/A vssd1 vssd1 vccd1 vccd1 _4451_/A sky130_fd_sc_hd__buf_2
XFILLER_78_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7227_ _7854_/CLK _7227_/D vssd1 vssd1 vccd1 vccd1 _7227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7158_ _7685_/CLK _7158_/D vssd1 vssd1 vccd1 vccd1 _7158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7089_ _7070_/X _7089_/B vssd1 vssd1 vccd1 vccd1 _7090_/A sky130_fd_sc_hd__and2b_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3106_ clkbuf_0__3106_/X vssd1 vssd1 vccd1 vccd1 _6347__429/A sky130_fd_sc_hd__clkbuf_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4790_ _4790_/A vssd1 vssd1 vccd1 vccd1 _7283_/D sky130_fd_sc_hd__clkbuf_1
X_3810_ _3907_/B _4111_/A _4394_/A vssd1 vssd1 vccd1 vccd1 _4919_/A sky130_fd_sc_hd__or3b_1
Xclkbuf_1_1_0__3310_ clkbuf_0__3310_/X vssd1 vssd1 vccd1 vccd1 _6825__24/A sky130_fd_sc_hd__clkbuf_4
X_3741_ _3721_/X _7737_/Q _3741_/S vssd1 vssd1 vccd1 vccd1 _3742_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3672_ _7823_/Q vssd1 vssd1 vccd1 vccd1 _3672_/X sky130_fd_sc_hd__buf_4
X_5411_ _7518_/Q vssd1 vssd1 vccd1 vccd1 _5520_/A sky130_fd_sc_hd__buf_2
Xoutput103 _5126_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[19] sky130_fd_sc_hd__buf_2
Xoutput114 _5091_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[3] sky130_fd_sc_hd__buf_2
Xoutput125 _5041_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[12] sky130_fd_sc_hd__buf_2
X_5342_ _7158_/Q _4998_/A _5274_/A _5317_/B vssd1 vssd1 vccd1 vccd1 _5343_/B sky130_fd_sc_hd__o211a_1
Xoutput136 _5063_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[22] sky130_fd_sc_hd__buf_2
Xoutput147 _5021_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[3] sky130_fd_sc_hd__buf_2
Xoutput158 _4997_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_stb_o sky130_fd_sc_hd__buf_2
Xclkbuf_0__3140_ _6513_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3140_/X sky130_fd_sc_hd__clkbuf_16
X_5273_ _5270_/X _7153_/Q _5262_/X _5266_/X _7121_/Q vssd1 vssd1 vccd1 vccd1 _7121_/D
+ sky130_fd_sc_hd__o32a_1
Xoutput169 _5197_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[17] sky130_fd_sc_hd__buf_2
X_7012_ _7821_/Q _7013_/S _7011_/X _7003_/X vssd1 vssd1 vccd1 vccd1 _7820_/D sky130_fd_sc_hd__o211a_1
XFILLER_114_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4224_ _7473_/Q vssd1 vssd1 vccd1 vccd1 _4224_/X sky130_fd_sc_hd__buf_4
X_4155_ _4399_/A vssd1 vssd1 vccd1 vccd1 _4155_/X sky130_fd_sc_hd__buf_2
XFILLER_110_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4086_ _4066_/X _7596_/Q _4088_/S vssd1 vssd1 vccd1 vccd1 _4087_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7845_ _7845_/CLK _7845_/D vssd1 vssd1 vccd1 vccd1 _7845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7776_ _7776_/CLK _7776_/D vssd1 vssd1 vccd1 vccd1 _7776_/Q sky130_fd_sc_hd__dfxtp_1
X_4988_ _4988_/A vssd1 vssd1 vccd1 vccd1 _7109_/D sky130_fd_sc_hd__clkbuf_1
X_3939_ _3938_/X _7655_/Q _3942_/S vssd1 vssd1 vccd1 vccd1 _3940_/A sky130_fd_sc_hd__mux2_1
X_6727_ _7687_/Q _5996_/A _6723_/C _6726_/X vssd1 vssd1 vccd1 vccd1 _7687_/D sky130_fd_sc_hd__a31o_1
X_6658_ _6684_/A vssd1 vssd1 vccd1 vccd1 _6658_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5609_ _7183_/Q _7364_/Q _7720_/Q _7260_/Q _5486_/X _5426_/X vssd1 vssd1 vccd1 vccd1
+ _5609_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6589_ _7674_/Q vssd1 vssd1 vccd1 vccd1 _6595_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput27 caravel_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 _5234_/B sky130_fd_sc_hd__clkbuf_1
Xinput16 caravel_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 _5211_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_52_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput38 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 _5105_/A sky130_fd_sc_hd__buf_4
Xinput49 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 _5096_/A sky130_fd_sc_hd__buf_6
XFILLER_6_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5960_ _5953_/X _5955_/X _5958_/X _5959_/X vssd1 vssd1 vccd1 vccd1 _5960_/X sky130_fd_sc_hd__o211a_1
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5891_ _5891_/A vssd1 vssd1 vccd1 vccd1 _7340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4911_ _4817_/X _7232_/Q _4911_/S vssd1 vssd1 vccd1 vccd1 _4912_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7630_ _7630_/CLK _7630_/D vssd1 vssd1 vccd1 vccd1 _7630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4842_ _4842_/A vssd1 vssd1 vccd1 vccd1 _7263_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7561_ _7561_/CLK _7561_/D vssd1 vssd1 vccd1 vccd1 _7561_/Q sky130_fd_sc_hd__dfxtp_1
X_4773_ _4713_/X _7290_/Q _4777_/S vssd1 vssd1 vccd1 vccd1 _4774_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7492_ _7492_/CLK _7492_/D vssd1 vssd1 vccd1 vccd1 _7492_/Q sky130_fd_sc_hd__dfxtp_1
X_3724_ _3724_/A _3927_/B _3927_/C _3678_/A vssd1 vssd1 vccd1 vccd1 _4614_/D sky130_fd_sc_hd__or4b_4
X_3655_ _7768_/Q _3649_/X _3667_/S vssd1 vssd1 vccd1 vccd1 _3656_/A sky130_fd_sc_hd__mux2_1
X_3586_ _3650_/A vssd1 vssd1 vccd1 vccd1 _4424_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5325_ _5325_/A vssd1 vssd1 vccd1 vccd1 _7151_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3086_ clkbuf_0__3086_/X vssd1 vssd1 vccd1 vccd1 _6287__399/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3123_ _6426_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3123_/X sky130_fd_sc_hd__clkbuf_16
X_5256_ _5358_/A vssd1 vssd1 vccd1 vccd1 _5256_/X sky130_fd_sc_hd__buf_1
XFILLER_102_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4207_ _4167_/X _7549_/Q _4211_/S vssd1 vssd1 vccd1 vccd1 _4208_/A sky130_fd_sc_hd__mux2_1
X_5187_ _5187_/A vssd1 vssd1 vccd1 vccd1 _5187_/X sky130_fd_sc_hd__buf_2
XFILLER_83_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4138_ _4138_/A vssd1 vssd1 vccd1 vccd1 _7576_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4069_ _7822_/Q vssd1 vssd1 vccd1 vccd1 _4069_/X sky130_fd_sc_hd__buf_2
XFILLER_44_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7828_ _7829_/CLK _7828_/D vssd1 vssd1 vccd1 vccd1 _7828_/Q sky130_fd_sc_hd__dfxtp_1
X_7759_ _7759_/CLK _7759_/D vssd1 vssd1 vccd1 vccd1 _7759_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2769_ _5789_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2769_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7873__200 vssd1 vssd1 vccd1 vccd1 _7873__200/HI core0Index[7] sky130_fd_sc_hd__conb_1
XFILLER_79_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6791__171 _6792__172/A vssd1 vssd1 vccd1 vccd1 _7738_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5845__299 _5845__299/A vssd1 vssd1 vccd1 vccd1 _7316_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5110_ _5110_/A vssd1 vssd1 vccd1 vccd1 _5110_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _7626_/Q _7618_/Q _7610_/Q _7602_/Q _5935_/X _5937_/X vssd1 vssd1 vccd1 vccd1
+ _6090_/X sky130_fd_sc_hd__mux4_2
X_5041_ _5041_/A vssd1 vssd1 vccd1 vccd1 _5041_/X sky130_fd_sc_hd__clkbuf_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_26_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6992_ _6860_/Y _6861_/X _6991_/X _6250_/C _6250_/B vssd1 vssd1 vccd1 vccd1 _6993_/D
+ sky130_fd_sc_hd__o2111a_1
X_5943_ _7571_/Q _7381_/Q _7729_/Q _7627_/Q _5942_/X _4465_/X vssd1 vssd1 vccd1 vccd1
+ _5943_/X sky130_fd_sc_hd__mux4_1
X_5874_ _5874_/A _5892_/B vssd1 vssd1 vccd1 vccd1 _5890_/S sky130_fd_sc_hd__nand2_2
X_7613_ _7613_/CLK _7613_/D vssd1 vssd1 vccd1 vccd1 _7613_/Q sky130_fd_sc_hd__dfxtp_1
X_4825_ _4825_/A vssd1 vssd1 vccd1 vccd1 _7270_/D sky130_fd_sc_hd__clkbuf_1
X_7544_ _7544_/CLK _7544_/D vssd1 vssd1 vccd1 vccd1 _7544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4756_ _4756_/A vssd1 vssd1 vccd1 vccd1 _7298_/D sky130_fd_sc_hd__clkbuf_1
X_3707_ _3706_/X _7750_/Q _3713_/S vssd1 vssd1 vccd1 vccd1 _3708_/A sky130_fd_sc_hd__mux2_1
X_7475_ _7821_/CLK _7475_/D vssd1 vssd1 vccd1 vccd1 _7475_/Q sky130_fd_sc_hd__dfxtp_1
X_4687_ _4901_/A _4901_/B _4731_/C _4847_/B vssd1 vssd1 vccd1 vccd1 _4703_/S sky130_fd_sc_hd__or4_4
X_3638_ _3638_/A vssd1 vssd1 vccd1 vccd1 _7774_/D sky130_fd_sc_hd__clkbuf_1
X_6426_ _6432_/A vssd1 vssd1 vccd1 vccd1 _6426_/X sky130_fd_sc_hd__buf_1
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3569_ _7824_/Q vssd1 vssd1 vccd1 vccd1 _3944_/A sky130_fd_sc_hd__clkbuf_4
X_6371__448 _6371__448/A vssd1 vssd1 vccd1 vccd1 _7511_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3138_ clkbuf_0__3138_/X vssd1 vssd1 vccd1 vccd1 _6506__74/A sky130_fd_sc_hd__clkbuf_4
X_5308_ _5308_/A vssd1 vssd1 vccd1 vccd1 _5308_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3106_ _6342_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3106_/X sky130_fd_sc_hd__clkbuf_16
X_6288_ _6294_/A vssd1 vssd1 vccd1 vccd1 _6288_/X sky130_fd_sc_hd__buf_1
XFILLER_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5239_ _5239_/A vssd1 vssd1 vccd1 vccd1 _5338_/A sky130_fd_sc_hd__buf_2
XFILLER_102_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4610_ _4262_/X _7390_/Q _4612_/S vssd1 vssd1 vccd1 vccd1 _4611_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5590_ _5590_/A _5590_/B vssd1 vssd1 vccd1 vccd1 _5590_/X sky130_fd_sc_hd__and2_1
XFILLER_116_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4541_ _3745_/A _4614_/B _4614_/A vssd1 vssd1 vccd1 vccd1 _4668_/B sky130_fd_sc_hd__and3b_2
X_7260_ _7260_/CLK _7260_/D vssd1 vssd1 vccd1 vccd1 _7260_/Q sky130_fd_sc_hd__dfxtp_1
X_4472_ _4472_/A vssd1 vssd1 vccd1 vccd1 _7456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7191_ _7839_/CLK _7191_/D vssd1 vssd1 vccd1 vccd1 _7191_/Q sky130_fd_sc_hd__dfxtp_1
X_6211_ _6933_/A _6930_/A _6233_/D vssd1 vssd1 vccd1 vccd1 _6884_/A sky130_fd_sc_hd__nand3_1
XFILLER_112_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6142_ _6142_/A vssd1 vssd1 vccd1 vccd1 _6142_/X sky130_fd_sc_hd__buf_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6073_ _7577_/Q _7387_/Q _7735_/Q _7633_/Q _5998_/A _4450_/A vssd1 vssd1 vccd1 vccd1
+ _6073_/X sky130_fd_sc_hd__mux4_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5081_/B vssd1 vssd1 vccd1 vccd1 _5033_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_29 _5085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_18 _5214_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6798__177 _6798__177/A vssd1 vssd1 vccd1 vccd1 _7744_/CLK sky130_fd_sc_hd__inv_2
X_6975_ _7811_/Q vssd1 vssd1 vccd1 vccd1 _6975_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5787__253 _5788__254/A vssd1 vssd1 vccd1 vccd1 _7270_/CLK sky130_fd_sc_hd__inv_2
X_5857_ _5872_/S vssd1 vssd1 vccd1 vccd1 _5866_/S sky130_fd_sc_hd__buf_2
XFILLER_70_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4808_ _7474_/Q vssd1 vssd1 vccd1 vccd1 _4808_/X sky130_fd_sc_hd__buf_2
XFILLER_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4739_ _4716_/X _7305_/Q _4741_/S vssd1 vssd1 vccd1 vccd1 _4740_/A sky130_fd_sc_hd__mux2_1
X_7527_ _7527_/CLK _7527_/D vssd1 vssd1 vccd1 vccd1 _7527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7458_ _7458_/CLK _7458_/D vssd1 vssd1 vccd1 vccd1 _7458_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7389_ _7389_/CLK _7389_/D vssd1 vssd1 vccd1 vccd1 _7389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5711_ _5711_/A vssd1 vssd1 vccd1 vccd1 _7216_/D sky130_fd_sc_hd__clkbuf_1
X_3972_ _4131_/A _4424_/A _3991_/C vssd1 vssd1 vccd1 vccd1 _3973_/B sky130_fd_sc_hd__nand3_2
X_6691_ _6688_/X _6689_/X _6690_/X vssd1 vssd1 vccd1 vccd1 _7676_/D sky130_fd_sc_hd__a21oi_1
X_5642_ _5642_/A vssd1 vssd1 vccd1 vccd1 _7193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5573_ _7584_/Q _7568_/Q _7552_/Q _7544_/Q _5512_/X _5513_/X vssd1 vssd1 vccd1 vccd1
+ _5573_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4524_ _4539_/S vssd1 vssd1 vccd1 vccd1 _4533_/S sky130_fd_sc_hd__buf_2
X_7312_ _7312_/CLK _7312_/D vssd1 vssd1 vccd1 vccd1 _7312_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_116_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4455_ _6325_/A _4455_/B vssd1 vssd1 vccd1 vccd1 _4455_/Y sky130_fd_sc_hd__nor2_1
X_7243_ _7243_/CLK _7243_/D vssd1 vssd1 vccd1 vccd1 _7243_/Q sky130_fd_sc_hd__dfxtp_1
X_4386_ _4386_/A vssd1 vssd1 vccd1 vccd1 _7489_/D sky130_fd_sc_hd__clkbuf_1
X_7174_ _7174_/CLK _7174_/D vssd1 vssd1 vccd1 vccd1 _7174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6056_ _7726_/Q _7710_/Q _7429_/Q _7491_/Q _6024_/X _5998_/X vssd1 vssd1 vccd1 vccd1
+ _6056_/X sky130_fd_sc_hd__mux4_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _5007_/A vssd1 vssd1 vccd1 vccd1 _5007_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3122_ clkbuf_0__3122_/X vssd1 vssd1 vccd1 vccd1 _6422__486/A sky130_fd_sc_hd__clkbuf_4
X_6958_ _6943_/X _6919_/X _6889_/B vssd1 vssd1 vccd1 vccd1 _6958_/X sky130_fd_sc_hd__a21o_1
X_5909_ _5909_/A vssd1 vssd1 vccd1 vccd1 _7348_/D sky130_fd_sc_hd__clkbuf_1
X_6889_ _7843_/Q _6889_/B vssd1 vssd1 vccd1 vccd1 _6892_/C sky130_fd_sc_hd__xor2_1
XFILLER_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6418__484 _6418__484/A vssd1 vssd1 vccd1 vccd1 _7549_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__2768_ clkbuf_0__2768_/X vssd1 vssd1 vccd1 vccd1 _5785__251/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4240_ _7539_/Q _4239_/X _4240_/S vssd1 vssd1 vccd1 vccd1 _4241_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4171_ _4170_/X _7564_/Q _4174_/S vssd1 vssd1 vccd1 vccd1 _4172_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7792_ _7792_/CLK _7792_/D vssd1 vssd1 vccd1 vccd1 _7792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3955_ _3970_/S vssd1 vssd1 vccd1 vccd1 _3964_/S sky130_fd_sc_hd__buf_2
XFILLER_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6674_ _6672_/X _6673_/X _6665_/X vssd1 vssd1 vccd1 vccd1 _7672_/D sky130_fd_sc_hd__a21oi_1
X_3886_ _4280_/A _4194_/A _4194_/B vssd1 vssd1 vccd1 vccd1 _4919_/B sky130_fd_sc_hd__or3b_2
X_5625_ _5620_/X _5624_/X _5434_/A vssd1 vssd1 vccd1 vccd1 _5625_/Y sky130_fd_sc_hd__a21oi_1
X_5556_ _5554_/X _5555_/X _5575_/S vssd1 vssd1 vccd1 vccd1 _5556_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4507_ _7440_/Q _4213_/X _4515_/S vssd1 vssd1 vccd1 vccd1 _4508_/A sky130_fd_sc_hd__mux2_1
X_5487_ _7689_/Q _7278_/Q _7161_/Q _7270_/Q _5521_/A _5486_/X vssd1 vssd1 vccd1 vccd1
+ _5487_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4438_ _7459_/Q vssd1 vssd1 vccd1 vccd1 _6051_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7226_ _7226_/CLK _7226_/D vssd1 vssd1 vccd1 vccd1 _7226_/Q sky130_fd_sc_hd__dfxtp_1
X_7157_ _7687_/CLK _7157_/D vssd1 vssd1 vccd1 vccd1 _7157_/Q sky130_fd_sc_hd__dfxtp_1
X_4369_ _4167_/X _7496_/Q _4373_/S vssd1 vssd1 vccd1 vccd1 _4370_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7088_ _7851_/Q _7024_/A _7100_/C vssd1 vssd1 vccd1 vccd1 _7089_/B sky130_fd_sc_hd__mux2_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6493__63 _6494__64/A vssd1 vssd1 vccd1 vccd1 _7608_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6039_ _7368_/Q _5931_/X _6038_/X _5996_/X vssd1 vssd1 vccd1 vccd1 _7368_/D sky130_fd_sc_hd__o211a_1
XFILLER_27_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3105_ clkbuf_0__3105_/X vssd1 vssd1 vccd1 vccd1 _6339__422/A sky130_fd_sc_hd__clkbuf_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6466__522 _6468__524/A vssd1 vssd1 vccd1 vccd1 _7587_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2766_ clkbuf_0__2766_/X vssd1 vssd1 vccd1 vccd1 _5776__244/A sky130_fd_sc_hd__clkbuf_16
XFILLER_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3740_ _3740_/A vssd1 vssd1 vccd1 vccd1 _7738_/D sky130_fd_sc_hd__clkbuf_1
X_6755__142 _6757__144/A vssd1 vssd1 vccd1 vccd1 _7709_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3671_ _3671_/A vssd1 vssd1 vccd1 vccd1 _7763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5410_ _5405_/X _5406_/X _5432_/S vssd1 vssd1 vccd1 vccd1 _5410_/X sky130_fd_sc_hd__mux2_1
Xoutput115 _5093_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[4] sky130_fd_sc_hd__buf_2
Xoutput104 _5086_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[1] sky130_fd_sc_hd__buf_2
X_5341_ _5317_/B _5336_/Y _5343_/A vssd1 vssd1 vccd1 vccd1 _7157_/D sky130_fd_sc_hd__a21oi_1
X_7890__217 vssd1 vssd1 vccd1 vccd1 _7890__217/HI manufacturerID[9] sky130_fd_sc_hd__conb_1
Xoutput159 _4999_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_we_o sky130_fd_sc_hd__buf_2
Xoutput126 _5043_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[13] sky130_fd_sc_hd__buf_2
Xoutput148 _5023_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[4] sky130_fd_sc_hd__buf_2
Xoutput137 _5065_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[23] sky130_fd_sc_hd__buf_2
X_5272_ _5270_/X _7152_/Q _5262_/X _5266_/X _7120_/Q vssd1 vssd1 vccd1 vccd1 _7120_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_99_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7011_ _6996_/A _6997_/A _7820_/Q vssd1 vssd1 vccd1 vccd1 _7011_/X sky130_fd_sc_hd__a21o_1
XFILLER_101_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4223_ _4223_/A vssd1 vssd1 vccd1 vccd1 _7545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4154_ _4154_/A vssd1 vssd1 vccd1 vccd1 _7570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4085_ _4085_/A vssd1 vssd1 vccd1 vccd1 _7597_/D sky130_fd_sc_hd__clkbuf_1
X_7844_ _7845_/CLK _7844_/D vssd1 vssd1 vccd1 vccd1 _7844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7775_ _7775_/CLK _7775_/D vssd1 vssd1 vccd1 vccd1 _7775_/Q sky130_fd_sc_hd__dfxtp_1
X_6726_ _6737_/S _6726_/B _6726_/C vssd1 vssd1 vccd1 vccd1 _6726_/X sky130_fd_sc_hd__and3_1
X_4987_ _7109_/Q _4417_/A _4987_/S vssd1 vssd1 vccd1 vccd1 _4988_/A sky130_fd_sc_hd__mux2_1
X_3938_ _3938_/A vssd1 vssd1 vccd1 vccd1 _3938_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_109_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6657_ _6657_/A vssd1 vssd1 vccd1 vccd1 _6684_/A sky130_fd_sc_hd__clkbuf_2
X_3869_ _3884_/S vssd1 vssd1 vccd1 vccd1 _3878_/S sky130_fd_sc_hd__buf_2
X_6588_ _6588_/A _6588_/B _6588_/C _6588_/D vssd1 vssd1 vccd1 vccd1 _6588_/X sky130_fd_sc_hd__and4_1
X_5608_ _7848_/Q vssd1 vssd1 vccd1 vccd1 _6872_/A sky130_fd_sc_hd__buf_2
X_5539_ _7582_/Q _7566_/Q _7550_/Q _7542_/Q _5502_/X _5521_/X vssd1 vssd1 vccd1 vccd1
+ _5539_/X sky130_fd_sc_hd__mux4_1
X_6335__419 _6335__419/A vssd1 vssd1 vccd1 vccd1 _7482_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_15_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7154_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_6548__107 _6548__107/A vssd1 vssd1 vccd1 vccd1 _7652_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7209_ _5246_/A _7209_/D vssd1 vssd1 vccd1 vccd1 _7209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5914__310 _5916__312/A vssd1 vssd1 vccd1 vccd1 _7351_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6268__384 _6268__384/A vssd1 vssd1 vccd1 vccd1 _7437_/CLK sky130_fd_sc_hd__inv_2
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput28 caravel_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_2
Xinput17 caravel_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 _5213_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput39 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 _5107_/A sky130_fd_sc_hd__buf_4
XFILLER_2_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5890_ _5064_/A _7340_/Q _5890_/S vssd1 vssd1 vccd1 vccd1 _5891_/A sky130_fd_sc_hd__mux2_1
X_4910_ _4910_/A vssd1 vssd1 vccd1 vccd1 _7233_/D sky130_fd_sc_hd__clkbuf_1
X_4841_ _4820_/X _7263_/Q _4845_/S vssd1 vssd1 vccd1 vccd1 _4842_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7560_ _7560_/CLK _7560_/D vssd1 vssd1 vccd1 vccd1 _7560_/Q sky130_fd_sc_hd__dfxtp_1
X_4772_ _4772_/A vssd1 vssd1 vccd1 vccd1 _7291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7491_ _7491_/CLK _7491_/D vssd1 vssd1 vccd1 vccd1 _7491_/Q sky130_fd_sc_hd__dfxtp_1
X_3723_ _3723_/A vssd1 vssd1 vccd1 vccd1 _7745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3654_ _3676_/S vssd1 vssd1 vccd1 vccd1 _3667_/S sky130_fd_sc_hd__buf_2
X_5781__248 _5782__249/A vssd1 vssd1 vccd1 vccd1 _7265_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3585_ _3585_/A vssd1 vssd1 vccd1 vccd1 _3724_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6373_ _6373_/A vssd1 vssd1 vccd1 vccd1 _6373_/X sky130_fd_sc_hd__buf_1
X_5324_ _7096_/A _7151_/Q _5328_/S vssd1 vssd1 vccd1 vccd1 _5325_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3085_ clkbuf_0__3085_/X vssd1 vssd1 vccd1 vccd1 _6277__390/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3122_ _6420_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3122_/X sky130_fd_sc_hd__clkbuf_16
X_5255_ _5382_/A vssd1 vssd1 vccd1 vccd1 _5255_/X sky130_fd_sc_hd__buf_1
X_4206_ _4206_/A vssd1 vssd1 vccd1 vccd1 _7550_/D sky130_fd_sc_hd__clkbuf_1
X_5186_ _7130_/Q _5173_/X input7/X _5177_/X _5185_/X vssd1 vssd1 vccd1 vccd1 _5186_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_110_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4137_ _4054_/X _7576_/Q _4141_/S vssd1 vssd1 vccd1 vccd1 _4138_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4068_ _4068_/A vssd1 vssd1 vccd1 vccd1 _7604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6109__328 _6110__329/A vssd1 vssd1 vccd1 vccd1 _7377_/CLK sky130_fd_sc_hd__inv_2
X_7827_ _7829_/CLK _7827_/D vssd1 vssd1 vccd1 vccd1 _7827_/Q sky130_fd_sc_hd__dfxtp_1
X_7758_ _7758_/CLK _7758_/D vssd1 vssd1 vccd1 vccd1 _7758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6709_ _6707_/X _6708_/X _6690_/X vssd1 vssd1 vccd1 vccd1 _7682_/D sky130_fd_sc_hd__a21oi_1
Xclkbuf_0__2768_ _5783_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2768_/X sky130_fd_sc_hd__clkbuf_16
X_7689_ _7689_/CLK _7689_/D vssd1 vssd1 vccd1 vccd1 _7689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5357__189 _5357__189/A vssd1 vssd1 vccd1 vccd1 _7161_/CLK sky130_fd_sc_hd__inv_2
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5040_/A _5044_/B vssd1 vssd1 vccd1 vccd1 _5041_/A sky130_fd_sc_hd__or2_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6991_ _6991_/A _6991_/B _6991_/C vssd1 vssd1 vccd1 vccd1 _6991_/X sky130_fd_sc_hd__and3_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5942_ _6011_/A vssd1 vssd1 vccd1 vccd1 _5942_/X sky130_fd_sc_hd__buf_4
XFILLER_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5873_ _5873_/A vssd1 vssd1 vccd1 vccd1 _7332_/D sky130_fd_sc_hd__clkbuf_1
X_6800__179 _6800__179/A vssd1 vssd1 vccd1 vccd1 _7746_/CLK sky130_fd_sc_hd__inv_2
XFILLER_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4824_ _4823_/X _7270_/Q _4827_/S vssd1 vssd1 vccd1 vccd1 _4825_/A sky130_fd_sc_hd__mux2_1
X_7612_ _7612_/CLK _7612_/D vssd1 vssd1 vccd1 vccd1 _7612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7543_ _7543_/CLK _7543_/D vssd1 vssd1 vccd1 vccd1 _7543_/Q sky130_fd_sc_hd__dfxtp_1
X_4755_ _4713_/X _7298_/Q _4759_/S vssd1 vssd1 vccd1 vccd1 _4756_/A sky130_fd_sc_hd__mux2_1
X_7896__223 vssd1 vssd1 vccd1 vccd1 _7896__223/HI partID[9] sky130_fd_sc_hd__conb_1
X_3706_ _3935_/A vssd1 vssd1 vccd1 vccd1 _3706_/X sky130_fd_sc_hd__clkbuf_2
X_7474_ _7474_/CLK _7474_/D vssd1 vssd1 vccd1 vccd1 _7474_/Q sky130_fd_sc_hd__dfxtp_1
X_4686_ _4686_/A _4865_/B vssd1 vssd1 vccd1 vccd1 _4847_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3637_ _3558_/X _7774_/Q _3641_/S vssd1 vssd1 vccd1 vccd1 _3638_/A sky130_fd_sc_hd__mux2_1
X_3568_ _3568_/A vssd1 vssd1 vccd1 vccd1 _7833_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3137_ clkbuf_0__3137_/X vssd1 vssd1 vccd1 vccd1 _6498__67/A sky130_fd_sc_hd__clkbuf_4
X_5307_ _5307_/A vssd1 vssd1 vccd1 vccd1 _5307_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3105_ _6336_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3105_/X sky130_fd_sc_hd__clkbuf_16
X_5238_ _5145_/X _7228_/Q _5682_/B _7203_/Q _5237_/X vssd1 vssd1 vccd1 vccd1 _5238_/X
+ sky130_fd_sc_hd__a221o_4
X_6412__479 _6412__479/A vssd1 vssd1 vccd1 vccd1 _7544_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5169_ _7191_/Q _5175_/B _5171_/C vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__and3_1
XFILLER_56_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6736__129 _6736__129/A vssd1 vssd1 vccd1 vccd1 _7695_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_wb_clk_i _7474_/CLK vssd1 vssd1 vccd1 vccd1 _7799_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4540_ _4540_/A vssd1 vssd1 vccd1 vccd1 _7424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4471_ _4393_/X _7456_/Q _4479_/S vssd1 vssd1 vccd1 vccd1 _4472_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7190_ _7839_/CLK _7190_/D vssd1 vssd1 vccd1 vccd1 _7190_/Q sky130_fd_sc_hd__dfxtp_1
X_6210_ _7799_/Q vssd1 vssd1 vccd1 vccd1 _6930_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _7625_/Q _7617_/Q _7609_/Q _7601_/Q _6024_/X _5998_/X vssd1 vssd1 vccd1 vccd1
+ _6072_/X sky130_fd_sc_hd__mux4_2
X_5023_ _5023_/A vssd1 vssd1 vccd1 vccd1 _5023_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_19 _5156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6974_ _6983_/A _6974_/B vssd1 vssd1 vccd1 vccd1 _6974_/Y sky130_fd_sc_hd__nor2_1
X_5925_ _5925_/A vssd1 vssd1 vccd1 vccd1 _5925_/X sky130_fd_sc_hd__buf_1
XFILLER_53_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5856_ _5856_/A _5892_/B vssd1 vssd1 vccd1 vccd1 _5872_/S sky130_fd_sc_hd__nand2_2
XFILLER_80_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4807_ _4807_/A vssd1 vssd1 vccd1 vccd1 _7276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7526_ _7526_/CLK _7526_/D vssd1 vssd1 vccd1 vccd1 _7526_/Q sky130_fd_sc_hd__dfxtp_1
X_4738_ _4738_/A vssd1 vssd1 vccd1 vccd1 _7306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4669_ _4684_/S vssd1 vssd1 vccd1 vccd1 _4678_/S sky130_fd_sc_hd__buf_2
X_7457_ _7457_/CLK _7457_/D vssd1 vssd1 vccd1 vccd1 _7457_/Q sky130_fd_sc_hd__dfxtp_1
X_7388_ _7388_/CLK _7388_/D vssd1 vssd1 vccd1 vccd1 _7388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6460__517 _6462__519/A vssd1 vssd1 vccd1 vccd1 _7582_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3971_ _3971_/A vssd1 vssd1 vccd1 vccd1 _7643_/D sky130_fd_sc_hd__clkbuf_1
X_5710_ _7216_/Q _5114_/A _5714_/S vssd1 vssd1 vccd1 vccd1 _5711_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6690_ _6690_/A vssd1 vssd1 vccd1 vccd1 _6690_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5641_ _5645_/A _5641_/B vssd1 vssd1 vccd1 vccd1 _5642_/A sky130_fd_sc_hd__or2_1
X_5572_ _5570_/X _5571_/X _5572_/S vssd1 vssd1 vccd1 vccd1 _5572_/X sky130_fd_sc_hd__mux2_1
X_4523_ _4632_/A _4523_/B vssd1 vssd1 vccd1 vccd1 _4539_/S sky130_fd_sc_hd__nand2_2
X_7311_ _7311_/CLK _7311_/D vssd1 vssd1 vccd1 vccd1 _7311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7242_ _7242_/CLK _7242_/D vssd1 vssd1 vccd1 vccd1 _7242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4454_ _4436_/X _4455_/B _4453_/Y vssd1 vssd1 vccd1 vccd1 _7461_/D sky130_fd_sc_hd__o21a_1
X_4385_ _7489_/Q _3941_/A _4385_/S vssd1 vssd1 vccd1 vccd1 _4386_/A sky130_fd_sc_hd__mux2_1
X_7173_ _7173_/CLK _7173_/D vssd1 vssd1 vccd1 vccd1 _7173_/Q sky130_fd_sc_hd__dfxtp_1
X_6124_ _6130_/A vssd1 vssd1 vccd1 vccd1 _6124_/X sky130_fd_sc_hd__buf_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6055_ _7369_/Q _5931_/X _6054_/X _5996_/X vssd1 vssd1 vccd1 vccd1 _7369_/D sky130_fd_sc_hd__o211a_1
XFILLER_85_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _5874_/A _5087_/B vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__and2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6957_ _7806_/Q _6969_/B vssd1 vssd1 vccd1 vccd1 _6957_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3121_ clkbuf_0__3121_/X vssd1 vssd1 vccd1 vccd1 _6444_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5908_ _7348_/Q _5081_/A _5908_/S vssd1 vssd1 vccd1 vccd1 _5909_/A sky130_fd_sc_hd__mux2_1
X_6888_ _7841_/Q _6888_/B vssd1 vssd1 vccd1 vccd1 _6892_/B sky130_fd_sc_hd__xor2_1
XFILLER_14_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7509_ _7509_/CLK _7509_/D vssd1 vssd1 vccd1 vccd1 _7509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2767_ clkbuf_0__2767_/X vssd1 vssd1 vccd1 vccd1 _5782__249/A sky130_fd_sc_hd__clkbuf_4
XFILLER_45_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6384__459 _6384__459/A vssd1 vssd1 vccd1 vccd1 _7522_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6425__489 _6425__489/A vssd1 vssd1 vccd1 vccd1 _7554_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4170_ _4414_/A vssd1 vssd1 vccd1 vccd1 _4170_/X sky130_fd_sc_hd__buf_2
XFILLER_96_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6541__102 _6543__104/A vssd1 vssd1 vccd1 vccd1 _7647_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7791_ _7791_/CLK _7791_/D vssd1 vssd1 vccd1 vccd1 _7791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3954_ _4668_/A _4632_/B vssd1 vssd1 vccd1 vccd1 _3970_/S sky130_fd_sc_hd__nand2_2
X_6673_ _6677_/A _6714_/C _6600_/B vssd1 vssd1 vccd1 vccd1 _6673_/X sky130_fd_sc_hd__or3b_1
X_3885_ _3885_/A vssd1 vssd1 vccd1 vccd1 _7697_/D sky130_fd_sc_hd__clkbuf_1
X_5745__219 _5745__219/A vssd1 vssd1 vccd1 vccd1 _7236_/CLK sky130_fd_sc_hd__inv_2
X_5624_ _5613_/A _5621_/X _5623_/X vssd1 vssd1 vccd1 vccd1 _5624_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5555_ _7514_/Q _7506_/Q _7445_/Q _7437_/Q _5512_/X _5506_/X vssd1 vssd1 vccd1 vccd1
+ _5555_/X sky130_fd_sc_hd__mux4_2
XFILLER_117_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4506_ _4521_/S vssd1 vssd1 vccd1 vccd1 _4515_/S sky130_fd_sc_hd__buf_2
X_5486_ _5518_/A vssd1 vssd1 vccd1 vccd1 _5486_/X sky130_fd_sc_hd__clkbuf_8
X_7225_ _7333_/CLK _7225_/D vssd1 vssd1 vccd1 vccd1 _7225_/Q sky130_fd_sc_hd__dfxtp_1
X_4437_ _7460_/Q vssd1 vssd1 vccd1 vccd1 _4452_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7156_ _7331_/CLK _7156_/D vssd1 vssd1 vccd1 vccd1 _7156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ _4368_/A vssd1 vssd1 vccd1 vccd1 _7497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7087_ _7087_/A vssd1 vssd1 vccd1 vccd1 _7850_/D sky130_fd_sc_hd__clkbuf_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _4301_/A vssd1 vssd1 vccd1 vccd1 _4300_/A sky130_fd_sc_hd__buf_6
XFILLER_100_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6038_ _5932_/X _6026_/X _6037_/X _5993_/X vssd1 vssd1 vccd1 vccd1 _6038_/X sky130_fd_sc_hd__a211o_2
XFILLER_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3104_ clkbuf_0__3104_/X vssd1 vssd1 vccd1 vccd1 _6335__419/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6390__463 _6391__464/A vssd1 vssd1 vccd1 vccd1 _7526_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5850__303 _5851__304/A vssd1 vssd1 vccd1 vccd1 _7320_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3670_ _7763_/Q _3669_/X _3676_/S vssd1 vssd1 vccd1 vccd1 _3671_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput105 _5128_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[20] sky130_fd_sc_hd__buf_2
Xoutput116 _5095_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[5] sky130_fd_sc_hd__buf_2
X_5340_ _5187_/X _5682_/C _7228_/D vssd1 vssd1 vccd1 vccd1 _5343_/A sky130_fd_sc_hd__a21oi_2
XFILLER_99_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput138 _5067_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[24] sky130_fd_sc_hd__buf_2
Xoutput127 _5045_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[14] sky130_fd_sc_hd__buf_2
Xoutput149 _5026_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_114_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5271_ _5270_/X _7151_/Q _5262_/X _5266_/X _7119_/Q vssd1 vssd1 vccd1 vccd1 _7119_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4222_ _7545_/Q _4221_/X _4231_/S vssd1 vssd1 vccd1 vccd1 _4223_/A sky130_fd_sc_hd__mux2_1
X_7010_ _7820_/Q _7013_/S _7009_/X _7003_/X vssd1 vssd1 vccd1 vccd1 _7819_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4153_ _4149_/X _7570_/Q _4165_/S vssd1 vssd1 vccd1 vccd1 _4154_/A sky130_fd_sc_hd__mux2_1
X_4084_ _4063_/X _7597_/Q _4088_/S vssd1 vssd1 vccd1 vccd1 _4085_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7843_ _7845_/CLK _7843_/D vssd1 vssd1 vccd1 vccd1 _7843_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7774_ _7774_/CLK _7774_/D vssd1 vssd1 vccd1 vccd1 _7774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4986_ _4986_/A vssd1 vssd1 vccd1 vccd1 _7110_/D sky130_fd_sc_hd__clkbuf_1
X_3937_ _3937_/A vssd1 vssd1 vccd1 vccd1 _7656_/D sky130_fd_sc_hd__clkbuf_1
X_6725_ _7687_/Q _6725_/B _6725_/C _6725_/D vssd1 vssd1 vccd1 vccd1 _6726_/C sky130_fd_sc_hd__and4b_1
XFILLER_32_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6656_ _6679_/A vssd1 vssd1 vccd1 vccd1 _6656_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3868_ _4901_/A _4901_/B _4731_/C _4955_/A vssd1 vssd1 vccd1 vccd1 _3884_/S sky130_fd_sc_hd__or4_4
X_6587_ _7851_/Q _6677_/B vssd1 vssd1 vccd1 vccd1 _6588_/D sky130_fd_sc_hd__xor2_1
X_5607_ _5455_/X _5604_/X _5606_/X vssd1 vssd1 vccd1 vccd1 _7190_/D sky130_fd_sc_hd__a21o_1
X_3799_ _3794_/X _4303_/B _3791_/B _4303_/D vssd1 vssd1 vccd1 vccd1 _3800_/B sky130_fd_sc_hd__o22a_1
X_5538_ _5536_/X _5537_/X _5575_/S vssd1 vssd1 vccd1 vccd1 _5538_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3299_ clkbuf_0__3299_/X vssd1 vssd1 vccd1 vccd1 _6769__154/A sky130_fd_sc_hd__clkbuf_4
X_7208_ _7477_/CLK _7208_/D vssd1 vssd1 vccd1 vccd1 _7208_/Q sky130_fd_sc_hd__dfxtp_1
X_5469_ _5466_/X _5468_/X _5403_/A vssd1 vssd1 vccd1 vccd1 _5469_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7139_ _7339_/CLK _7139_/D vssd1 vssd1 vccd1 vccd1 _7139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 caravel_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 _5218_/B sky130_fd_sc_hd__clkbuf_1
Xinput29 caravel_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_2
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6275__389 _6275__389/A vssd1 vssd1 vccd1 vccd1 _7442_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5815__275 _5819__279/A vssd1 vssd1 vccd1 vccd1 _7292_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4840_ _4840_/A vssd1 vssd1 vccd1 vccd1 _7264_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _4710_/X _7291_/Q _4777_/S vssd1 vssd1 vccd1 vccd1 _4772_/A sky130_fd_sc_hd__mux2_1
X_7490_ _7490_/CLK _7490_/D vssd1 vssd1 vccd1 vccd1 _7490_/Q sky130_fd_sc_hd__dfxtp_1
X_3722_ _3721_/X _7745_/Q _3722_/S vssd1 vssd1 vccd1 vccd1 _3723_/A sky130_fd_sc_hd__mux2_1
X_3653_ _4578_/A _3653_/B _4431_/B vssd1 vssd1 vccd1 vccd1 _3676_/S sky130_fd_sc_hd__and3_2
XFILLER_9_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5323_ _5323_/A vssd1 vssd1 vccd1 vccd1 _7150_/D sky130_fd_sc_hd__clkbuf_1
X_3584_ _4614_/A _4614_/B _4614_/C vssd1 vssd1 vccd1 vccd1 _3653_/B sky130_fd_sc_hd__and3b_2
Xclkbuf_1_1_0__3084_ clkbuf_0__3084_/X vssd1 vssd1 vccd1 vccd1 _6275__389/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3121_ _6419_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3121_/X sky130_fd_sc_hd__clkbuf_16
X_5185_ _7197_/Q _5189_/B _5185_/C vssd1 vssd1 vccd1 vccd1 _5185_/X sky130_fd_sc_hd__and3_1
X_4205_ _4164_/X _7550_/Q _4205_/S vssd1 vssd1 vccd1 vccd1 _4206_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4136_ _4136_/A vssd1 vssd1 vccd1 vccd1 _7577_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4067_ _4066_/X _7604_/Q _4070_/S vssd1 vssd1 vccd1 vccd1 _4068_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7826_ _7826_/CLK _7826_/D vssd1 vssd1 vccd1 vccd1 _7826_/Q sky130_fd_sc_hd__dfxtp_2
X_6341__424 _6341__424/A vssd1 vssd1 vccd1 vccd1 _7487_/CLK sky130_fd_sc_hd__inv_2
X_7757_ _7757_/CLK _7757_/D vssd1 vssd1 vccd1 vccd1 _7757_/Q sky130_fd_sc_hd__dfxtp_1
X_4969_ _4236_/X _7161_/Q _4971_/S vssd1 vssd1 vccd1 vccd1 _4970_/A sky130_fd_sc_hd__mux2_1
X_6708_ _6708_/A _6708_/B _6714_/C vssd1 vssd1 vccd1 vccd1 _6708_/X sky130_fd_sc_hd__or3_1
Xclkbuf_0__2767_ _5777_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2767_/X sky130_fd_sc_hd__clkbuf_16
X_7688_ _7688_/CLK _7688_/D vssd1 vssd1 vccd1 vccd1 _7688_/Q sky130_fd_sc_hd__dfxtp_1
X_6554__112 _6555__113/A vssd1 vssd1 vccd1 vccd1 _7657_/CLK sky130_fd_sc_hd__inv_2
X_6639_ _6679_/A vssd1 vssd1 vccd1 vccd1 _6640_/C sky130_fd_sc_hd__buf_2
XFILLER_22_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2449_ clkbuf_0__2449_/X vssd1 vssd1 vccd1 vccd1 _5374__203/A sky130_fd_sc_hd__clkbuf_4
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6990_ _6213_/Y _6214_/X _6866_/B _6989_/X _6866_/A vssd1 vssd1 vccd1 vccd1 _6993_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5941_ _7619_/Q _7611_/Q _7603_/Q _7595_/Q _5939_/X _5940_/X vssd1 vssd1 vccd1 vccd1
+ _5941_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5872_ _5047_/A _7332_/Q _5872_/S vssd1 vssd1 vccd1 vccd1 _5873_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6479__533 _6480__534/A vssd1 vssd1 vccd1 vccd1 _7598_/CLK sky130_fd_sc_hd__inv_2
X_4823_ _7469_/Q vssd1 vssd1 vccd1 vccd1 _4823_/X sky130_fd_sc_hd__buf_2
X_7611_ _7611_/CLK _7611_/D vssd1 vssd1 vccd1 vccd1 _7611_/Q sky130_fd_sc_hd__dfxtp_1
X_7542_ _7542_/CLK _7542_/D vssd1 vssd1 vccd1 vccd1 _7542_/Q sky130_fd_sc_hd__dfxtp_1
X_4754_ _4754_/A vssd1 vssd1 vccd1 vccd1 _7299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3705_ _3705_/A vssd1 vssd1 vccd1 vccd1 _7751_/D sky130_fd_sc_hd__clkbuf_1
X_7473_ _7473_/CLK _7473_/D vssd1 vssd1 vccd1 vccd1 _7473_/Q sky130_fd_sc_hd__dfxtp_1
X_4685_ _4685_/A vssd1 vssd1 vccd1 vccd1 _7349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3636_ _3636_/A vssd1 vssd1 vccd1 vccd1 _7775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3567_ _3566_/X _7833_/Q _3567_/S vssd1 vssd1 vccd1 vccd1 _3568_/A sky130_fd_sc_hd__mux2_1
X_6355_ _6379_/A vssd1 vssd1 vccd1 vccd1 _6355_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3136_ clkbuf_0__3136_/X vssd1 vssd1 vccd1 vccd1 _6494__64/A sky130_fd_sc_hd__clkbuf_4
X_5306_ _5303_/X _7341_/Q _5299_/X _5300_/X _7141_/Q vssd1 vssd1 vccd1 vccd1 _7141_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6768__153 _6768__153/A vssd1 vssd1 vccd1 vccd1 _7720_/CLK sky130_fd_sc_hd__inv_2
X_5237_ input35/X input2/X _5138_/D vssd1 vssd1 vccd1 vccd1 _5237_/X sky130_fd_sc_hd__o21a_4
XFILLER_115_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3104_ _6330_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3104_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_102_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6115__333 _6116__334/A vssd1 vssd1 vccd1 vccd1 _7382_/CLK sky130_fd_sc_hd__inv_2
X_5168_ _7123_/Q _5159_/X input31/X _5163_/X _5167_/X vssd1 vssd1 vccd1 vccd1 _5168_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_84_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5099_ _5099_/A vssd1 vssd1 vccd1 vccd1 _5099_/X sky130_fd_sc_hd__clkbuf_1
X_4119_ _3820_/X _7584_/Q _4123_/S vssd1 vssd1 vccd1 vccd1 _4120_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7809_ _7812_/CLK _7809_/D vssd1 vssd1 vccd1 vccd1 _7809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__2998_ clkbuf_0__2998_/X vssd1 vssd1 vccd1 vccd1 _6178__379/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5363__194 _5363__194/A vssd1 vssd1 vccd1 vccd1 _7166_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5927__321 _5929__323/A vssd1 vssd1 vccd1 vccd1 _7362_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4470_ _4485_/S vssd1 vssd1 vccd1 vccd1 _4479_/S sky130_fd_sc_hd__buf_2
X_7856__230 vssd1 vssd1 vccd1 vccd1 core1Index[0] _7856__230/LO sky130_fd_sc_hd__conb_1
XFILLER_112_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _7370_/Q _6631_/B _6070_/X _5996_/X vssd1 vssd1 vccd1 vccd1 _7370_/D sky130_fd_sc_hd__o211a_1
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _7024_/A _5022_/B vssd1 vssd1 vccd1 vccd1 _5023_/A sky130_fd_sc_hd__or2_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6973_ _6969_/Y _6972_/X _6954_/A vssd1 vssd1 vccd1 vccd1 _7810_/D sky130_fd_sc_hd__a21oi_1
XFILLER_81_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4806_ _4803_/X _7276_/Q _4818_/S vssd1 vssd1 vccd1 vccd1 _4807_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7525_ _7525_/CLK _7525_/D vssd1 vssd1 vccd1 vccd1 _7525_/Q sky130_fd_sc_hd__dfxtp_1
X_4737_ _4713_/X _7306_/Q _4741_/S vssd1 vssd1 vccd1 vccd1 _4738_/A sky130_fd_sc_hd__mux2_1
X_4668_ _4668_/A _4668_/B vssd1 vssd1 vccd1 vccd1 _4684_/S sky130_fd_sc_hd__nand2_2
X_7456_ _7456_/CLK _7456_/D vssd1 vssd1 vccd1 vccd1 _7456_/Q sky130_fd_sc_hd__dfxtp_1
X_3619_ _3619_/A vssd1 vssd1 vccd1 vccd1 _7782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6407_ _6413_/A vssd1 vssd1 vccd1 vccd1 _6407_/X sky130_fd_sc_hd__buf_1
X_4599_ _4599_/A vssd1 vssd1 vccd1 vccd1 _7396_/D sky130_fd_sc_hd__clkbuf_1
X_7387_ _7387_/CLK _7387_/D vssd1 vssd1 vccd1 vccd1 _7387_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3119_ clkbuf_0__3119_/X vssd1 vssd1 vccd1 vccd1 _6409__476/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6269_ _6269_/A vssd1 vssd1 vccd1 vccd1 _6269_/X sky130_fd_sc_hd__buf_1
XFILLER_0_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5794__259 _5794__259/A vssd1 vssd1 vccd1 vccd1 _7276_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3970_ _3950_/X _7643_/Q _3970_/S vssd1 vssd1 vccd1 vccd1 _3971_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5640_ _7846_/Q _5672_/D _5638_/X _7193_/Q _5639_/X vssd1 vssd1 vccd1 vccd1 _5641_/B
+ sky130_fd_sc_hd__a32o_1
X_5571_ _7693_/Q _7282_/Q _7165_/Q _7274_/Q _5472_/A _5508_/X vssd1 vssd1 vccd1 vccd1
+ _5571_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7310_ _7310_/CLK _7310_/D vssd1 vssd1 vccd1 vccd1 _7310_/Q sky130_fd_sc_hd__dfxtp_1
X_4522_ _4522_/A vssd1 vssd1 vccd1 vccd1 _7433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4453_ _4436_/X _4455_/B _6325_/A vssd1 vssd1 vccd1 vccd1 _4453_/Y sky130_fd_sc_hd__a21oi_1
X_7241_ _7241_/CLK _7241_/D vssd1 vssd1 vccd1 vccd1 _7241_/Q sky130_fd_sc_hd__dfxtp_1
X_4384_ _4384_/A vssd1 vssd1 vccd1 vccd1 _7490_/D sky130_fd_sc_hd__clkbuf_1
X_7172_ _7172_/CLK _7172_/D vssd1 vssd1 vccd1 vccd1 _7172_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6054_ _5932_/X _6044_/X _6053_/X _5993_/X vssd1 vssd1 vccd1 vccd1 _6054_/X sky130_fd_sc_hd__a211o_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5142_/B vssd1 vssd1 vccd1 vccd1 _5087_/B sky130_fd_sc_hd__clkbuf_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6811__12 _6812__13/A vssd1 vssd1 vccd1 vccd1 _7754_/CLK sky130_fd_sc_hd__inv_2
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6956_ _6972_/B vssd1 vssd1 vccd1 vccd1 _6969_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0_0__3120_ clkbuf_0__3120_/X vssd1 vssd1 vccd1 vccd1 _6418__484/A sky130_fd_sc_hd__clkbuf_4
X_5907_ _5907_/A vssd1 vssd1 vccd1 vccd1 _7347_/D sky130_fd_sc_hd__clkbuf_1
X_6887_ _6887_/A _6887_/B _6887_/C vssd1 vssd1 vccd1 vccd1 _6893_/C sky130_fd_sc_hd__or3_1
XFILLER_14_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7508_ _7508_/CLK _7508_/D vssd1 vssd1 vccd1 vccd1 _7508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7439_ _7439_/CLK _7439_/D vssd1 vssd1 vccd1 vccd1 _7439_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2449_ _5370_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2449_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_115_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6128__343 _6129__344/A vssd1 vssd1 vccd1 vccd1 _7392_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6645__116 _6645__116/A vssd1 vssd1 vccd1 vccd1 _7663_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7790_ _7790_/CLK _7790_/D vssd1 vssd1 vccd1 vccd1 _7790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3953_ _4614_/A _4614_/B _4614_/C vssd1 vssd1 vccd1 vccd1 _4632_/B sky130_fd_sc_hd__and3_2
XFILLER_51_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6672_ _6640_/C _6661_/X _6598_/Y vssd1 vssd1 vccd1 vccd1 _6672_/X sky130_fd_sc_hd__a21o_1
X_3884_ _3840_/X _7697_/Q _3884_/S vssd1 vssd1 vccd1 vccd1 _3885_/A sky130_fd_sc_hd__mux2_1
X_5623_ _5466_/X _5622_/X _5404_/A vssd1 vssd1 vccd1 vccd1 _5623_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5554_ _7241_/Q _7172_/Q _7482_/Q _7249_/Q _5479_/X _5508_/X vssd1 vssd1 vccd1 vccd1
+ _5554_/X sky130_fd_sc_hd__mux4_1
X_5485_ _5611_/S _5485_/B vssd1 vssd1 vccd1 vccd1 _5485_/X sky130_fd_sc_hd__and2_1
X_4505_ _4865_/A _4865_/B _4505_/C vssd1 vssd1 vccd1 vccd1 _4521_/S sky130_fd_sc_hd__and3_2
X_7224_ _7224_/CLK _7224_/D vssd1 vssd1 vccd1 vccd1 _7224_/Q sky130_fd_sc_hd__dfxtp_1
X_4436_ _5964_/A vssd1 vssd1 vccd1 vccd1 _4436_/X sky130_fd_sc_hd__buf_2
X_7155_ _7331_/CLK _7155_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
X_4367_ _4164_/X _7497_/Q _4367_/S vssd1 vssd1 vccd1 vccd1 _4368_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7086_ _7070_/X _7086_/B vssd1 vssd1 vccd1 vccd1 _7087_/A sky130_fd_sc_hd__and2b_1
XFILLER_58_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _7518_/Q vssd1 vssd1 vccd1 vccd1 _4301_/A sky130_fd_sc_hd__buf_4
X_6037_ _6030_/X _6035_/X _6036_/X vssd1 vssd1 vccd1 vccd1 _6037_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2998_ _6173_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2998_/X sky130_fd_sc_hd__clkbuf_16
X_6939_ _6939_/A vssd1 vssd1 vccd1 vccd1 _6939_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6431__494 _6431__494/A vssd1 vssd1 vccd1 vccd1 _7559_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6473__528 _6474__529/A vssd1 vssd1 vccd1 vccd1 _7593_/CLK sky130_fd_sc_hd__inv_2
Xoutput106 _5130_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[21] sky130_fd_sc_hd__buf_2
Xoutput139 _5070_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[25] sky130_fd_sc_hd__buf_2
Xoutput128 _5048_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[15] sky130_fd_sc_hd__buf_2
Xoutput117 _5097_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[6] sky130_fd_sc_hd__buf_2
X_5270_ _5303_/A vssd1 vssd1 vccd1 vccd1 _5270_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4221_ _7474_/Q vssd1 vssd1 vccd1 vccd1 _4221_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4152_ _4174_/S vssd1 vssd1 vccd1 vccd1 _4165_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4083_ _4083_/A vssd1 vssd1 vccd1 vccd1 _7598_/D sky130_fd_sc_hd__clkbuf_1
X_6762__148 _6763__149/A vssd1 vssd1 vccd1 vccd1 _7715_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5751__224 _5751__224/A vssd1 vssd1 vccd1 vccd1 _7241_/CLK sky130_fd_sc_hd__inv_2
X_7842_ _7845_/CLK _7842_/D vssd1 vssd1 vccd1 vccd1 _7842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7773_ _7773_/CLK _7773_/D vssd1 vssd1 vccd1 vccd1 _7773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4985_ _7110_/Q _4414_/A _4987_/S vssd1 vssd1 vccd1 vccd1 _4986_/A sky130_fd_sc_hd__mux2_1
X_3936_ _3935_/X _7656_/Q _3942_/S vssd1 vssd1 vccd1 vccd1 _3937_/A sky130_fd_sc_hd__mux2_1
X_6724_ _6724_/A vssd1 vssd1 vccd1 vccd1 _7686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6655_ _6705_/D vssd1 vssd1 vccd1 vccd1 _6711_/D sky130_fd_sc_hd__clkbuf_2
X_3867_ _4194_/A _4280_/A _4286_/B vssd1 vssd1 vccd1 vccd1 _4955_/A sky130_fd_sc_hd__or3_2
X_6586_ _7673_/Q _6621_/B vssd1 vssd1 vccd1 vccd1 _6677_/B sky130_fd_sc_hd__xnor2_1
X_5606_ _7190_/Q _5453_/A _5680_/A vssd1 vssd1 vccd1 vccd1 _5606_/X sky130_fd_sc_hd__a21o_1
X_3798_ _7526_/Q _7521_/Q vssd1 vssd1 vccd1 vccd1 _4303_/D sky130_fd_sc_hd__xnor2_1
XFILLER_11_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5537_ _7513_/Q _7505_/Q _7444_/Q _7436_/Q _5512_/X _5513_/X vssd1 vssd1 vccd1 vccd1
+ _5537_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_1_1_0__3298_ clkbuf_0__3298_/X vssd1 vssd1 vccd1 vccd1 _6760__146/A sky130_fd_sc_hd__clkbuf_4
X_7207_ _7477_/CLK _7207_/D vssd1 vssd1 vccd1 vccd1 _7207_/Q sky130_fd_sc_hd__dfxtp_1
X_5468_ _7177_/Q _7358_/Q _7714_/Q _7254_/Q _4301_/A _5467_/X vssd1 vssd1 vccd1 vccd1
+ _5468_/X sky130_fd_sc_hd__mux4_2
X_5399_ _7224_/Q _5493_/A _5399_/C _5399_/D vssd1 vssd1 vccd1 vccd1 _5401_/C sky130_fd_sc_hd__or4_4
XFILLER_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4419_ _4419_/A vssd1 vssd1 vccd1 vccd1 _7478_/D sky130_fd_sc_hd__clkbuf_1
X_7138_ _7339_/CLK _7138_/D vssd1 vssd1 vccd1 vccd1 _7138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7069_ _7069_/A vssd1 vssd1 vccd1 vccd1 _7845_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7838_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput19 caravel_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 _5220_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_10_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5921__316 _5924__319/A vssd1 vssd1 vccd1 vccd1 _7357_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4770_ _4770_/A vssd1 vssd1 vccd1 vccd1 _7292_/D sky130_fd_sc_hd__clkbuf_1
X_3721_ _3950_/A vssd1 vssd1 vccd1 vccd1 _3721_/X sky130_fd_sc_hd__clkbuf_2
X_3652_ _4578_/B vssd1 vssd1 vccd1 vccd1 _4431_/B sky130_fd_sc_hd__clkbuf_2
X_3583_ _7464_/Q vssd1 vssd1 vccd1 vccd1 _4614_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5322_ _7100_/A _7150_/Q _5328_/S vssd1 vssd1 vccd1 vccd1 _5323_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3083_ clkbuf_0__3083_/X vssd1 vssd1 vccd1 vccd1 _6294_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3120_ _6413_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3120_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_88_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5184_ _7129_/Q _5173_/X input6/X _5177_/X _5183_/X vssd1 vssd1 vccd1 vccd1 _5184_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_68_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4204_ _4204_/A vssd1 vssd1 vccd1 vccd1 _7551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4135_ _4051_/X _7577_/Q _4141_/S vssd1 vssd1 vccd1 vccd1 _4136_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4066_ _7823_/Q vssd1 vssd1 vccd1 vccd1 _4066_/X sky130_fd_sc_hd__buf_2
X_7825_ _7825_/CLK _7825_/D vssd1 vssd1 vccd1 vccd1 _7825_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7756_ _7756_/CLK _7756_/D vssd1 vssd1 vccd1 vccd1 _7756_/Q sky130_fd_sc_hd__dfxtp_1
X_4968_ _4968_/A vssd1 vssd1 vccd1 vccd1 _7162_/D sky130_fd_sc_hd__clkbuf_1
X_7687_ _7687_/CLK _7687_/D vssd1 vssd1 vccd1 vccd1 _7687_/Q sky130_fd_sc_hd__dfxtp_1
X_6707_ _6679_/X _6684_/X _7682_/Q vssd1 vssd1 vccd1 vccd1 _6707_/X sky130_fd_sc_hd__a21bo_1
X_3919_ _3919_/A vssd1 vssd1 vccd1 vccd1 _7664_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__2766_ _5771_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2766_/X sky130_fd_sc_hd__clkbuf_16
X_4899_ _4826_/X _7237_/Q _4899_/S vssd1 vssd1 vccd1 vccd1 _4900_/A sky130_fd_sc_hd__mux2_1
X_6638_ _5951_/A _6630_/X _6637_/A _6725_/C vssd1 vssd1 vccd1 vccd1 _6679_/A sky130_fd_sc_hd__a211o_2
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6569_ _6569_/A vssd1 vssd1 vccd1 vccd1 _6613_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2448_ clkbuf_0__2448_/X vssd1 vssd1 vccd1 vccd1 _5369__199/A sky130_fd_sc_hd__clkbuf_4
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7880__207 vssd1 vssd1 vccd1 vccd1 _7880__207/HI core1Index[7] sky130_fd_sc_hd__conb_1
XFILLER_70_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6281__394 _6281__394/A vssd1 vssd1 vccd1 vccd1 _7447_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5821__280 _5824__283/A vssd1 vssd1 vccd1 vccd1 _7297_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5940_ _5998_/A vssd1 vssd1 vccd1 vccd1 _5940_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5871_ _5871_/A vssd1 vssd1 vccd1 vccd1 _7331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7610_ _7610_/CLK _7610_/D vssd1 vssd1 vccd1 vccd1 _7610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4822_ _4822_/A vssd1 vssd1 vccd1 vccd1 _7271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4753_ _4710_/X _7299_/Q _4759_/S vssd1 vssd1 vccd1 vccd1 _4754_/A sky130_fd_sc_hd__mux2_1
X_7541_ _7541_/CLK _7541_/D vssd1 vssd1 vccd1 vccd1 _7541_/Q sky130_fd_sc_hd__dfxtp_1
X_3704_ _3703_/X _7751_/Q _3713_/S vssd1 vssd1 vccd1 vccd1 _3705_/A sky130_fd_sc_hd__mux2_1
X_7472_ _7473_/CLK _7472_/D vssd1 vssd1 vccd1 vccd1 _7472_/Q sky130_fd_sc_hd__dfxtp_1
X_4684_ _3675_/X _7349_/Q _4684_/S vssd1 vssd1 vccd1 vccd1 _4685_/A sky130_fd_sc_hd__mux2_1
X_3635_ _3554_/X _7775_/Q _3641_/S vssd1 vssd1 vccd1 vccd1 _3636_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3566_ _3941_/A vssd1 vssd1 vccd1 vccd1 _3566_/X sky130_fd_sc_hd__clkbuf_4
X_6354_ _6385_/A vssd1 vssd1 vccd1 vccd1 _6354_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3135_ clkbuf_0__3135_/X vssd1 vssd1 vccd1 vccd1 _6488__59/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5305_ _5303_/X _7340_/Q _5299_/X _5300_/X _7140_/Q vssd1 vssd1 vccd1 vccd1 _7140_/D
+ sky130_fd_sc_hd__o32a_1
X_6818__18 _6818__18/A vssd1 vssd1 vccd1 vccd1 _7760_/CLK sky130_fd_sc_hd__inv_2
X_5236_ _7108_/Q _5236_/B vssd1 vssd1 vccd1 vccd1 _5682_/B sky130_fd_sc_hd__and2_1
XFILLER_69_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5167_ _7190_/Q _5175_/B _5171_/C vssd1 vssd1 vccd1 vccd1 _5167_/X sky130_fd_sc_hd__and3_1
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5098_ _5098_/A _5098_/B vssd1 vssd1 vccd1 vccd1 _5099_/A sky130_fd_sc_hd__and2_1
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4118_ _4118_/A vssd1 vssd1 vccd1 vccd1 _7585_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4049_ _4046_/X _7610_/Q _4061_/S vssd1 vssd1 vccd1 vccd1 _4050_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6775__158 _6776__159/A vssd1 vssd1 vccd1 vccd1 _7725_/CLK sky130_fd_sc_hd__inv_2
X_7808_ _7808_/CLK _7808_/D vssd1 vssd1 vccd1 vccd1 _7808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7739_ _7739_/CLK _7739_/D vssd1 vssd1 vccd1 vccd1 _7739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6122__338 _6122__338/A vssd1 vssd1 vccd1 vccd1 _7387_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2997_ clkbuf_0__2997_/X vssd1 vssd1 vccd1 vccd1 _6172__374/A sky130_fd_sc_hd__clkbuf_4
XFILLER_4_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6070_ _5932_/A _6060_/X _6069_/X _5993_/X vssd1 vssd1 vccd1 vccd1 _6070_/X sky130_fd_sc_hd__a211o_2
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5021_/A vssd1 vssd1 vccd1 vccd1 _5021_/X sky130_fd_sc_hd__clkbuf_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6972_ _6972_/A _6972_/B _6974_/B vssd1 vssd1 vccd1 vccd1 _6972_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4805_ _4827_/S vssd1 vssd1 vccd1 vccd1 _4818_/S sky130_fd_sc_hd__buf_2
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7524_ _7524_/CLK _7524_/D vssd1 vssd1 vccd1 vccd1 _7524_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4736_ _4736_/A vssd1 vssd1 vccd1 vccd1 _7307_/D sky130_fd_sc_hd__clkbuf_1
X_7455_ _7455_/CLK _7455_/D vssd1 vssd1 vccd1 vccd1 _7455_/Q sky130_fd_sc_hd__dfxtp_1
X_4667_ _4667_/A vssd1 vssd1 vccd1 vccd1 _7357_/D sky130_fd_sc_hd__clkbuf_1
X_3618_ _3558_/X _7782_/Q _3622_/S vssd1 vssd1 vccd1 vccd1 _3619_/A sky130_fd_sc_hd__mux2_1
X_7386_ _7386_/CLK _7386_/D vssd1 vssd1 vccd1 vccd1 _7386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4598_ _4242_/X _7396_/Q _4606_/S vssd1 vssd1 vccd1 vccd1 _4599_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3118_ clkbuf_0__3118_/X vssd1 vssd1 vccd1 vccd1 _6404__472/A sky130_fd_sc_hd__clkbuf_4
X_3549_ _4243_/A _4028_/A vssd1 vssd1 vccd1 vccd1 _3579_/S sky130_fd_sc_hd__or2_2
Xclkbuf_1_0_0__2782_ clkbuf_0__2782_/X vssd1 vssd1 vccd1 vccd1 _5855__307/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5219_ _7140_/Q _5215_/X _5216_/X _5218_/X vssd1 vssd1 vccd1 vccd1 _5219_/X sky130_fd_sc_hd__o22a_4
XFILLER_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6199_ _6228_/B vssd1 vssd1 vccd1 vccd1 _6233_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7886__213 vssd1 vssd1 vccd1 vccd1 _7886__213/HI manufacturerID[5] sky130_fd_sc_hd__conb_1
XFILLER_85_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5570_ _7298_/Q _7290_/Q _7266_/Q _7114_/Q _4301_/A _5467_/X vssd1 vssd1 vccd1 vccd1
+ _5570_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4521_ _7433_/Q _4239_/X _4521_/S vssd1 vssd1 vccd1 vccd1 _4522_/A sky130_fd_sc_hd__mux2_1
X_4452_ _4452_/A _4459_/A vssd1 vssd1 vccd1 vccd1 _4455_/B sky130_fd_sc_hd__and2_1
X_7240_ _7240_/CLK _7240_/D vssd1 vssd1 vccd1 vccd1 _7240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4383_ _7490_/Q _3938_/A _4385_/S vssd1 vssd1 vccd1 vccd1 _4384_/A sky130_fd_sc_hd__mux2_1
X_7171_ _7171_/CLK _7171_/D vssd1 vssd1 vccd1 vccd1 _7171_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6048_/X _6052_/X _6036_/X vssd1 vssd1 vccd1 vccd1 _6053_/X sky130_fd_sc_hd__o21a_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5004_/A vssd1 vssd1 vccd1 vccd1 _5142_/B sky130_fd_sc_hd__buf_2
XFILLER_85_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _6952_/Y _6953_/X _6954_/X vssd1 vssd1 vccd1 vccd1 _7805_/D sky130_fd_sc_hd__a21oi_1
XFILLER_26_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5906_ _7347_/Q _5079_/A _5908_/S vssd1 vssd1 vccd1 vccd1 _5907_/A sky130_fd_sc_hd__mux2_1
X_6886_ _7842_/Q _6194_/A _6232_/A _7847_/Q vssd1 vssd1 vccd1 vccd1 _6887_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4719_ _7471_/Q vssd1 vssd1 vccd1 vccd1 _4719_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7507_ _7507_/CLK _7507_/D vssd1 vssd1 vccd1 vccd1 _7507_/Q sky130_fd_sc_hd__dfxtp_1
X_5699_ _7211_/Q _5103_/A _5703_/S vssd1 vssd1 vccd1 vccd1 _5700_/A sky130_fd_sc_hd__mux2_1
X_7438_ _7438_/CLK _7438_/D vssd1 vssd1 vccd1 vccd1 _7438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7369_ _7838_/CLK _7369_/D vssd1 vssd1 vccd1 vccd1 _7369_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2448_ _5364_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2448_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_115_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2765_ clkbuf_0__2765_/X vssd1 vssd1 vccd1 vccd1 _5770__239/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3317_ clkbuf_0__3317_/X vssd1 vssd1 vccd1 vccd1 _7035__54/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6174__375 _6177__378/A vssd1 vssd1 vccd1 vccd1 _7427_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6740_ _6746_/A vssd1 vssd1 vccd1 vccd1 _6740_/X sky130_fd_sc_hd__buf_1
XFILLER_90_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3952_ _3952_/A vssd1 vssd1 vccd1 vccd1 _7651_/D sky130_fd_sc_hd__clkbuf_1
X_6671_ _6667_/Y _6670_/X _5970_/X vssd1 vssd1 vccd1 vccd1 _7671_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3883_ _3883_/A vssd1 vssd1 vccd1 vccd1 _7698_/D sky130_fd_sc_hd__clkbuf_1
X_5622_ _7695_/Q _7284_/Q _7167_/Q _7276_/Q _4296_/A _4302_/B vssd1 vssd1 vccd1 vccd1
+ _5622_/X sky130_fd_sc_hd__mux4_1
X_5553_ _5551_/X _5552_/X _5572_/S vssd1 vssd1 vccd1 vccd1 _5553_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4504_ _4504_/A vssd1 vssd1 vccd1 vccd1 _7441_/D sky130_fd_sc_hd__clkbuf_1
X_5484_ _7294_/Q _7286_/Q _7262_/Q _7110_/Q _5518_/A _4296_/A vssd1 vssd1 vccd1 vccd1
+ _5485_/B sky130_fd_sc_hd__mux4_2
X_7223_ _7339_/CLK _7223_/D vssd1 vssd1 vccd1 vccd1 _7223_/Q sky130_fd_sc_hd__dfxtp_1
X_4435_ _7461_/Q vssd1 vssd1 vccd1 vccd1 _5964_/A sky130_fd_sc_hd__buf_2
X_7154_ _7154_/CLK _7154_/D vssd1 vssd1 vccd1 vccd1 _7154_/Q sky130_fd_sc_hd__dfxtp_1
X_4366_ _4366_/A vssd1 vssd1 vccd1 vccd1 _7498_/D sky130_fd_sc_hd__clkbuf_1
X_6105_ _6111_/A vssd1 vssd1 vccd1 vccd1 _6105_/X sky130_fd_sc_hd__buf_1
XFILLER_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7085_ _5565_/X _7026_/A _7100_/C vssd1 vssd1 vccd1 vccd1 _7086_/B sky130_fd_sc_hd__mux2_1
XFILLER_58_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _4297_/A vssd1 vssd1 vccd1 vccd1 _4312_/A sky130_fd_sc_hd__buf_2
X_6036_ _7460_/Q vssd1 vssd1 vccd1 vccd1 _6036_/X sky130_fd_sc_hd__clkbuf_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2997_ _6167_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2997_/X sky130_fd_sc_hd__clkbuf_16
X_6938_ _7801_/Q _6952_/B vssd1 vssd1 vccd1 vccd1 _6938_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6869_ _6869_/A _6869_/B vssd1 vssd1 vccd1 vccd1 _6870_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6484__55 _6486__57/A vssd1 vssd1 vccd1 vccd1 _7600_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6651__121 _6651__121/A vssd1 vssd1 vccd1 vccd1 _7668_/CLK sky130_fd_sc_hd__inv_2
Xoutput107 _5132_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[22] sky130_fd_sc_hd__buf_2
Xoutput129 _5050_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[16] sky130_fd_sc_hd__buf_2
Xoutput118 _5099_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[7] sky130_fd_sc_hd__buf_2
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4220_ _4220_/A vssd1 vssd1 vccd1 vccd1 _7546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4151_ _4767_/A _4217_/B vssd1 vssd1 vccd1 vccd1 _4174_/S sky130_fd_sc_hd__nand2_4
XFILLER_95_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4082_ _4060_/X _7598_/Q _4082_/S vssd1 vssd1 vccd1 vccd1 _4083_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7841_ _7845_/CLK _7841_/D vssd1 vssd1 vccd1 vccd1 _7841_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6408__475 _6409__476/A vssd1 vssd1 vccd1 vccd1 _7540_/CLK sky130_fd_sc_hd__inv_2
X_7772_ _7772_/CLK _7772_/D vssd1 vssd1 vccd1 vccd1 _7772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4984_ _4984_/A vssd1 vssd1 vccd1 vccd1 _7111_/D sky130_fd_sc_hd__clkbuf_1
X_3935_ _3935_/A vssd1 vssd1 vccd1 vccd1 _3935_/X sky130_fd_sc_hd__clkbuf_4
X_6723_ _6723_/A _6723_/B _6723_/C vssd1 vssd1 vccd1 vccd1 _6724_/A sky130_fd_sc_hd__and3_1
Xclkbuf_0__2782_ _5852_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2782_/X sky130_fd_sc_hd__clkbuf_16
X_6654_ _6676_/A _6657_/A vssd1 vssd1 vccd1 vccd1 _6705_/D sky130_fd_sc_hd__and2b_1
XFILLER_109_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5605_ _7060_/A vssd1 vssd1 vccd1 vccd1 _5680_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3866_ _4285_/A _4285_/B vssd1 vssd1 vccd1 vccd1 _4286_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6585_ _6580_/X _6581_/Y _6582_/X _6584_/Y vssd1 vssd1 vccd1 vccd1 _6588_/C sky130_fd_sc_hd__o211a_1
X_3797_ _3794_/X _4303_/B _4304_/B _3796_/X vssd1 vssd1 vccd1 vccd1 _3800_/A sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_1_1_0__3297_ clkbuf_0__3297_/X vssd1 vssd1 vccd1 vccd1 _6753__140/A sky130_fd_sc_hd__clkbuf_4
X_5536_ _7240_/Q _7171_/Q _7481_/Q _7248_/Q _5479_/X _5518_/X vssd1 vssd1 vccd1 vccd1
+ _5536_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5467_ _5479_/A vssd1 vssd1 vccd1 vccd1 _5467_/X sky130_fd_sc_hd__buf_4
XFILLER_117_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7206_ _7477_/CLK _7206_/D vssd1 vssd1 vccd1 vccd1 _7206_/Q sky130_fd_sc_hd__dfxtp_1
X_4418_ _4417_/X _7478_/Q _4418_/S vssd1 vssd1 vccd1 vccd1 _4419_/A sky130_fd_sc_hd__mux2_1
X_5398_ _7225_/Q _7215_/Q _5458_/C _7214_/Q vssd1 vssd1 vccd1 vccd1 _5399_/D sky130_fd_sc_hd__or4b_1
XFILLER_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7137_ _7339_/CLK _7137_/D vssd1 vssd1 vccd1 vccd1 _7137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4349_ _4164_/X _7505_/Q _4349_/S vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7068_ _7048_/X _7068_/B vssd1 vssd1 vccd1 vccd1 _7069_/A sky130_fd_sc_hd__and2b_1
XFILLER_101_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6019_ _5932_/X _6004_/X _6018_/X _5993_/X vssd1 vssd1 vccd1 vccd1 _6019_/X sky130_fd_sc_hd__a211o_2
XFILLER_27_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3720_ _3720_/A vssd1 vssd1 vccd1 vccd1 _7746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3651_ _3927_/A _3927_/B vssd1 vssd1 vccd1 vccd1 _4578_/B sky130_fd_sc_hd__nor2_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3582_ _7465_/Q vssd1 vssd1 vccd1 vccd1 _4614_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5321_ _5321_/A vssd1 vssd1 vccd1 vccd1 _7149_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3082_ clkbuf_0__3082_/X vssd1 vssd1 vccd1 vccd1 _6266__382/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5183_ _7196_/Q _5189_/B _5185_/C vssd1 vssd1 vccd1 vccd1 _5183_/X sky130_fd_sc_hd__and3_1
X_4203_ _4161_/X _7551_/Q _4205_/S vssd1 vssd1 vccd1 vccd1 _4204_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4134_ _4134_/A vssd1 vssd1 vccd1 vccd1 _7578_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4065_ _4065_/A vssd1 vssd1 vccd1 vccd1 _7605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7824_ _7825_/CLK _7824_/D vssd1 vssd1 vccd1 vccd1 _7824_/Q sky130_fd_sc_hd__dfxtp_1
X_7755_ _7755_/CLK _7755_/D vssd1 vssd1 vccd1 vccd1 _7755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4967_ _4233_/X _7162_/Q _4971_/S vssd1 vssd1 vccd1 vccd1 _4968_/A sky130_fd_sc_hd__mux2_1
X_7686_ _7687_/CLK _7686_/D vssd1 vssd1 vccd1 vccd1 _7686_/Q sky130_fd_sc_hd__dfxtp_1
X_6706_ _6704_/Y _6705_/X _5970_/X vssd1 vssd1 vccd1 vccd1 _7681_/D sky130_fd_sc_hd__o21a_1
X_3918_ _3828_/X _7664_/Q _3918_/S vssd1 vssd1 vccd1 vccd1 _3919_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__2765_ _5765_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2765_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_32_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4898_ _4898_/A vssd1 vssd1 vccd1 vccd1 _7238_/D sky130_fd_sc_hd__clkbuf_1
X_6637_ _6637_/A _6637_/B vssd1 vssd1 vccd1 vccd1 _6640_/B sky130_fd_sc_hd__nand2_1
X_3849_ _3706_/X _7710_/Q _3853_/S vssd1 vssd1 vccd1 vccd1 _3850_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6568_ _6594_/A vssd1 vssd1 vccd1 vccd1 _6613_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5519_ _7239_/Q _7170_/Q _7480_/Q _7247_/Q _5479_/X _5518_/X vssd1 vssd1 vccd1 vccd1
+ _5519_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3317_ _6857_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3317_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_87_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__2447_ clkbuf_0__2447_/X vssd1 vssd1 vccd1 vccd1 _5362__193/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6850__44 _6850__44/A vssd1 vssd1 vccd1 vccd1 _7786_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5375__204 _5375__204/A vssd1 vssd1 vccd1 vccd1 _7176_/CLK sky130_fd_sc_hd__inv_2
X_5870_ _5044_/A hold3/A _5872_/S vssd1 vssd1 vccd1 vccd1 _5871_/A sky130_fd_sc_hd__mux2_1
X_4821_ _4820_/X _7271_/Q _4827_/S vssd1 vssd1 vccd1 vccd1 _4822_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4752_ _4752_/A vssd1 vssd1 vccd1 vccd1 _7300_/D sky130_fd_sc_hd__clkbuf_1
X_7540_ _7540_/CLK _7540_/D vssd1 vssd1 vccd1 vccd1 _7540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4683_ _4683_/A vssd1 vssd1 vccd1 vccd1 _7350_/D sky130_fd_sc_hd__clkbuf_1
X_3703_ _3932_/A vssd1 vssd1 vccd1 vccd1 _3703_/X sky130_fd_sc_hd__clkbuf_2
X_7471_ _7473_/CLK _7471_/D vssd1 vssd1 vccd1 vccd1 _7471_/Q sky130_fd_sc_hd__dfxtp_1
X_3634_ _3634_/A vssd1 vssd1 vccd1 vccd1 _7776_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3134_ clkbuf_0__3134_/X vssd1 vssd1 vccd1 vccd1 _6501_/A sky130_fd_sc_hd__clkbuf_4
X_3565_ _7825_/Q vssd1 vssd1 vccd1 vccd1 _3941_/A sky130_fd_sc_hd__buf_2
XFILLER_115_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5304_ _5303_/X _7339_/Q _5299_/X _5300_/X _7139_/Q vssd1 vssd1 vccd1 vccd1 _7139_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_103_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5235_ _7148_/Q _5199_/A _5204_/A _5234_/X vssd1 vssd1 vccd1 vccd1 _5235_/X sky130_fd_sc_hd__o22a_4
XFILLER_88_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5166_ _7122_/Q _5159_/X input30/X _5163_/X _5165_/X vssd1 vssd1 vccd1 vccd1 _5166_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5097_ _5097_/A vssd1 vssd1 vccd1 vccd1 _5097_/X sky130_fd_sc_hd__clkbuf_1
X_4117_ _3816_/X _7585_/Q _4123_/S vssd1 vssd1 vccd1 vccd1 _4118_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4048_ _4070_/S vssd1 vssd1 vccd1 vccd1 _4061_/S sky130_fd_sc_hd__buf_2
XFILLER_83_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5999_ _7723_/Q _7707_/Q _7426_/Q _7488_/Q _5933_/X _5998_/X vssd1 vssd1 vccd1 vccd1
+ _5999_/X sky130_fd_sc_hd__mux4_1
X_7807_ _7812_/CLK _7807_/D vssd1 vssd1 vccd1 vccd1 _7807_/Q sky130_fd_sc_hd__dfxtp_1
X_7738_ _7738_/CLK _7738_/D vssd1 vssd1 vccd1 vccd1 _7738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7669_ _7845_/CLK _7669_/D vssd1 vssd1 vccd1 vccd1 _7669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__2996_ clkbuf_0__2996_/X vssd1 vssd1 vccd1 vccd1 _6163__366/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6505__73 _6506__74/A vssd1 vssd1 vccd1 vccd1 _7618_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _7092_/A _5022_/B vssd1 vssd1 vccd1 vccd1 _5021_/A sky130_fd_sc_hd__or2_1
XFILLER_112_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6823__22 _6825__24/A vssd1 vssd1 vccd1 vccd1 _7764_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6971_ _6983_/B vssd1 vssd1 vccd1 vccd1 _6974_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4804_ _4955_/B _4847_/B vssd1 vssd1 vccd1 vccd1 _4827_/S sky130_fd_sc_hd__or2_2
X_7523_ _7523_/CLK _7523_/D vssd1 vssd1 vccd1 vccd1 _7523_/Q sky130_fd_sc_hd__dfxtp_1
X_4735_ _4710_/X _7307_/Q _4741_/S vssd1 vssd1 vccd1 vccd1 _4736_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7454_ _7454_/CLK _7454_/D vssd1 vssd1 vccd1 vccd1 _7454_/Q sky130_fd_sc_hd__dfxtp_1
X_4666_ _4417_/X _7357_/Q _4666_/S vssd1 vssd1 vccd1 vccd1 _4667_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4597_ _4612_/S vssd1 vssd1 vccd1 vccd1 _4606_/S sky130_fd_sc_hd__buf_2
X_7385_ _7385_/CLK _7385_/D vssd1 vssd1 vccd1 vccd1 _7385_/Q sky130_fd_sc_hd__dfxtp_1
X_3617_ _3617_/A vssd1 vssd1 vccd1 vccd1 _7783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3548_ _6325_/A _3630_/D _4434_/A vssd1 vssd1 vccd1 vccd1 _4028_/A sky130_fd_sc_hd__or3b_4
X_6336_ _6348_/A vssd1 vssd1 vccd1 vccd1 _6336_/X sky130_fd_sc_hd__buf_1
XFILLER_88_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__2781_ clkbuf_0__2781_/X vssd1 vssd1 vccd1 vccd1 _5851__304/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5218_ _5217_/X _5218_/B vssd1 vssd1 vccd1 vccd1 _5218_/X sky130_fd_sc_hd__and2b_1
X_6198_ _7803_/Q _6245_/A _6245_/B vssd1 vssd1 vccd1 vccd1 _6883_/A sky130_fd_sc_hd__nand3_2
XFILLER_57_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5149_ _5149_/A vssd1 vssd1 vccd1 vccd1 _5236_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6781__163 _6782__164/A vssd1 vssd1 vccd1 vccd1 _7730_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4520_ _4520_/A vssd1 vssd1 vccd1 vccd1 _7434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4451_ _4451_/A _4457_/A _4457_/B vssd1 vssd1 vccd1 vccd1 _4459_/A sky130_fd_sc_hd__and3_1
X_7170_ _7170_/CLK _7170_/D vssd1 vssd1 vccd1 vccd1 _7170_/Q sky130_fd_sc_hd__dfxtp_1
X_4382_ _4382_/A vssd1 vssd1 vccd1 vccd1 _7491_/D sky130_fd_sc_hd__clkbuf_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6052_ _6005_/X _6049_/X _6051_/X _5959_/X vssd1 vssd1 vccd1 vccd1 _6052_/X sky130_fd_sc_hd__o211a_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5003_/A vssd1 vssd1 vccd1 vccd1 _5003_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6954_ _6954_/A vssd1 vssd1 vccd1 vccd1 _6954_/X sky130_fd_sc_hd__clkbuf_2
X_5905_ _5905_/A vssd1 vssd1 vccd1 vccd1 _7346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6885_ _7846_/Q _6883_/Y _6884_/Y _5584_/X vssd1 vssd1 vccd1 vccd1 _6887_/B sky130_fd_sc_hd__a22o_1
XFILLER_34_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5698_ _5698_/A vssd1 vssd1 vccd1 vccd1 _7210_/D sky130_fd_sc_hd__clkbuf_1
X_4718_ _4718_/A vssd1 vssd1 vccd1 vccd1 _7313_/D sky130_fd_sc_hd__clkbuf_1
X_7506_ _7506_/CLK _7506_/D vssd1 vssd1 vccd1 vccd1 _7506_/Q sky130_fd_sc_hd__dfxtp_1
X_4649_ _4649_/A vssd1 vssd1 vccd1 vccd1 _7373_/D sky130_fd_sc_hd__clkbuf_1
X_7437_ _7437_/CLK _7437_/D vssd1 vssd1 vccd1 vccd1 _7437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7368_ _7838_/CLK _7368_/D vssd1 vssd1 vccd1 vccd1 _7368_/Q sky130_fd_sc_hd__dfxtp_1
X_5841__295 _5843__297/A vssd1 vssd1 vccd1 vccd1 _7312_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__2447_ _5358_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2447_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7299_ _7299_/CLK _7299_/D vssd1 vssd1 vccd1 vccd1 _7299_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__2764_ clkbuf_0__2764_/X vssd1 vssd1 vccd1 vccd1 _5771_/A sky130_fd_sc_hd__clkbuf_4
X_6319_ _7819_/Q _6319_/B vssd1 vssd1 vccd1 vccd1 _6320_/A sky130_fd_sc_hd__and2_1
XFILLER_89_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7348_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_76_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3316_ clkbuf_0__3316_/X vssd1 vssd1 vccd1 vccd1 _6856__49/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6788__169 _6788__169/A vssd1 vssd1 vccd1 vccd1 _7736_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6135__349 _6135__349/A vssd1 vssd1 vccd1 vccd1 _7398_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6443__504 _6443__504/A vssd1 vssd1 vccd1 vccd1 _7569_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3951_ _3950_/X _7651_/Q _3951_/S vssd1 vssd1 vccd1 vccd1 _3952_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6670_ _6711_/A _6670_/B _6670_/C _6711_/D vssd1 vssd1 vccd1 vccd1 _6670_/X sky130_fd_sc_hd__and4_1
X_3882_ _3836_/X _7698_/Q _3884_/S vssd1 vssd1 vccd1 vccd1 _3883_/A sky130_fd_sc_hd__mux2_1
X_5621_ _7300_/Q _7292_/Q _7268_/Q _7116_/Q _5413_/X _5416_/X vssd1 vssd1 vccd1 vccd1
+ _5621_/X sky130_fd_sc_hd__mux4_2
X_5552_ _7305_/Q _7233_/Q _7701_/Q _7321_/Q _5472_/A _5508_/X vssd1 vssd1 vccd1 vccd1
+ _5552_/X sky130_fd_sc_hd__mux4_1
X_4503_ _4417_/X _7441_/Q _4503_/S vssd1 vssd1 vccd1 vccd1 _4504_/A sky130_fd_sc_hd__mux2_1
X_6337__420 _6339__422/A vssd1 vssd1 vccd1 vccd1 _7483_/CLK sky130_fd_sc_hd__inv_2
X_5483_ _5480_/X _5482_/X _5572_/S vssd1 vssd1 vccd1 vccd1 _5483_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7222_ _7339_/CLK _7222_/D vssd1 vssd1 vccd1 vccd1 _7222_/Q sky130_fd_sc_hd__dfxtp_1
X_4434_ _4434_/A _4434_/B vssd1 vssd1 vccd1 vccd1 _7462_/D sky130_fd_sc_hd__nor2_1
X_7153_ _7339_/CLK _7153_/D vssd1 vssd1 vccd1 vccd1 _7153_/Q sky130_fd_sc_hd__dfxtp_1
X_4365_ _4161_/X _7498_/Q _4367_/S vssd1 vssd1 vccd1 vccd1 _4366_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__3108_ clkbuf_0__3108_/X vssd1 vssd1 vccd1 vccd1 _6373_/A sky130_fd_sc_hd__clkbuf_16
X_7084_ _7084_/A vssd1 vssd1 vccd1 vccd1 _7849_/D sky130_fd_sc_hd__clkbuf_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6035_ _4451_/A _6032_/X _6034_/X _5964_/X vssd1 vssd1 vccd1 vccd1 _6035_/X sky130_fd_sc_hd__o211a_1
XFILLER_100_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _4296_/A vssd1 vssd1 vccd1 vccd1 _4297_/A sky130_fd_sc_hd__clkbuf_4
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__2996_ _6161_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2996_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_81_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6937_ _6972_/B vssd1 vssd1 vccd1 vccd1 _6952_/B sky130_fd_sc_hd__clkbuf_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6868_ _6897_/A _6997_/A vssd1 vssd1 vccd1 vccd1 _6943_/A sky130_fd_sc_hd__or2_1
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__2816_ clkbuf_0__2816_/X vssd1 vssd1 vccd1 vccd1 _5929__323/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput108 _5134_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[23] sky130_fd_sc_hd__buf_2
Xoutput119 _5102_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[8] sky130_fd_sc_hd__buf_2
XFILLER_56_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4150_ _4286_/B _4150_/B _4865_/A vssd1 vssd1 vccd1 vccd1 _4767_/A sky130_fd_sc_hd__and3b_4
XFILLER_95_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4081_ _4081_/A vssd1 vssd1 vccd1 vccd1 _7599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7840_ _7840_/CLK _7840_/D vssd1 vssd1 vccd1 vccd1 _7840_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7771_ _7771_/CLK _7771_/D vssd1 vssd1 vccd1 vccd1 _7771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4983_ _7111_/Q _4411_/A _4987_/S vssd1 vssd1 vccd1 vccd1 _4984_/A sky130_fd_sc_hd__mux2_1
X_6722_ _6637_/A _6668_/B _6725_/D _6726_/B vssd1 vssd1 vccd1 vccd1 _6723_/C sky130_fd_sc_hd__o31ai_1
X_3934_ _3934_/A vssd1 vssd1 vccd1 vccd1 _7657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__2781_ _5846_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2781_/X sky130_fd_sc_hd__clkbuf_16
X_6653_ _6901_/A _6714_/A vssd1 vssd1 vccd1 vccd1 _6657_/A sky130_fd_sc_hd__nand2_1
X_3865_ _3865_/A vssd1 vssd1 vccd1 vccd1 _4285_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5604_ _5584_/X _5394_/Y _5448_/X _5603_/X vssd1 vssd1 vccd1 vccd1 _5604_/X sky130_fd_sc_hd__a22o_1
X_6584_ _7854_/Q _6584_/B vssd1 vssd1 vccd1 vccd1 _6584_/Y sky130_fd_sc_hd__xnor2_1
X_3796_ _7518_/Q _7523_/Q vssd1 vssd1 vccd1 vccd1 _3796_/X sky130_fd_sc_hd__and2b_1
X_5535_ _5533_/X _5534_/X _5575_/S vssd1 vssd1 vccd1 vccd1 _5535_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5466_ _5516_/A vssd1 vssd1 vccd1 vccd1 _5466_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7205_ _7839_/CLK _7205_/D vssd1 vssd1 vccd1 vccd1 _7205_/Q sky130_fd_sc_hd__dfxtp_1
X_4417_ _4417_/A vssd1 vssd1 vccd1 vccd1 _4417_/X sky130_fd_sc_hd__clkbuf_2
X_5397_ _7204_/Q vssd1 vssd1 vccd1 vccd1 _5462_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7136_ _7336_/CLK _7136_/D vssd1 vssd1 vccd1 vccd1 _7136_/Q sky130_fd_sc_hd__dfxtp_1
X_7871__198 vssd1 vssd1 vccd1 vccd1 _7871__198/HI core0Index[5] sky130_fd_sc_hd__conb_1
X_4348_ _4348_/A vssd1 vssd1 vccd1 vccd1 _7506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7067_ _5036_/A _6249_/A _7067_/S vssd1 vssd1 vccd1 vccd1 _7068_/B sky130_fd_sc_hd__mux2_1
XFILLER_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4279_ _4279_/A vssd1 vssd1 vccd1 vccd1 _7526_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6018_ _6010_/X _6017_/X _4452_/A vssd1 vssd1 vccd1 vccd1 _6018_/X sky130_fd_sc_hd__o21a_1
XFILLER_27_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2394_ clkbuf_0__2394_/X vssd1 vssd1 vccd1 vccd1 _5259__187/A sky130_fd_sc_hd__clkbuf_4
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5359__190 _5363__194/A vssd1 vssd1 vccd1 vccd1 _7162_/CLK sky130_fd_sc_hd__inv_2
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_33_wb_clk_i _7474_/CLK vssd1 vssd1 vccd1 vccd1 _7812_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_111_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3650_ _3650_/A vssd1 vssd1 vccd1 vccd1 _3927_/B sky130_fd_sc_hd__inv_2
X_3581_ _4009_/A vssd1 vssd1 vccd1 vccd1 _4614_/A sky130_fd_sc_hd__clkbuf_1
X_6293__404 _6293__404/A vssd1 vssd1 vccd1 vccd1 _7457_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5320_ _7016_/A _7149_/Q _5328_/S vssd1 vssd1 vccd1 vccd1 _5321_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4202_ _4202_/A vssd1 vssd1 vccd1 vccd1 _7552_/D sky130_fd_sc_hd__clkbuf_1
X_5182_ _7128_/Q _5173_/X input5/X _5177_/X _5181_/X vssd1 vssd1 vccd1 vccd1 _5182_/X
+ sky130_fd_sc_hd__a221o_4
X_6414__480 _6418__484/A vssd1 vssd1 vccd1 vccd1 _7545_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4133_ _4046_/X _7578_/Q _4141_/S vssd1 vssd1 vccd1 vccd1 _4134_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4064_ _4063_/X _7605_/Q _4070_/S vssd1 vssd1 vccd1 vccd1 _4065_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7823_ _7825_/CLK _7823_/D vssd1 vssd1 vccd1 vccd1 _7823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7754_ _7754_/CLK _7754_/D vssd1 vssd1 vccd1 vccd1 _7754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6705_ _6705_/A _6705_/B _6705_/C _6705_/D vssd1 vssd1 vccd1 vccd1 _6705_/X sky130_fd_sc_hd__and4_1
X_4966_ _4966_/A vssd1 vssd1 vccd1 vccd1 _7163_/D sky130_fd_sc_hd__clkbuf_1
X_7685_ _7685_/CLK _7685_/D vssd1 vssd1 vccd1 vccd1 _7685_/Q sky130_fd_sc_hd__dfxtp_1
X_3917_ _3917_/A vssd1 vssd1 vccd1 vccd1 _7665_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__2764_ _5764_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2764_/X sky130_fd_sc_hd__clkbuf_16
X_4897_ _4823_/X _7238_/Q _4899_/S vssd1 vssd1 vccd1 vccd1 _4898_/A sky130_fd_sc_hd__mux2_1
X_6636_ _6725_/B vssd1 vssd1 vccd1 vccd1 _6637_/A sky130_fd_sc_hd__inv_2
X_3848_ _3848_/A vssd1 vssd1 vccd1 vccd1 _7711_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6456__514 _6456__514/A vssd1 vssd1 vccd1 vccd1 _7579_/CLK sky130_fd_sc_hd__inv_2
X_6567_ _6711_/B _6711_/C _5661_/X vssd1 vssd1 vccd1 vccd1 _6567_/Y sky130_fd_sc_hd__a21oi_1
X_3779_ _3718_/X _7722_/Q _3781_/S vssd1 vssd1 vccd1 vccd1 _3780_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5518_ _5518_/A vssd1 vssd1 vccd1 vccd1 _5518_/X sky130_fd_sc_hd__buf_4
Xclkbuf_0__3316_ _6851_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3316_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_105_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5449_ _7040_/A _5437_/A _5448_/X _5338_/A vssd1 vssd1 vccd1 vccd1 _5647_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7119_ _7687_/CLK _7119_/D vssd1 vssd1 vccd1 vccd1 _7119_/Q sky130_fd_sc_hd__dfxtp_1
X_6745__134 _6745__134/A vssd1 vssd1 vccd1 vccd1 _7701_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6517__82 _6519__84/A vssd1 vssd1 vccd1 vccd1 _7627_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6835__31 _6836__32/A vssd1 vssd1 vccd1 vccd1 _7773_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4820_ _7470_/Q vssd1 vssd1 vccd1 vccd1 _4820_/X sky130_fd_sc_hd__buf_2
XFILLER_33_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4751_ _4705_/X _7300_/Q _4759_/S vssd1 vssd1 vccd1 vccd1 _4752_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4682_ _3672_/X _7350_/Q _4684_/S vssd1 vssd1 vccd1 vccd1 _4683_/A sky130_fd_sc_hd__mux2_1
X_3702_ _3702_/A vssd1 vssd1 vccd1 vccd1 _7752_/D sky130_fd_sc_hd__clkbuf_1
X_7470_ _7818_/CLK _7470_/D vssd1 vssd1 vccd1 vccd1 _7470_/Q sky130_fd_sc_hd__dfxtp_1
X_3633_ _3505_/X _7776_/Q _3641_/S vssd1 vssd1 vccd1 vccd1 _3634_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3133_ clkbuf_0__3133_/X vssd1 vssd1 vccd1 vccd1 _6770_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3564_ _3564_/A vssd1 vssd1 vccd1 vccd1 _7834_/D sky130_fd_sc_hd__clkbuf_1
X_5303_ _5303_/A vssd1 vssd1 vccd1 vccd1 _5303_/X sky130_fd_sc_hd__clkbuf_2
X_5234_ _5200_/X _5234_/B vssd1 vssd1 vccd1 vccd1 _5234_/X sky130_fd_sc_hd__and2b_1
XFILLER_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5165_ _7189_/Q _5175_/B _5171_/C vssd1 vssd1 vccd1 vccd1 _5165_/X sky130_fd_sc_hd__and3_1
XFILLER_68_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4116_ _4116_/A vssd1 vssd1 vccd1 vccd1 _7586_/D sky130_fd_sc_hd__clkbuf_1
X_5096_ _5096_/A _5098_/B vssd1 vssd1 vccd1 vccd1 _5097_/A sky130_fd_sc_hd__and2_1
XFILLER_83_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4047_ _4614_/D _4072_/B vssd1 vssd1 vccd1 vccd1 _4070_/S sky130_fd_sc_hd__or2_2
XFILLER_17_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6804__6 _6807__9/A vssd1 vssd1 vccd1 vccd1 _7748_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7806_ _7808_/CLK _7806_/D vssd1 vssd1 vccd1 vccd1 _7806_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _5998_/A vssd1 vssd1 vccd1 vccd1 _5998_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__2779_ clkbuf_0__2779_/X vssd1 vssd1 vccd1 vccd1 _5838__293/A sky130_fd_sc_hd__clkbuf_4
X_7737_ _7737_/CLK _7737_/D vssd1 vssd1 vccd1 vccd1 _7737_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2816_ _5925_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2816_/X sky130_fd_sc_hd__clkbuf_16
X_4949_ _4233_/X _7170_/Q _4953_/S vssd1 vssd1 vccd1 vccd1 _4950_/A sky130_fd_sc_hd__mux2_1
X_7668_ _7668_/CLK _7668_/D vssd1 vssd1 vccd1 vccd1 _7668_/Q sky130_fd_sc_hd__dfxtp_1
X_6619_ _7843_/Q _6705_/B _6705_/C vssd1 vssd1 vccd1 vccd1 _6619_/X sky130_fd_sc_hd__and3_1
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7599_ _7599_/CLK _7599_/D vssd1 vssd1 vccd1 vccd1 _7599_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__2995_ clkbuf_0__2995_/X vssd1 vssd1 vccd1 vccd1 _6160__364/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6331__415 _6333__417/A vssd1 vssd1 vccd1 vccd1 _7478_/CLK sky130_fd_sc_hd__inv_2
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6970_ _6859_/A _6997_/A _6900_/B vssd1 vssd1 vccd1 vccd1 _6983_/B sky130_fd_sc_hd__o21bai_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7863__237 vssd1 vssd1 vccd1 vccd1 partID[11] _7863__237/LO sky130_fd_sc_hd__conb_1
XFILLER_80_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5852_ _5852_/A vssd1 vssd1 vccd1 vccd1 _5852_/X sky130_fd_sc_hd__buf_1
XFILLER_22_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6264__380 _6266__382/A vssd1 vssd1 vccd1 vccd1 _7433_/CLK sky130_fd_sc_hd__inv_2
X_4803_ _7475_/Q vssd1 vssd1 vccd1 vccd1 _4803_/X sky130_fd_sc_hd__buf_2
X_5783_ _5789_/A vssd1 vssd1 vccd1 vccd1 _5783_/X sky130_fd_sc_hd__buf_1
XFILLER_119_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4734_ _4734_/A vssd1 vssd1 vccd1 vccd1 _7308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7522_ _7522_/CLK _7522_/D vssd1 vssd1 vccd1 vccd1 _7522_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_107_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7453_ _7453_/CLK _7453_/D vssd1 vssd1 vccd1 vccd1 _7453_/Q sky130_fd_sc_hd__dfxtp_1
X_4665_ _4665_/A vssd1 vssd1 vccd1 vccd1 _7358_/D sky130_fd_sc_hd__clkbuf_1
X_7384_ _7384_/CLK _7384_/D vssd1 vssd1 vccd1 vccd1 _7384_/Q sky130_fd_sc_hd__dfxtp_1
X_3616_ _3554_/X _7783_/Q _3622_/S vssd1 vssd1 vccd1 vccd1 _3617_/A sky130_fd_sc_hd__mux2_1
X_4596_ _4596_/A _4632_/B vssd1 vssd1 vccd1 vccd1 _4612_/S sky130_fd_sc_hd__nand2_2
Xclkbuf_1_1_0__3116_ clkbuf_0__3116_/X vssd1 vssd1 vccd1 vccd1 _6393__465/A sky130_fd_sc_hd__clkbuf_4
X_3547_ _3585_/A _3650_/A vssd1 vssd1 vccd1 vccd1 _4434_/A sky130_fd_sc_hd__and2_1
XFILLER_1_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__2780_ clkbuf_0__2780_/X vssd1 vssd1 vccd1 vccd1 _5843__297/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__2394_ _5256_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2394_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5217_ _5217_/A vssd1 vssd1 vccd1 vccd1 _5217_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6197_ _6197_/A vssd1 vssd1 vccd1 vccd1 _6245_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5148_ _5200_/A vssd1 vssd1 vccd1 vccd1 _5161_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5079_ _5079_/A _5081_/B vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__or2_1
XFILLER_57_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6427__490 _6428__491/A vssd1 vssd1 vccd1 vccd1 _7555_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5747__220 _5749__222/A vssd1 vssd1 vccd1 vccd1 _7237_/CLK sky130_fd_sc_hd__inv_2
X_4450_ _4450_/A _7477_/Q _6328_/C vssd1 vssd1 vccd1 vccd1 _4457_/B sky130_fd_sc_hd__and3_1
X_4381_ _7491_/Q _3935_/A _4385_/S vssd1 vssd1 vccd1 vccd1 _4382_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _6051_/A _6051_/B vssd1 vssd1 vccd1 vccd1 _6051_/X sky130_fd_sc_hd__or2_1
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5856_/A _5002_/B vssd1 vssd1 vccd1 vccd1 _5003_/A sky130_fd_sc_hd__and2_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6953_ _6943_/X _6939_/X _6249_/B vssd1 vssd1 vccd1 vccd1 _6953_/X sky130_fd_sc_hd__a21o_1
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5904_ _7346_/Q _5077_/A _5908_/S vssd1 vssd1 vccd1 vccd1 _5905_/A sky130_fd_sc_hd__mux2_1
X_6884_ _6884_/A _6884_/B vssd1 vssd1 vccd1 vccd1 _6884_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5697_ _7210_/Q _5101_/A _5703_/S vssd1 vssd1 vccd1 vccd1 _5698_/A sky130_fd_sc_hd__mux2_1
X_4717_ _4716_/X _7313_/Q _4720_/S vssd1 vssd1 vccd1 vccd1 _4718_/A sky130_fd_sc_hd__mux2_1
X_7505_ _7505_/CLK _7505_/D vssd1 vssd1 vccd1 vccd1 _7505_/Q sky130_fd_sc_hd__dfxtp_1
X_4648_ _3675_/X _7373_/Q _4648_/S vssd1 vssd1 vccd1 vccd1 _4649_/A sky130_fd_sc_hd__mux2_1
X_7436_ _7436_/CLK _7436_/D vssd1 vssd1 vccd1 vccd1 _7436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4579_ _4594_/S vssd1 vssd1 vccd1 vccd1 _4588_/S sky130_fd_sc_hd__clkbuf_2
X_7367_ _7838_/CLK _7367_/D vssd1 vssd1 vccd1 vccd1 _7367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6318_ _6318_/A vssd1 vssd1 vccd1 vccd1 _7472_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__2763_ clkbuf_0__2763_/X vssd1 vssd1 vccd1 vccd1 _5762__233/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7298_ _7298_/CLK _7298_/D vssd1 vssd1 vccd1 vccd1 _7298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6249_ _6249_/A _6249_/B vssd1 vssd1 vccd1 vccd1 _6250_/C sky130_fd_sc_hd__xor2_1
XFILLER_39_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6496__65 _6500__69/A vssd1 vssd1 vccd1 vccd1 _7610_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3315_ clkbuf_0__3315_/X vssd1 vssd1 vccd1 vccd1 _6850__44/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3950_ _3950_/A vssd1 vssd1 vccd1 vccd1 _3950_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_16_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3881_ _3881_/A vssd1 vssd1 vccd1 vccd1 _7699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5620_ _5613_/A _5617_/X _5619_/X vssd1 vssd1 vccd1 vccd1 _5620_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5551_ _7665_/Q _7498_/Q _7453_/Q _7313_/Q _5481_/X _5506_/X vssd1 vssd1 vccd1 vccd1
+ _5551_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6732__125 _6733__126/A vssd1 vssd1 vccd1 vccd1 _7691_/CLK sky130_fd_sc_hd__inv_2
X_4502_ _4502_/A vssd1 vssd1 vccd1 vccd1 _7442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7221_ _7336_/CLK _7221_/D vssd1 vssd1 vccd1 vccd1 _7221_/Q sky130_fd_sc_hd__dfxtp_1
X_5482_ _7302_/Q _7230_/Q _7698_/Q _7318_/Q _5479_/A _5481_/X vssd1 vssd1 vccd1 vccd1
+ _5482_/X sky130_fd_sc_hd__mux4_1
X_4433_ _3724_/A _4424_/C _4421_/X vssd1 vssd1 vccd1 vccd1 _4434_/B sky130_fd_sc_hd__o21ai_1
XFILLER_6_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7152_ _7154_/CLK _7152_/D vssd1 vssd1 vccd1 vccd1 _7152_/Q sky130_fd_sc_hd__dfxtp_1
X_4364_ _4364_/A vssd1 vssd1 vccd1 vccd1 _7499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6103_ _7372_/Q _6631_/B _6102_/X _5996_/A vssd1 vssd1 vccd1 vccd1 _7372_/D sky130_fd_sc_hd__o211a_1
X_7083_ _7106_/A _7083_/B vssd1 vssd1 vccd1 vccd1 _7084_/A sky130_fd_sc_hd__or2_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4295_ _5479_/A vssd1 vssd1 vccd1 vccd1 _4296_/A sky130_fd_sc_hd__buf_4
X_6034_ _6079_/A _6034_/B vssd1 vssd1 vccd1 vccd1 _6034_/X sky130_fd_sc_hd__or2_1
XFILLER_98_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6936_ _6933_/Y _6934_/X _6935_/X vssd1 vssd1 vccd1 vccd1 _7800_/D sky130_fd_sc_hd__a21oi_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2995_ _6155_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2995_/X sky130_fd_sc_hd__clkbuf_16
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6867_ _6993_/A _6867_/B _6867_/C _6867_/D vssd1 vssd1 vccd1 vccd1 _6997_/A sky130_fd_sc_hd__and4_2
X_7876__203 vssd1 vssd1 vccd1 vccd1 _7876__203/HI core1Index[3] sky130_fd_sc_hd__conb_1
X_7419_ _7419_/CLK _7419_/D vssd1 vssd1 vccd1 vccd1 _7419_/Q sky130_fd_sc_hd__dfxtp_1
X_6277__390 _6277__390/A vssd1 vssd1 vccd1 vccd1 _7443_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__2815_ clkbuf_0__2815_/X vssd1 vssd1 vccd1 vccd1 _5924__319/A sky130_fd_sc_hd__clkbuf_4
XFILLER_104_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6794__174 _6794__174/A vssd1 vssd1 vccd1 vccd1 _7741_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6141__354 _6141__354/A vssd1 vssd1 vccd1 vccd1 _7403_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput109 _5136_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[24] sky130_fd_sc_hd__buf_2
XFILLER_95_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4080_ _4057_/X _7599_/Q _4082_/S vssd1 vssd1 vccd1 vccd1 _4081_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7770_ _7770_/CLK _7770_/D vssd1 vssd1 vccd1 vccd1 _7770_/Q sky130_fd_sc_hd__dfxtp_1
X_4982_ _4982_/A vssd1 vssd1 vccd1 vccd1 _7112_/D sky130_fd_sc_hd__clkbuf_1
X_6721_ _6718_/A _6726_/B _7686_/Q vssd1 vssd1 vccd1 vccd1 _6723_/B sky130_fd_sc_hd__a21o_1
X_3933_ _3932_/X _7657_/Q _3942_/S vssd1 vssd1 vccd1 vccd1 _3934_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_3_wb_clk_i _7826_/CLK vssd1 vssd1 vccd1 vccd1 _5246_/A sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__2780_ _5840_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2780_/X sky130_fd_sc_hd__clkbuf_16
X_6652_ _6630_/B _6652_/B _6652_/C vssd1 vssd1 vccd1 vccd1 _6676_/A sky130_fd_sc_hd__and3b_1
X_3864_ _3805_/A _3588_/A _5239_/A vssd1 vssd1 vccd1 vccd1 _4280_/A sky130_fd_sc_hd__a21o_1
XFILLER_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5603_ _5396_/A _7077_/A _5602_/X _6396_/B vssd1 vssd1 vccd1 vccd1 _5603_/X sky130_fd_sc_hd__a31o_1
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6583_ _7670_/Q _6583_/B vssd1 vssd1 vccd1 vccd1 _6584_/B sky130_fd_sc_hd__xor2_1
X_3795_ _7525_/Q _7520_/Q vssd1 vssd1 vccd1 vccd1 _4303_/B sky130_fd_sc_hd__xnor2_1
X_5534_ _7304_/Q _7232_/Q _7700_/Q _7320_/Q _5472_/A _5508_/X vssd1 vssd1 vccd1 vccd1
+ _5534_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_1_1_0__3295_ clkbuf_0__3295_/X vssd1 vssd1 vccd1 vccd1 _6743__132/A sky130_fd_sc_hd__clkbuf_4
X_5465_ _7580_/Q _7564_/Q _7548_/Q _7540_/Q _4300_/A _4297_/A vssd1 vssd1 vccd1 vccd1
+ _5465_/X sky130_fd_sc_hd__mux4_2
X_6157__361 _6158__362/A vssd1 vssd1 vccd1 vccd1 _7413_/CLK sky130_fd_sc_hd__inv_2
X_7204_ _7826_/CLK _7204_/D vssd1 vssd1 vccd1 vccd1 _7204_/Q sky130_fd_sc_hd__dfxtp_1
X_4416_ _4416_/A vssd1 vssd1 vccd1 vccd1 _7479_/D sky130_fd_sc_hd__clkbuf_1
X_7135_ _7336_/CLK _7135_/D vssd1 vssd1 vccd1 vccd1 _7135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5396_ _5396_/A _7077_/A vssd1 vssd1 vccd1 vccd1 _5492_/A sky130_fd_sc_hd__nand2_1
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4347_ _4161_/X _7506_/Q _4349_/S vssd1 vssd1 vccd1 vccd1 _4348_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7066_ _7066_/A vssd1 vssd1 vccd1 vccd1 _7844_/D sky130_fd_sc_hd__clkbuf_1
X_4278_ _6394_/C _4278_/B _4278_/C vssd1 vssd1 vccd1 vccd1 _4279_/A sky130_fd_sc_hd__and3_1
X_6017_ _4451_/A _6012_/X _6016_/X _5964_/X vssd1 vssd1 vccd1 vccd1 _6017_/X sky130_fd_sc_hd__o211a_1
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__2393_ clkbuf_0__2393_/X vssd1 vssd1 vccd1 vccd1 _5376_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6919_ _6919_/A vssd1 vssd1 vccd1 vccd1 _6919_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3580_ _3580_/A vssd1 vssd1 vccd1 vccd1 _7830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4201_ _4158_/X _7552_/Q _4205_/S vssd1 vssd1 vccd1 vccd1 _4202_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5181_ _7195_/Q _5189_/B _5185_/C vssd1 vssd1 vccd1 vccd1 _5181_/X sky130_fd_sc_hd__and3_1
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4132_ _4147_/S vssd1 vssd1 vccd1 vccd1 _4141_/S sky130_fd_sc_hd__clkbuf_2
X_4063_ _7824_/Q vssd1 vssd1 vccd1 vccd1 _4063_/X sky130_fd_sc_hd__buf_2
XFILLER_83_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7822_ _7825_/CLK _7822_/D vssd1 vssd1 vccd1 vccd1 _7822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7753_ _7753_/CLK _7753_/D vssd1 vssd1 vccd1 vccd1 _7753_/Q sky130_fd_sc_hd__dfxtp_1
X_6380__455 _6381__456/A vssd1 vssd1 vccd1 vccd1 _7518_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4965_ _4230_/X _7163_/Q _4965_/S vssd1 vssd1 vccd1 vccd1 _4966_/A sky130_fd_sc_hd__mux2_1
X_6704_ _6656_/X _6658_/X _7681_/Q vssd1 vssd1 vccd1 vccd1 _6704_/Y sky130_fd_sc_hd__a21boi_1
X_3916_ _3824_/X _7665_/Q _3918_/S vssd1 vssd1 vccd1 vccd1 _3917_/A sky130_fd_sc_hd__mux2_1
X_7684_ _7684_/CLK _7684_/D vssd1 vssd1 vccd1 vccd1 _7684_/Q sky130_fd_sc_hd__dfxtp_1
X_6421__485 _6422__486/A vssd1 vssd1 vccd1 vccd1 _7550_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__2763_ _5758_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2763_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_20_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4896_ _4896_/A vssd1 vssd1 vccd1 vccd1 _7239_/D sky130_fd_sc_hd__clkbuf_1
X_6635_ _6635_/A vssd1 vssd1 vccd1 vccd1 _7659_/D sky130_fd_sc_hd__clkbuf_1
X_3847_ _3703_/X _7711_/Q _3853_/S vssd1 vssd1 vccd1 vccd1 _3848_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6566_ _7841_/Q _6711_/B _6711_/C vssd1 vssd1 vccd1 vccd1 _6566_/X sky130_fd_sc_hd__and3_1
X_3778_ _3778_/A vssd1 vssd1 vccd1 vccd1 _7723_/D sky130_fd_sc_hd__clkbuf_1
X_5517_ _5514_/X _5515_/X _5578_/S vssd1 vssd1 vccd1 vccd1 _5517_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3315_ _6845_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3315_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_3_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5448_ _5493_/C _5677_/B _5440_/X _5394_/C vssd1 vssd1 vccd1 vccd1 _5448_/X sky130_fd_sc_hd__o211a_1
XFILLER_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7118_ _7154_/CLK _7118_/D vssd1 vssd1 vccd1 vccd1 _7118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7049_ _7406_/Q _7077_/B vssd1 vssd1 vccd1 vccd1 _7074_/S sky130_fd_sc_hd__nand2_2
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5741__215 _5743__217/A vssd1 vssd1 vccd1 vccd1 _7232_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _4765_/S vssd1 vssd1 vccd1 vccd1 _4759_/S sky130_fd_sc_hd__buf_2
X_4681_ _4681_/A vssd1 vssd1 vccd1 vccd1 _7351_/D sky130_fd_sc_hd__clkbuf_1
X_3701_ _3698_/X _7752_/Q _3713_/S vssd1 vssd1 vccd1 vccd1 _3702_/A sky130_fd_sc_hd__mux2_1
X_3632_ _3647_/S vssd1 vssd1 vccd1 vccd1 _3641_/S sky130_fd_sc_hd__buf_2
X_6420_ _6444_/A vssd1 vssd1 vccd1 vccd1 _6420_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3132_ clkbuf_0__3132_/X vssd1 vssd1 vccd1 vccd1 _6478__532/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5302_ _5295_/X _7338_/Q _5299_/X _5300_/X _7138_/Q vssd1 vssd1 vccd1 vccd1 _7138_/D
+ sky130_fd_sc_hd__o32a_1
X_3563_ _3562_/X _7834_/Q _3567_/S vssd1 vssd1 vccd1 vccd1 _3564_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6282_ _6282_/A vssd1 vssd1 vccd1 vccd1 _6282_/X sky130_fd_sc_hd__buf_1
X_5233_ _7147_/Q _5199_/A _5204_/A _5232_/X vssd1 vssd1 vccd1 vccd1 _5233_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5164_ _5200_/A vssd1 vssd1 vccd1 vccd1 _5175_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4115_ _3784_/X _7586_/Q _4123_/S vssd1 vssd1 vccd1 vccd1 _4116_/A sky130_fd_sc_hd__mux2_1
X_5095_ _5095_/A vssd1 vssd1 vccd1 vccd1 _5095_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4046_ _7829_/Q vssd1 vssd1 vccd1 vccd1 _4046_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7805_ _7808_/CLK _7805_/D vssd1 vssd1 vccd1 vccd1 _7805_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _7366_/Q _5931_/X _5994_/X _5996_/X vssd1 vssd1 vccd1 vccd1 _7366_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_1_1_0__2778_ clkbuf_0__2778_/X vssd1 vssd1 vccd1 vccd1 _5830__286/A sky130_fd_sc_hd__clkbuf_4
X_7736_ _7736_/CLK _7736_/D vssd1 vssd1 vccd1 vccd1 _7736_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2815_ _5919_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2815_/X sky130_fd_sc_hd__clkbuf_16
X_4948_ _4948_/A vssd1 vssd1 vccd1 vccd1 _7171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7667_ _7667_/CLK _7667_/D vssd1 vssd1 vccd1 vccd1 _7667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4879_ _7246_/Q _4414_/A _4881_/S vssd1 vssd1 vccd1 vccd1 _4880_/A sky130_fd_sc_hd__mux2_1
X_6618_ _6594_/A _6569_/A _6617_/D _7681_/Q vssd1 vssd1 vccd1 vccd1 _6705_/C sky130_fd_sc_hd__a31o_1
XFILLER_116_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7598_ _7598_/CLK _7598_/D vssd1 vssd1 vccd1 vccd1 _7598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2994_ clkbuf_0__2994_/X vssd1 vssd1 vccd1 vccd1 _6263_/A sky130_fd_sc_hd__clkbuf_4
X_5805__267 _5805__267/A vssd1 vssd1 vccd1 vccd1 _7284_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4802_ _4802_/A vssd1 vssd1 vccd1 vccd1 _7277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4733_ _4705_/X _7308_/Q _4741_/S vssd1 vssd1 vccd1 vccd1 _4734_/A sky130_fd_sc_hd__mux2_1
X_7521_ _7521_/CLK _7521_/D vssd1 vssd1 vccd1 vccd1 _7521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7452_ _7452_/CLK _7452_/D vssd1 vssd1 vccd1 vccd1 _7452_/Q sky130_fd_sc_hd__dfxtp_1
X_4664_ _4414_/X _7358_/Q _4666_/S vssd1 vssd1 vccd1 vccd1 _4665_/A sky130_fd_sc_hd__mux2_1
X_4595_ _4595_/A vssd1 vssd1 vccd1 vccd1 _7397_/D sky130_fd_sc_hd__clkbuf_1
X_3615_ _3615_/A vssd1 vssd1 vccd1 vccd1 _7784_/D sky130_fd_sc_hd__clkbuf_1
X_7383_ _7383_/CLK _7383_/D vssd1 vssd1 vccd1 vccd1 _7383_/Q sky130_fd_sc_hd__dfxtp_1
X_3546_ _5676_/B _7476_/Q vssd1 vssd1 vccd1 vccd1 _3650_/A sky130_fd_sc_hd__and2b_1
Xclkbuf_1_1_0__3115_ clkbuf_0__3115_/X vssd1 vssd1 vccd1 vccd1 _6391__464/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__2393_ _5255_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2393_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5216_ _5216_/A vssd1 vssd1 vccd1 vccd1 _5216_/X sky130_fd_sc_hd__buf_2
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6511__78 _6512__79/A vssd1 vssd1 vccd1 vccd1 _7623_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6196_ _6228_/B vssd1 vssd1 vccd1 vccd1 _6245_/A sky130_fd_sc_hd__clkbuf_2
X_6271__385 _6273__387/A vssd1 vssd1 vccd1 vccd1 _7438_/CLK sky130_fd_sc_hd__inv_2
X_5147_ _7108_/Q vssd1 vssd1 vccd1 vccd1 _5200_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5078_ _5078_/A vssd1 vssd1 vccd1 vccd1 _5078_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4029_ _4044_/S vssd1 vssd1 vccd1 vccd1 _4038_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7719_ _7719_/CLK _7719_/D vssd1 vssd1 vccd1 vccd1 _7719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6393__465 _6393__465/A vssd1 vssd1 vccd1 vccd1 _7528_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5853__305 _5855__307/A vssd1 vssd1 vccd1 vccd1 _7322_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5259__187 _5259__187/A vssd1 vssd1 vccd1 vccd1 _7116_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4380_ _4380_/A vssd1 vssd1 vccd1 vccd1 _7492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6050_ _7591_/Q _7559_/Q _7834_/Q _7535_/Q _6013_/X _6014_/X vssd1 vssd1 vccd1 vccd1
+ _6051_/B sky130_fd_sc_hd__mux4_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5001_/A vssd1 vssd1 vccd1 vccd1 _5001_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6952_ _7805_/Q _6952_/B vssd1 vssd1 vccd1 vccd1 _6952_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5903_ _5903_/A vssd1 vssd1 vccd1 vccd1 _7345_/D sky130_fd_sc_hd__clkbuf_1
X_6883_ _6883_/A _6883_/B vssd1 vssd1 vccd1 vccd1 _6883_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5834_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5834_/X sky130_fd_sc_hd__buf_1
XFILLER_34_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5765_ _5771_/A vssd1 vssd1 vccd1 vccd1 _5765_/X sky130_fd_sc_hd__buf_1
X_5696_ _5696_/A vssd1 vssd1 vccd1 vccd1 _7209_/D sky130_fd_sc_hd__clkbuf_1
X_4716_ _7472_/Q vssd1 vssd1 vccd1 vccd1 _4716_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7504_ _7504_/CLK _7504_/D vssd1 vssd1 vccd1 vccd1 _7504_/Q sky130_fd_sc_hd__dfxtp_1
X_4647_ _4647_/A vssd1 vssd1 vccd1 vccd1 _7374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7435_ _7435_/CLK _7435_/D vssd1 vssd1 vccd1 vccd1 _7435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7366_ _7845_/CLK _7366_/D vssd1 vssd1 vccd1 vccd1 _7366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4578_ _4578_/A _4578_/B _4668_/B vssd1 vssd1 vccd1 vccd1 _4594_/S sky130_fd_sc_hd__and3_2
X_6317_ _7818_/Q _6319_/B vssd1 vssd1 vccd1 vccd1 _6318_/A sky130_fd_sc_hd__and2_1
XFILLER_116_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3529_ _7462_/Q vssd1 vssd1 vccd1 vccd1 _3585_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7297_ _7297_/CLK _7297_/D vssd1 vssd1 vccd1 vccd1 _7297_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__2762_ clkbuf_0__2762_/X vssd1 vssd1 vccd1 vccd1 _5755__227/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6248_ _7805_/Q _6248_/B vssd1 vssd1 vccd1 vccd1 _6249_/B sky130_fd_sc_hd__xor2_4
X_5917__313 _5918__314/A vssd1 vssd1 vccd1 vccd1 _7354_/CLK sky130_fd_sc_hd__inv_2
X_6179_ _7016_/A _3588_/X _7070_/A vssd1 vssd1 vccd1 vccd1 _7003_/A sky130_fd_sc_hd__a21oi_4
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3314_ clkbuf_0__3314_/X vssd1 vssd1 vccd1 vccd1 _6842__37/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7226_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3880_ _3832_/X _7699_/Q _3884_/S vssd1 vssd1 vccd1 vccd1 _3881_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5550_ _5548_/X _5549_/X _5569_/S vssd1 vssd1 vccd1 vccd1 _5550_/X sky130_fd_sc_hd__mux2_1
X_5481_ _5520_/A vssd1 vssd1 vccd1 vccd1 _5481_/X sky130_fd_sc_hd__buf_6
X_4501_ _4414_/X _7442_/Q _4503_/S vssd1 vssd1 vccd1 vccd1 _4502_/A sky130_fd_sc_hd__mux2_1
X_7220_ _7336_/CLK _7220_/D vssd1 vssd1 vccd1 vccd1 _7220_/Q sky130_fd_sc_hd__dfxtp_1
X_4432_ _3630_/D _4434_/A _4431_/Y vssd1 vssd1 vccd1 vccd1 _7463_/D sky130_fd_sc_hd__o21a_1
XFILLER_6_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7151_ _7344_/CLK _7151_/D vssd1 vssd1 vccd1 vccd1 _7151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4363_ _4158_/X _7499_/Q _4367_/S vssd1 vssd1 vccd1 vccd1 _4364_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6102_ _5932_/A _6092_/X _6101_/X _5993_/A vssd1 vssd1 vccd1 vccd1 _6102_/X sky130_fd_sc_hd__a211o_2
X_7082_ _5584_/X _7028_/A _7105_/C vssd1 vssd1 vccd1 vccd1 _7083_/B sky130_fd_sc_hd__mux2_1
XFILLER_59_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ _7519_/Q vssd1 vssd1 vccd1 vccd1 _5479_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6033_ _7392_/Q _7376_/Q _7646_/Q _7638_/Q _6013_/X _6014_/X vssd1 vssd1 vccd1 vccd1
+ _6034_/B sky130_fd_sc_hd__mux4_1
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6344__426 _6347__429/A vssd1 vssd1 vccd1 vccd1 _7489_/CLK sky130_fd_sc_hd__inv_2
X_6935_ _6954_/A vssd1 vssd1 vccd1 vccd1 _6935_/X sky130_fd_sc_hd__clkbuf_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2994_ _6154_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2994_/X sky130_fd_sc_hd__clkbuf_16
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6866_ _6866_/A _6866_/B vssd1 vssd1 vccd1 vccd1 _6867_/D sky130_fd_sc_hd__and2_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5679_ _5679_/A _5679_/B vssd1 vssd1 vccd1 vccd1 _5679_/Y sky130_fd_sc_hd__nand2_1
X_7418_ _7418_/CLK _7418_/D vssd1 vssd1 vccd1 vccd1 _7418_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__2814_ clkbuf_0__2814_/X vssd1 vssd1 vccd1 vccd1 _5918__314/A sky130_fd_sc_hd__clkbuf_4
X_7349_ _7349_/CLK _7349_/D vssd1 vssd1 vccd1 vccd1 _7349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput92 _7159_/Q vssd1 vssd1 vccd1 vccd1 caravel_uart_tx sky130_fd_sc_hd__buf_2
XFILLER_76_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5790__255 _5792__257/A vssd1 vssd1 vccd1 vccd1 _7272_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4981_ _7112_/Q _4408_/A _4987_/S vssd1 vssd1 vccd1 vccd1 _4982_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3932_ _3932_/A vssd1 vssd1 vccd1 vccd1 _3932_/X sky130_fd_sc_hd__clkbuf_4
X_6720_ _6720_/A vssd1 vssd1 vccd1 vccd1 _7685_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7899__226 vssd1 vssd1 vccd1 vccd1 _7899__226/HI versionID[0] sky130_fd_sc_hd__conb_1
X_3863_ _4111_/A vssd1 vssd1 vccd1 vccd1 _4731_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6582_ _7855_/Q _6583_/B vssd1 vssd1 vccd1 vccd1 _6582_/X sky130_fd_sc_hd__xor2_1
X_5602_ _5593_/X _5601_/X _5602_/S vssd1 vssd1 vccd1 vccd1 _5602_/X sky130_fd_sc_hd__mux2_2
XFILLER_118_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3794_ _7524_/Q _7523_/Q vssd1 vssd1 vccd1 vccd1 _3794_/X sky130_fd_sc_hd__and2_1
X_5533_ _7664_/Q _7497_/Q _7452_/Q _7312_/Q _5481_/X _5506_/X vssd1 vssd1 vccd1 vccd1
+ _5533_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3294_ clkbuf_0__3294_/X vssd1 vssd1 vccd1 vccd1 _6746_/A sky130_fd_sc_hd__clkbuf_4
X_5464_ _7522_/Q vssd1 vssd1 vccd1 vccd1 _5602_/S sky130_fd_sc_hd__buf_2
X_7203_ _7407_/CLK _7203_/D vssd1 vssd1 vccd1 vccd1 _7203_/Q sky130_fd_sc_hd__dfxtp_2
X_5395_ _5463_/A _5446_/A vssd1 vssd1 vccd1 vccd1 _7077_/A sky130_fd_sc_hd__nor2_1
X_4415_ _4414_/X _7479_/Q _4418_/S vssd1 vssd1 vccd1 vccd1 _4416_/A sky130_fd_sc_hd__mux2_1
X_7134_ _7336_/CLK _7134_/D vssd1 vssd1 vccd1 vccd1 _7134_/Q sky130_fd_sc_hd__dfxtp_1
X_4346_ _4346_/A vssd1 vssd1 vccd1 vccd1 _7507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7065_ _7048_/X _7065_/B vssd1 vssd1 vccd1 vccd1 _7066_/A sky130_fd_sc_hd__and2b_1
X_4277_ _7529_/Q _3791_/B _5461_/A _4901_/B vssd1 vssd1 vccd1 vccd1 _4278_/C sky130_fd_sc_hd__a31o_1
X_6016_ _6016_/A _6016_/B vssd1 vssd1 vccd1 vccd1 _6016_/X sky130_fd_sc_hd__or2_1
XFILLER_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__2392_ clkbuf_0__2392_/X vssd1 vssd1 vccd1 vccd1 _5254__184/A sky130_fd_sc_hd__clkbuf_4
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7033__52 _7035__54/A vssd1 vssd1 vccd1 vccd1 _7831_/CLK sky130_fd_sc_hd__inv_2
X_6918_ _6918_/A _6933_/B vssd1 vssd1 vccd1 vccd1 _6918_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6529__92 _6529__92/A vssd1 vssd1 vccd1 vccd1 _7637_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6847__41 _6848__42/A vssd1 vssd1 vccd1 vccd1 _7783_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5366__196 _5368__198/A vssd1 vssd1 vccd1 vccd1 _7168_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4200_ _4200_/A vssd1 vssd1 vccd1 vccd1 _7553_/D sky130_fd_sc_hd__clkbuf_1
X_5180_ _7127_/Q _5173_/X input4/X _5177_/X _5179_/X vssd1 vssd1 vccd1 vccd1 _5180_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4131_ _4131_/A _4614_/B _4614_/C _4131_/D vssd1 vssd1 vccd1 vccd1 _4147_/S sky130_fd_sc_hd__or4_4
XFILLER_3_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4062_ _4062_/A vssd1 vssd1 vccd1 vccd1 _7606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7821_ _7821_/CLK _7821_/D vssd1 vssd1 vccd1 vccd1 _7821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7752_ _7752_/CLK _7752_/D vssd1 vssd1 vccd1 vccd1 _7752_/Q sky130_fd_sc_hd__dfxtp_1
X_4964_ _4964_/A vssd1 vssd1 vccd1 vccd1 _7164_/D sky130_fd_sc_hd__clkbuf_1
X_6703_ _6701_/X _6702_/X _6690_/X vssd1 vssd1 vccd1 vccd1 _7680_/D sky130_fd_sc_hd__a21oi_1
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3915_ _3915_/A vssd1 vssd1 vccd1 vccd1 _7666_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__2762_ _5752_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2762_/X sky130_fd_sc_hd__clkbuf_16
X_7683_ _7684_/CLK _7683_/D vssd1 vssd1 vccd1 vccd1 _7683_/Q sky130_fd_sc_hd__dfxtp_1
X_4895_ _4820_/X _7239_/Q _4899_/S vssd1 vssd1 vccd1 vccd1 _4896_/A sky130_fd_sc_hd__mux2_1
X_6634_ _6723_/A _6634_/B _6637_/B vssd1 vssd1 vccd1 vccd1 _6635_/A sky130_fd_sc_hd__and3_1
X_3846_ _3846_/A vssd1 vssd1 vccd1 vccd1 _7712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6565_ _7682_/Q _6609_/B _7683_/Q vssd1 vssd1 vccd1 vccd1 _6711_/C sky130_fd_sc_hd__a21o_1
X_3777_ _3715_/X _7723_/Q _3781_/S vssd1 vssd1 vccd1 vccd1 _3778_/A sky130_fd_sc_hd__mux2_1
X_5516_ _5516_/A vssd1 vssd1 vccd1 vccd1 _5578_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_118_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3314_ _6839_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3314_/X sky130_fd_sc_hd__clkbuf_16
X_5447_ _5493_/A _5493_/B _5493_/D _5462_/A vssd1 vssd1 vccd1 vccd1 _5677_/B sky130_fd_sc_hd__or4b_1
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7117_ _7687_/CLK _7117_/D vssd1 vssd1 vccd1 vccd1 _7117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4329_ _4161_/X _7514_/Q _4331_/S vssd1 vssd1 vccd1 vccd1 _4330_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7048_ _7070_/A vssd1 vssd1 vccd1 vccd1 _7048_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6357__436 _6359__438/A vssd1 vssd1 vccd1 vccd1 _7499_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7036__1 _7039__4/A vssd1 vssd1 vccd1 vccd1 _7834_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _3722_/S vssd1 vssd1 vccd1 vccd1 _3713_/S sky130_fd_sc_hd__buf_2
XFILLER_14_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4680_ _3669_/X _7351_/Q _4684_/S vssd1 vssd1 vccd1 vccd1 _4681_/A sky130_fd_sc_hd__mux2_1
X_3631_ _3653_/B _4632_/A vssd1 vssd1 vccd1 vccd1 _3647_/S sky130_fd_sc_hd__nand2_2
X_3562_ _3938_/A vssd1 vssd1 vccd1 vccd1 _3562_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3131_ clkbuf_0__3131_/X vssd1 vssd1 vccd1 vccd1 _6474__529/A sky130_fd_sc_hd__clkbuf_4
X_5301_ _5295_/X _7337_/Q _5299_/X _5300_/X _7137_/Q vssd1 vssd1 vccd1 vccd1 _7137_/D
+ sky130_fd_sc_hd__o32a_1
X_6523__87 _6524__88/A vssd1 vssd1 vccd1 vccd1 _7632_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5232_ _5200_/X _5232_/B vssd1 vssd1 vccd1 vccd1 _5232_/X sky130_fd_sc_hd__and2b_1
X_5163_ _5177_/A vssd1 vssd1 vccd1 vccd1 _5163_/X sky130_fd_sc_hd__clkbuf_2
X_4114_ _4129_/S vssd1 vssd1 vccd1 vccd1 _4123_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_29_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5094_ _5094_/A _5098_/B vssd1 vssd1 vccd1 vccd1 _5095_/A sky130_fd_sc_hd__and2_1
XFILLER_84_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6841__36 _6842__37/A vssd1 vssd1 vccd1 vccd1 _7778_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4045_ _4045_/A vssd1 vssd1 vccd1 vccd1 _7611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7804_ _7808_/CLK _7804_/D vssd1 vssd1 vccd1 vccd1 _7804_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _5996_/A vssd1 vssd1 vccd1 vccd1 _5996_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2814_ _5913_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2814_/X sky130_fd_sc_hd__clkbuf_16
X_7735_ _7735_/CLK _7735_/D vssd1 vssd1 vccd1 vccd1 _7735_/Q sky130_fd_sc_hd__dfxtp_1
X_4947_ _4230_/X _7171_/Q _4947_/S vssd1 vssd1 vccd1 vccd1 _4948_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7666_ _7666_/CLK _7666_/D vssd1 vssd1 vccd1 vccd1 _7666_/Q sky130_fd_sc_hd__dfxtp_1
X_4878_ _4878_/A vssd1 vssd1 vccd1 vccd1 _7247_/D sky130_fd_sc_hd__clkbuf_1
X_6617_ _7681_/Q _6621_/B _6621_/C _6617_/D vssd1 vssd1 vccd1 vccd1 _6705_/B sky130_fd_sc_hd__nand4_1
X_3829_ _3828_/X _7716_/Q _3829_/S vssd1 vssd1 vccd1 vccd1 _3830_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5252__182 _5252__182/A vssd1 vssd1 vccd1 vccd1 _7111_/CLK sky130_fd_sc_hd__inv_2
X_7597_ _7597_/CLK _7597_/D vssd1 vssd1 vccd1 vccd1 _7597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_0 _7092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6439__500 _6443__504/A vssd1 vssd1 vccd1 vccd1 _7565_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4801_ _4728_/X _7277_/Q _4801_/S vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4732_ _4747_/S vssd1 vssd1 vccd1 vccd1 _4741_/S sky130_fd_sc_hd__buf_2
X_7520_ _7520_/CLK _7520_/D vssd1 vssd1 vccd1 vccd1 _7520_/Q sky130_fd_sc_hd__dfxtp_2
X_4663_ _4663_/A vssd1 vssd1 vccd1 vccd1 _7359_/D sky130_fd_sc_hd__clkbuf_1
X_7451_ _7451_/CLK _7451_/D vssd1 vssd1 vccd1 vccd1 _7451_/Q sky130_fd_sc_hd__dfxtp_1
X_3614_ _3505_/X _7784_/Q _3622_/S vssd1 vssd1 vccd1 vccd1 _3615_/A sky130_fd_sc_hd__mux2_1
X_4594_ _7397_/Q _3950_/A _4594_/S vssd1 vssd1 vccd1 vccd1 _4595_/A sky130_fd_sc_hd__mux2_1
X_7382_ _7382_/CLK _7382_/D vssd1 vssd1 vccd1 vccd1 _7382_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3114_ clkbuf_0__3114_/X vssd1 vssd1 vccd1 vccd1 _6392_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3545_ _3545_/A _3545_/B _3545_/C vssd1 vssd1 vccd1 vccd1 _5676_/B sky130_fd_sc_hd__and3_1
Xclkbuf_0__2392_ _5249_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2392_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5215_ _5215_/A vssd1 vssd1 vccd1 vccd1 _5215_/X sky130_fd_sc_hd__buf_2
XFILLER_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6195_ _6195_/A _6195_/B vssd1 vssd1 vccd1 vccd1 _6238_/A sky130_fd_sc_hd__xor2_1
X_5146_ _5177_/A vssd1 vssd1 vccd1 vccd1 _5146_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5077_ _5077_/A _5077_/B vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__or2_1
XFILLER_84_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4028_ _4028_/A _4072_/B vssd1 vssd1 vccd1 vccd1 _4044_/S sky130_fd_sc_hd__or2_2
XFILLER_84_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5979_ _6031_/A vssd1 vssd1 vccd1 vccd1 _5979_/X sky130_fd_sc_hd__buf_4
XFILLER_80_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5811__272 _5812__273/A vssd1 vssd1 vccd1 vccd1 _7289_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7718_ _7718_/CLK _7718_/D vssd1 vssd1 vccd1 vccd1 _7718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7649_ _7649_/CLK _7649_/D vssd1 vssd1 vccd1 vccd1 _7649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6434__496 _6435__497/A vssd1 vssd1 vccd1 vccd1 _7561_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5318_/A _5002_/B vssd1 vssd1 vccd1 vccd1 _5001_/A sky130_fd_sc_hd__and2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151__357 _6152__358/A vssd1 vssd1 vccd1 vccd1 _7409_/CLK sky130_fd_sc_hd__inv_2
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5754__226 _5755__227/A vssd1 vssd1 vccd1 vccd1 _7243_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6951_ _6949_/Y _6950_/X _6935_/X vssd1 vssd1 vccd1 vccd1 _7804_/D sky130_fd_sc_hd__a21oi_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5902_ _7345_/Q _5075_/A _5902_/S vssd1 vssd1 vccd1 vccd1 _5903_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6882_ _6882_/A _6882_/B _6882_/C _6222_/B vssd1 vssd1 vccd1 vccd1 _6887_/A sky130_fd_sc_hd__or4b_1
X_7867__194 vssd1 vssd1 vccd1 vccd1 _7867__194/HI core0Index[1] sky130_fd_sc_hd__conb_1
XFILLER_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5764_ _5795_/A vssd1 vssd1 vccd1 vccd1 _5764_/X sky130_fd_sc_hd__buf_1
X_7503_ _7503_/CLK _7503_/D vssd1 vssd1 vccd1 vccd1 _7503_/Q sky130_fd_sc_hd__dfxtp_1
X_5695_ _7209_/Q _5098_/A _5703_/S vssd1 vssd1 vccd1 vccd1 _5696_/A sky130_fd_sc_hd__mux2_1
X_4715_ _4715_/A vssd1 vssd1 vccd1 vccd1 _7314_/D sky130_fd_sc_hd__clkbuf_1
X_4646_ _3672_/X _7374_/Q _4648_/S vssd1 vssd1 vccd1 vccd1 _4647_/A sky130_fd_sc_hd__mux2_1
X_7434_ _7434_/CLK _7434_/D vssd1 vssd1 vccd1 vccd1 _7434_/Q sky130_fd_sc_hd__dfxtp_1
X_4577_ _4577_/A vssd1 vssd1 vccd1 vccd1 _7408_/D sky130_fd_sc_hd__clkbuf_1
X_7365_ _7679_/CLK _7365_/D vssd1 vssd1 vccd1 vccd1 _7365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6316_ _6316_/A vssd1 vssd1 vccd1 vccd1 _7471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3528_ _3678_/A vssd1 vssd1 vccd1 vccd1 _3630_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7296_ _7296_/CLK _7296_/D vssd1 vssd1 vccd1 vccd1 _7296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2761_ clkbuf_0__2761_/X vssd1 vssd1 vccd1 vccd1 _5751__224/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6247_ _6576_/A _6247_/B vssd1 vssd1 vccd1 vccd1 _6250_/B sky130_fd_sc_hd__xnor2_1
X_5129_ _7338_/Q _5131_/B vssd1 vssd1 vccd1 vccd1 _5130_/A sky130_fd_sc_hd__and2_1
XFILLER_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3313_ clkbuf_0__3313_/X vssd1 vssd1 vccd1 vccd1 _6838__34/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6289__400 _6292__403/A vssd1 vssd1 vccd1 vccd1 _7453_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5818__278 _5818__278/A vssd1 vssd1 vccd1 vccd1 _7295_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7901__228 vssd1 vssd1 vccd1 vccd1 _7901__228/HI versionID[2] sky130_fd_sc_hd__conb_1
XFILLER_117_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4500_ _4500_/A vssd1 vssd1 vccd1 vccd1 _7443_/D sky130_fd_sc_hd__clkbuf_1
X_5480_ _7662_/Q _7495_/Q _7450_/Q _7310_/Q _5518_/A _5479_/X vssd1 vssd1 vccd1 vccd1
+ _5480_/X sky130_fd_sc_hd__mux4_1
X_4431_ _6325_/A _4431_/B vssd1 vssd1 vccd1 vccd1 _4431_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7150_ _7154_/CLK _7150_/D vssd1 vssd1 vccd1 vccd1 _7150_/Q sky130_fd_sc_hd__dfxtp_1
X_4362_ _4362_/A vssd1 vssd1 vccd1 vccd1 _7500_/D sky130_fd_sc_hd__clkbuf_1
X_6101_ _6096_/X _6100_/X _6036_/X vssd1 vssd1 vccd1 vccd1 _6101_/X sky130_fd_sc_hd__o21a_1
X_7081_ _7081_/A vssd1 vssd1 vccd1 vccd1 _7848_/D sky130_fd_sc_hd__clkbuf_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _5611_/S vssd1 vssd1 vccd1 vccd1 _5613_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6032_ _7411_/Q _7352_/Q _7419_/Q _7400_/Q _6031_/X _6011_/X vssd1 vssd1 vccd1 vccd1
+ _6032_/X sky130_fd_sc_hd__mux4_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6934_ _6924_/X _6907_/X _6884_/Y vssd1 vssd1 vccd1 vccd1 _6934_/X sky130_fd_sc_hd__a21o_1
XFILLER_54_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6865_ _6213_/Y _6214_/X _6864_/X _6208_/B _6238_/A vssd1 vssd1 vccd1 vccd1 _6867_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7417_ _7417_/CLK _7417_/D vssd1 vssd1 vccd1 vccd1 _7417_/Q sky130_fd_sc_hd__dfxtp_1
X_5678_ _6901_/A _6326_/B _6325_/B vssd1 vssd1 vccd1 vccd1 _5735_/A sky130_fd_sc_hd__or3_1
X_4629_ _4629_/A vssd1 vssd1 vccd1 vccd1 _7382_/D sky130_fd_sc_hd__clkbuf_1
X_7348_ _7348_/CLK _7348_/D vssd1 vssd1 vccd1 vccd1 _7348_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__2813_ clkbuf_0__2813_/X vssd1 vssd1 vccd1 vccd1 _6111_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7279_ _7279_/CLK _7279_/D vssd1 vssd1 vccd1 vccd1 _7279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6284__396 _6287__399/A vssd1 vssd1 vccd1 vccd1 _7449_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3089_ clkbuf_0__3089_/X vssd1 vssd1 vccd1 vccd1 _6450_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput93 _5084_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[0] sky130_fd_sc_hd__buf_2
XFILLER_95_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4980_ _4980_/A vssd1 vssd1 vccd1 vccd1 _7113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3931_ _3931_/A vssd1 vssd1 vccd1 vccd1 _7658_/D sky130_fd_sc_hd__clkbuf_1
X_6304__411 _6306__413/A vssd1 vssd1 vccd1 vccd1 _7464_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3862_ _3907_/B vssd1 vssd1 vccd1 vccd1 _4901_/B sky130_fd_sc_hd__clkbuf_2
X_6581_ _6670_/B _6670_/C _7095_/B vssd1 vssd1 vccd1 vccd1 _6581_/Y sky130_fd_sc_hd__a21oi_1
X_5601_ _5595_/X _5597_/X _5600_/X _4291_/A vssd1 vssd1 vccd1 vccd1 _5601_/X sky130_fd_sc_hd__o22a_1
X_3793_ _3787_/X _4304_/B _4271_/A _4303_/C vssd1 vssd1 vccd1 vccd1 _3802_/A sky130_fd_sc_hd__a22o_1
X_5532_ _5530_/X _5531_/X _5569_/S vssd1 vssd1 vccd1 vccd1 _5532_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5463_ _5463_/A _5495_/A vssd1 vssd1 vccd1 vccd1 _5463_/Y sky130_fd_sc_hd__nor2_2
XFILLER_8_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7202_ _7407_/CLK _7202_/D vssd1 vssd1 vccd1 vccd1 _7202_/Q sky130_fd_sc_hd__dfxtp_1
X_5394_ _5463_/A _5682_/A _5394_/C vssd1 vssd1 vccd1 vccd1 _5394_/Y sky130_fd_sc_hd__nor3_1
X_4414_ _4414_/A vssd1 vssd1 vccd1 vccd1 _4414_/X sky130_fd_sc_hd__clkbuf_2
X_7133_ _7336_/CLK _7133_/D vssd1 vssd1 vccd1 vccd1 _7133_/Q sky130_fd_sc_hd__dfxtp_1
X_4345_ _4158_/X _7507_/Q _4349_/S vssd1 vssd1 vccd1 vccd1 _4346_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6350__431 _6353__434/A vssd1 vssd1 vccd1 vccd1 _7494_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7064_ _5038_/A _6242_/A _7067_/S vssd1 vssd1 vccd1 vccd1 _7065_/B sky130_fd_sc_hd__mux2_1
X_4276_ _6310_/A vssd1 vssd1 vccd1 vccd1 _6394_/C sky130_fd_sc_hd__buf_2
X_6015_ _7391_/Q _7375_/Q _7645_/Q _7637_/Q _6013_/X _6014_/X vssd1 vssd1 vccd1 vccd1
+ _6016_/B sky130_fd_sc_hd__mux4_2
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2391_ clkbuf_0__2391_/X vssd1 vssd1 vccd1 vccd1 _7039__4/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6917_ _6972_/B vssd1 vssd1 vccd1 vccd1 _6933_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6164__367 _6166__369/A vssd1 vssd1 vccd1 vccd1 _7419_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5767__236 _5769__238/A vssd1 vssd1 vccd1 vccd1 _7253_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7372_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_7859__233 vssd1 vssd1 vccd1 vccd1 partID[4] _7859__233/LO sky130_fd_sc_hd__conb_1
XFILLER_114_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4130_ _4130_/A vssd1 vssd1 vccd1 vccd1 _7579_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4061_ _4060_/X _7606_/Q _4061_/S vssd1 vssd1 vccd1 vccd1 _4062_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7820_ _7821_/CLK _7820_/D vssd1 vssd1 vccd1 vccd1 _7820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7751_ _7751_/CLK _7751_/D vssd1 vssd1 vccd1 vccd1 _7751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4963_ _4227_/X _7164_/Q _4965_/S vssd1 vssd1 vccd1 vccd1 _4964_/A sky130_fd_sc_hd__mux2_1
X_7682_ _7684_/CLK _7682_/D vssd1 vssd1 vccd1 vccd1 _7682_/Q sky130_fd_sc_hd__dfxtp_1
X_6702_ _6708_/A _6702_/B _6702_/C vssd1 vssd1 vccd1 vccd1 _6702_/X sky130_fd_sc_hd__or3_1
XFILLER_51_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3914_ _3820_/X _7666_/Q _3918_/S vssd1 vssd1 vccd1 vccd1 _3915_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__2761_ _5746_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2761_/X sky130_fd_sc_hd__clkbuf_16
X_6633_ _5993_/A _6630_/X _6725_/C vssd1 vssd1 vccd1 vccd1 _6637_/B sky130_fd_sc_hd__a21o_1
X_4894_ _4894_/A vssd1 vssd1 vccd1 vccd1 _7240_/D sky130_fd_sc_hd__clkbuf_1
X_3845_ _3698_/X _7712_/Q _3853_/S vssd1 vssd1 vccd1 vccd1 _3846_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6564_ _7683_/Q _7682_/Q _6609_/B vssd1 vssd1 vccd1 vccd1 _6711_/B sky130_fd_sc_hd__nand3_2
X_3776_ _3776_/A vssd1 vssd1 vccd1 vccd1 _7724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5515_ _7178_/Q _7359_/Q _7715_/Q _7255_/Q _5512_/X _5513_/X vssd1 vssd1 vccd1 vccd1
+ _5515_/X sky130_fd_sc_hd__mux4_1
X_6495_ _6501_/A vssd1 vssd1 vccd1 vccd1 _6495_/X sky130_fd_sc_hd__buf_1
XFILLER_106_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3313_ _6833_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3313_/X sky130_fd_sc_hd__clkbuf_16
X_5446_ _5446_/A _5446_/B vssd1 vssd1 vccd1 vccd1 _5493_/D sky130_fd_sc_hd__or2_1
XFILLER_99_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4328_ _4328_/A vssd1 vssd1 vccd1 vccd1 _7515_/D sky130_fd_sc_hd__clkbuf_1
X_7116_ _7116_/CLK _7116_/D vssd1 vssd1 vccd1 vccd1 _7116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7047_ _7047_/A vssd1 vssd1 vccd1 vccd1 _7839_/D sky130_fd_sc_hd__clkbuf_1
X_4259_ _7824_/Q vssd1 vssd1 vccd1 vccd1 _4259_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3630_ _3724_/A _4424_/C _3630_/C _3630_/D vssd1 vssd1 vccd1 vccd1 _4632_/A sky130_fd_sc_hd__and4b_4
X_3561_ _7826_/Q vssd1 vssd1 vccd1 vccd1 _3938_/A sky130_fd_sc_hd__clkbuf_4
X_5300_ _5308_/A vssd1 vssd1 vccd1 vccd1 _5300_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5231_ _7146_/Q _5199_/A _5204_/A _5230_/X vssd1 vssd1 vccd1 vccd1 _5231_/X sky130_fd_sc_hd__o22a_4
XFILLER_88_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5162_ _7121_/Q _5159_/X input29/X _5146_/X _5161_/X vssd1 vssd1 vccd1 vccd1 _5162_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_68_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5093_ _5093_/A vssd1 vssd1 vccd1 vccd1 _5093_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4113_ _4883_/A _4217_/B vssd1 vssd1 vccd1 vccd1 _4129_/S sky130_fd_sc_hd__nand2_2
XFILLER_96_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5837__292 _5838__293/A vssd1 vssd1 vccd1 vccd1 _7309_/CLK sky130_fd_sc_hd__inv_2
X_4044_ _3950_/X _7611_/Q _4044_/S vssd1 vssd1 vccd1 vccd1 _4045_/A sky130_fd_sc_hd__mux2_1
X_5911__309 _5911__309/A vssd1 vssd1 vccd1 vccd1 _7350_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7803_ _7808_/CLK _7803_/D vssd1 vssd1 vccd1 vccd1 _7803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__2813_ _5912_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2813_/X sky130_fd_sc_hd__clkbuf_16
X_5995_ _6737_/S vssd1 vssd1 vccd1 vccd1 _5996_/A sky130_fd_sc_hd__clkbuf_2
X_7734_ _7734_/CLK _7734_/D vssd1 vssd1 vccd1 vccd1 _7734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4946_ _4946_/A vssd1 vssd1 vccd1 vccd1 _7172_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7665_ _7665_/CLK _7665_/D vssd1 vssd1 vccd1 vccd1 _7665_/Q sky130_fd_sc_hd__dfxtp_1
X_4877_ _7247_/Q _4411_/A _4881_/S vssd1 vssd1 vccd1 vccd1 _4878_/A sky130_fd_sc_hd__mux2_1
X_6616_ _6189_/A _6708_/B _6702_/B _6242_/A vssd1 vssd1 vccd1 vccd1 _6616_/X sky130_fd_sc_hd__o2bb2a_1
X_3828_ _4408_/A vssd1 vssd1 vccd1 vccd1 _3828_/X sky130_fd_sc_hd__clkbuf_4
X_7596_ _7596_/CLK _7596_/D vssd1 vssd1 vccd1 vccd1 _7596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3759_ _3759_/A vssd1 vssd1 vccd1 vccd1 _7731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5429_ _5424_/X _5428_/X _5432_/S vssd1 vssd1 vccd1 vccd1 _5429_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_1 _3663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3089_ _6300_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3089_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6363__441 _6363__441/A vssd1 vssd1 vccd1 vccd1 _7504_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6648__119 _6648__119/A vssd1 vssd1 vccd1 vccd1 _7666_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4800_ _4800_/A vssd1 vssd1 vccd1 vccd1 _7278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4731_ _4901_/A _4901_/B _4731_/C _4919_/B vssd1 vssd1 vccd1 vccd1 _4747_/S sky130_fd_sc_hd__or4_4
X_4662_ _4411_/X _7359_/Q _4666_/S vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__mux2_1
X_7450_ _7450_/CLK _7450_/D vssd1 vssd1 vccd1 vccd1 _7450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3613_ _3628_/S vssd1 vssd1 vccd1 vccd1 _3622_/S sky130_fd_sc_hd__buf_2
X_6401_ _6413_/A vssd1 vssd1 vccd1 vccd1 _6401_/X sky130_fd_sc_hd__buf_1
X_4593_ _4593_/A vssd1 vssd1 vccd1 vccd1 _7398_/D sky130_fd_sc_hd__clkbuf_1
X_7381_ _7381_/CLK _7381_/D vssd1 vssd1 vccd1 vccd1 _7381_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3113_ clkbuf_0__3113_/X vssd1 vssd1 vccd1 vccd1 _6381__456/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3544_ _3927_/A _4447_/A _4424_/B _3542_/Y _3543_/X vssd1 vssd1 vccd1 vccd1 _3545_/C
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_0__2391_ _5248_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2391_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6263_ _6263_/A vssd1 vssd1 vccd1 vccd1 _6263_/X sky130_fd_sc_hd__buf_1
XFILLER_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5214_ _7139_/Q _5199_/X _5204_/X _5213_/X vssd1 vssd1 vccd1 vccd1 _5214_/X sky130_fd_sc_hd__o22a_4
XFILLER_88_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6194_ _6194_/A vssd1 vssd1 vccd1 vccd1 _6195_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5145_ _5187_/A vssd1 vssd1 vccd1 vccd1 _5145_/X sky130_fd_sc_hd__buf_2
XFILLER_96_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _5076_/A vssd1 vssd1 vccd1 vccd1 _5076_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4027_ _4027_/A vssd1 vssd1 vccd1 vccd1 _7619_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _6051_/A vssd1 vssd1 vccd1 vccd1 _5978_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7717_ _7717_/CLK _7717_/D vssd1 vssd1 vccd1 vccd1 _7717_/Q sky130_fd_sc_hd__dfxtp_1
X_4929_ _4230_/X _7179_/Q _4929_/S vssd1 vssd1 vccd1 vccd1 _4930_/A sky130_fd_sc_hd__mux2_1
X_7648_ _7648_/CLK _7648_/D vssd1 vssd1 vccd1 vccd1 _7648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7579_ _7579_/CLK _7579_/D vssd1 vssd1 vccd1 vccd1 _7579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6137__350 _6138__351/A vssd1 vssd1 vccd1 vccd1 _7399_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6950_ _6943_/X _6939_/X _6247_/B vssd1 vssd1 vccd1 vccd1 _6950_/X sky130_fd_sc_hd__a21o_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5901_ _5901_/A vssd1 vssd1 vccd1 vccd1 _7344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6881_ _7851_/Q _6881_/B vssd1 vssd1 vccd1 vccd1 _6882_/C sky130_fd_sc_hd__xnor2_1
XFILLER_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4714_ _4713_/X _7314_/Q _4720_/S vssd1 vssd1 vccd1 vccd1 _4715_/A sky130_fd_sc_hd__mux2_1
X_7502_ _7502_/CLK _7502_/D vssd1 vssd1 vccd1 vccd1 _7502_/Q sky130_fd_sc_hd__dfxtp_1
X_5694_ _5727_/A vssd1 vssd1 vccd1 vccd1 _5703_/S sky130_fd_sc_hd__buf_4
XFILLER_30_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4645_ _4645_/A vssd1 vssd1 vccd1 vccd1 _7375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7433_ _7433_/CLK _7433_/D vssd1 vssd1 vccd1 vccd1 _7433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4576_ _4265_/X _7408_/Q _4576_/S vssd1 vssd1 vccd1 vccd1 _4577_/A sky130_fd_sc_hd__mux2_1
X_7364_ _7364_/CLK _7364_/D vssd1 vssd1 vccd1 vccd1 _7364_/Q sky130_fd_sc_hd__dfxtp_1
X_3527_ _7463_/Q vssd1 vssd1 vccd1 vccd1 _3678_/A sky130_fd_sc_hd__clkbuf_2
X_6315_ _7817_/Q _6319_/B vssd1 vssd1 vccd1 vccd1 _6316_/A sky130_fd_sc_hd__and2_1
XFILLER_115_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2760_ clkbuf_0__2760_/X vssd1 vssd1 vccd1 vccd1 _5743__217/A sky130_fd_sc_hd__clkbuf_4
X_7295_ _7295_/CLK _7295_/D vssd1 vssd1 vccd1 vccd1 _7295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6246_ _6244_/Y _6883_/A _6248_/B vssd1 vssd1 vccd1 vccd1 _6247_/B sky130_fd_sc_hd__a21bo_1
X_5128_ _5128_/A vssd1 vssd1 vccd1 vccd1 _5128_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3312_ clkbuf_0__3312_/X vssd1 vssd1 vccd1 vccd1 _6857_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5059_ _5059_/A vssd1 vssd1 vccd1 vccd1 _5059_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5371__200 _5374__203/A vssd1 vssd1 vccd1 vccd1 _7172_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5924__319 _5924__319/A vssd1 vssd1 vccd1 vccd1 _7360_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_wb_clk_i _7474_/CLK vssd1 vssd1 vccd1 vccd1 _7818_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4430_ _3991_/C _4431_/B _4429_/Y vssd1 vssd1 vccd1 vccd1 _7464_/D sky130_fd_sc_hd__a21oi_1
X_5760__231 _5762__233/A vssd1 vssd1 vccd1 vccd1 _7248_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6100_ _6005_/X _6097_/X _6099_/X _5959_/A vssd1 vssd1 vccd1 vccd1 _6100_/X sky130_fd_sc_hd__o211a_1
X_4361_ _4155_/X _7500_/Q _4367_/S vssd1 vssd1 vccd1 vccd1 _4362_/A sky130_fd_sc_hd__mux2_1
X_7080_ _7070_/X _7080_/B vssd1 vssd1 vccd1 vccd1 _7081_/A sky130_fd_sc_hd__and2b_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4292_ _7520_/Q vssd1 vssd1 vccd1 vccd1 _5611_/S sky130_fd_sc_hd__buf_2
X_6031_ _6031_/A vssd1 vssd1 vccd1 vccd1 _6031_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6933_ _6933_/A _6933_/B vssd1 vssd1 vccd1 vccd1 _6933_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6864_ _6235_/Y _6236_/X _6225_/X _6991_/C _6229_/X vssd1 vssd1 vccd1 vccd1 _6864_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_62_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6795_ _6795_/A vssd1 vssd1 vccd1 vccd1 _6795_/X sky130_fd_sc_hd__buf_1
X_5746_ _5758_/A vssd1 vssd1 vccd1 vccd1 _5746_/X sky130_fd_sc_hd__buf_1
XFILLER_108_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5677_ _7040_/A _5677_/B vssd1 vssd1 vccd1 vccd1 _6325_/B sky130_fd_sc_hd__or2_2
X_7416_ _7416_/CLK _7416_/D vssd1 vssd1 vccd1 vccd1 _7416_/Q sky130_fd_sc_hd__dfxtp_1
X_4628_ _3672_/X _7382_/Q _4630_/S vssd1 vssd1 vccd1 vccd1 _4629_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__2389_ clkbuf_0__2389_/X vssd1 vssd1 vccd1 vccd1 _6832_/A sky130_fd_sc_hd__clkbuf_4
X_7347_ _7348_/CLK _7347_/D vssd1 vssd1 vccd1 vccd1 _7347_/Q sky130_fd_sc_hd__dfxtp_1
X_4559_ _4559_/A vssd1 vssd1 vccd1 vccd1 _7416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7278_ _7278_/CLK _7278_/D vssd1 vssd1 vccd1 vccd1 _7278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6229_ _7851_/Q _6890_/B vssd1 vssd1 vccd1 vccd1 _6229_/X sky130_fd_sc_hd__xor2_1
XFILLER_66_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3088_ clkbuf_0__3088_/X vssd1 vssd1 vccd1 vccd1 _6298__408/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5824__283 _5824__283/A vssd1 vssd1 vccd1 vccd1 _7300_/CLK sky130_fd_sc_hd__inv_2
Xoutput94 _5106_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[10] sky130_fd_sc_hd__buf_2
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5378__206 _5378__206/A vssd1 vssd1 vccd1 vccd1 _7178_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3930_ _3926_/X _7658_/Q _3942_/S vssd1 vssd1 vccd1 vccd1 _3931_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5831__287 _5833__289/A vssd1 vssd1 vccd1 vccd1 _7304_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3861_ _7527_/Q vssd1 vssd1 vccd1 vccd1 _4901_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6580_ _7095_/B _6670_/B _6670_/C vssd1 vssd1 vccd1 vccd1 _6580_/X sky130_fd_sc_hd__and3_1
X_5600_ _5598_/X _5599_/X _5611_/S vssd1 vssd1 vccd1 vccd1 _5600_/X sky130_fd_sc_hd__mux2_2
X_3792_ _7527_/Q _7522_/Q vssd1 vssd1 vccd1 vccd1 _4303_/C sky130_fd_sc_hd__xnor2_1
X_5531_ _7691_/Q _7280_/Q _7163_/Q _7272_/Q _5426_/A _4300_/A vssd1 vssd1 vccd1 vccd1
+ _5531_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_1_1_0__3292_ clkbuf_0__3292_/X vssd1 vssd1 vccd1 vccd1 _6736__129/A sky130_fd_sc_hd__clkbuf_4
X_7201_ _7329_/CLK _7201_/D vssd1 vssd1 vccd1 vccd1 _7201_/Q sky130_fd_sc_hd__dfxtp_1
X_5462_ _5462_/A _5462_/B _5493_/B _5462_/D vssd1 vssd1 vccd1 vccd1 _5495_/A sky130_fd_sc_hd__or4_1
XFILLER_99_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5393_ _7040_/B _5436_/A vssd1 vssd1 vccd1 vccd1 _5394_/C sky130_fd_sc_hd__or2_1
X_4413_ _4413_/A vssd1 vssd1 vccd1 vccd1 _7480_/D sky130_fd_sc_hd__clkbuf_1
X_7132_ _7224_/CLK _7132_/D vssd1 vssd1 vccd1 vccd1 _7132_/Q sky130_fd_sc_hd__dfxtp_1
X_4344_ _4344_/A vssd1 vssd1 vccd1 vccd1 _7508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7063_ _7063_/A vssd1 vssd1 vccd1 vccd1 _7843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6807__9 _6807__9/A vssd1 vssd1 vccd1 vccd1 _7751_/CLK sky130_fd_sc_hd__inv_2
X_6014_ _6031_/A vssd1 vssd1 vccd1 vccd1 _6014_/X sky130_fd_sc_hd__buf_2
X_4275_ _4901_/A _6308_/B _4278_/B _4979_/S vssd1 vssd1 vccd1 vccd1 _7527_/D sky130_fd_sc_hd__a31o_1
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2390_ clkbuf_0__2390_/X vssd1 vssd1 vccd1 vccd1 _5382_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6916_ _6916_/A _6916_/B vssd1 vssd1 vccd1 vccd1 _6972_/B sky130_fd_sc_hd__and2_1
XFILLER_35_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5729_ _5729_/A vssd1 vssd1 vccd1 vccd1 _7224_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6535__97 _6535__97/A vssd1 vssd1 vccd1 vccd1 _7642_/CLK sky130_fd_sc_hd__inv_2
X_5384__210 _5385__211/A vssd1 vssd1 vccd1 vccd1 _7182_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6853__46 _6855__48/A vssd1 vssd1 vccd1 vccd1 _7788_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4060_ _7825_/Q vssd1 vssd1 vccd1 vccd1 _4060_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7750_ _7750_/CLK _7750_/D vssd1 vssd1 vccd1 vccd1 _7750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4962_ _4962_/A vssd1 vssd1 vccd1 vccd1 _7165_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7681_ _7685_/CLK _7681_/D vssd1 vssd1 vccd1 vccd1 _7681_/Q sky130_fd_sc_hd__dfxtp_1
X_6701_ _6679_/X _6684_/X _7680_/Q vssd1 vssd1 vccd1 vccd1 _6701_/X sky130_fd_sc_hd__a21bo_1
Xclkbuf_0__2760_ _5740_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2760_/X sky130_fd_sc_hd__clkbuf_16
X_4893_ _4817_/X _7240_/Q _4893_/S vssd1 vssd1 vccd1 vccd1 _4894_/A sky130_fd_sc_hd__mux2_1
X_3913_ _3913_/A vssd1 vssd1 vccd1 vccd1 _7667_/D sky130_fd_sc_hd__clkbuf_1
X_6632_ _6668_/B vssd1 vssd1 vccd1 vccd1 _6725_/C sky130_fd_sc_hd__inv_2
X_3844_ _3859_/S vssd1 vssd1 vccd1 vccd1 _3853_/S sky130_fd_sc_hd__buf_2
X_6563_ _7681_/Q _6594_/A _6621_/C _6617_/D vssd1 vssd1 vccd1 vccd1 _6609_/B sky130_fd_sc_hd__and4_1
X_3775_ _3712_/X _7724_/Q _3775_/S vssd1 vssd1 vccd1 vccd1 _3776_/A sky130_fd_sc_hd__mux2_1
X_5514_ _7581_/Q _7565_/Q _7549_/Q _7541_/Q _5512_/X _5513_/X vssd1 vssd1 vccd1 vccd1
+ _5514_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3312_ _6832_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3312_/X sky130_fd_sc_hd__clkbuf_16
X_5445_ _5679_/A _5679_/B vssd1 vssd1 vccd1 vccd1 _7040_/A sky130_fd_sc_hd__or2b_1
X_7115_ _7115_/CLK _7115_/D vssd1 vssd1 vccd1 vccd1 _7115_/Q sky130_fd_sc_hd__dfxtp_1
X_5376_ _5376_/A vssd1 vssd1 vccd1 vccd1 _5376_/X sky130_fd_sc_hd__buf_1
XFILLER_113_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6784__165 _6788__169/A vssd1 vssd1 vccd1 vccd1 _7732_/CLK sky130_fd_sc_hd__inv_2
X_4327_ _4158_/X _7515_/Q _4331_/S vssd1 vssd1 vccd1 vccd1 _4328_/A sky130_fd_sc_hd__mux2_1
X_7046_ _5680_/A _7046_/B vssd1 vssd1 vccd1 vccd1 _7047_/A sky130_fd_sc_hd__and2b_1
X_4258_ _4258_/A vssd1 vssd1 vccd1 vccd1 _7534_/D sky130_fd_sc_hd__clkbuf_1
X_6170__372 _6172__374/A vssd1 vssd1 vccd1 vccd1 _7424_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6131__345 _6133__347/A vssd1 vssd1 vccd1 vccd1 _7394_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5773__241 _5775__243/A vssd1 vssd1 vccd1 vccd1 _7258_/CLK sky130_fd_sc_hd__inv_2
X_4189_ _4189_/A vssd1 vssd1 vccd1 vccd1 _7557_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7889__216 vssd1 vssd1 vccd1 vccd1 _7889__216/HI manufacturerID[8] sky130_fd_sc_hd__conb_1
XFILLER_19_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3560_ _3560_/A vssd1 vssd1 vccd1 vccd1 _7835_/D sky130_fd_sc_hd__clkbuf_1
X_6508__75 _6510__77/A vssd1 vssd1 vccd1 vccd1 _7620_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5230_ _5200_/X _5230_/B vssd1 vssd1 vccd1 vccd1 _5230_/X sky130_fd_sc_hd__and2b_1
X_5161_ _7188_/Q _5161_/B _5171_/C vssd1 vssd1 vccd1 vccd1 _5161_/X sky130_fd_sc_hd__and3_1
XFILLER_68_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5092_ _5092_/A _5098_/B vssd1 vssd1 vccd1 vccd1 _5093_/A sky130_fd_sc_hd__and2_1
XFILLER_68_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4112_ _4394_/B _4901_/C _4394_/A vssd1 vssd1 vccd1 vccd1 _4217_/B sky130_fd_sc_hd__and3b_4
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4043_ _4043_/A vssd1 vssd1 vccd1 vccd1 _7612_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5994_ _5932_/X _5977_/X _5992_/X _5993_/X vssd1 vssd1 vccd1 vccd1 _5994_/X sky130_fd_sc_hd__a211o_2
X_7802_ _7802_/CLK _7802_/D vssd1 vssd1 vccd1 vccd1 _7802_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__2775_ clkbuf_0__2775_/X vssd1 vssd1 vccd1 vccd1 _5825__284/A sky130_fd_sc_hd__clkbuf_4
X_7733_ _7733_/CLK _7733_/D vssd1 vssd1 vccd1 vccd1 _7733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4945_ _4227_/X _7172_/Q _4947_/S vssd1 vssd1 vccd1 vccd1 _4946_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4876_ _4876_/A vssd1 vssd1 vccd1 vccd1 _7248_/D sky130_fd_sc_hd__clkbuf_1
X_7664_ _7664_/CLK _7664_/D vssd1 vssd1 vccd1 vccd1 _7664_/Q sky130_fd_sc_hd__dfxtp_1
X_6615_ _6615_/A _6615_/B vssd1 vssd1 vccd1 vccd1 _6702_/B sky130_fd_sc_hd__nand2_1
X_3827_ _7471_/Q vssd1 vssd1 vccd1 vccd1 _4408_/A sky130_fd_sc_hd__buf_2
X_7595_ _7595_/CLK _7595_/D vssd1 vssd1 vccd1 vccd1 _7595_/Q sky130_fd_sc_hd__dfxtp_1
X_3758_ _3715_/X _7731_/Q _3762_/S vssd1 vssd1 vccd1 vccd1 _3759_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3689_ _3689_/A vssd1 vssd1 vccd1 vccd1 _7757_/D sky130_fd_sc_hd__clkbuf_1
X_5428_ _7301_/Q _7229_/Q _7697_/Q _7317_/Q _5426_/X _5427_/X vssd1 vssd1 vccd1 vccd1
+ _5428_/X sky130_fd_sc_hd__mux4_1
XFILLER_102_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_2 _7096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7029_ _7029_/A vssd1 vssd1 vccd1 vccd1 _7828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3088_ _6294_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3088_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_55_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6404__472 _6404__472/A vssd1 vssd1 vccd1 vccd1 _7537_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6177__378 _6177__378/A vssd1 vssd1 vccd1 vccd1 _7430_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6728__122 _6730__124/A vssd1 vssd1 vccd1 vccd1 _7688_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6446__506 _6448__508/A vssd1 vssd1 vccd1 vccd1 _7571_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4730_ _4730_/A vssd1 vssd1 vccd1 vccd1 _7309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4661_ _4661_/A vssd1 vssd1 vccd1 vccd1 _7360_/D sky130_fd_sc_hd__clkbuf_1
X_7380_ _7380_/CLK _7380_/D vssd1 vssd1 vccd1 vccd1 _7380_/Q sky130_fd_sc_hd__dfxtp_1
X_3612_ _4668_/A _3653_/B vssd1 vssd1 vccd1 vccd1 _3628_/S sky130_fd_sc_hd__nand2_2
X_4592_ _7398_/Q _3947_/A _4594_/S vssd1 vssd1 vccd1 vccd1 _4593_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3112_ clkbuf_0__3112_/X vssd1 vssd1 vccd1 vccd1 _6378__454/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3543_ _7465_/Q _3535_/A _4424_/B _4448_/B vssd1 vssd1 vccd1 vccd1 _3543_/X sky130_fd_sc_hd__a31o_1
Xclkbuf_0__2390_ _5247_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2390_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_89_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6262_ _6262_/A vssd1 vssd1 vccd1 vccd1 _7432_/D sky130_fd_sc_hd__clkbuf_1
X_5213_ _5206_/X _5213_/B vssd1 vssd1 vccd1 vccd1 _5213_/X sky130_fd_sc_hd__and2b_1
XFILLER_103_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6193_ _7807_/Q _6193_/B vssd1 vssd1 vccd1 vccd1 _6194_/A sky130_fd_sc_hd__xnor2_1
X_5144_ _5144_/A vssd1 vssd1 vccd1 vccd1 _5187_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5075_ _5075_/A _5077_/B vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__or2_1
XFILLER_111_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4026_ _3950_/X _7619_/Q _4026_/S vssd1 vssd1 vccd1 vccd1 _4027_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5977_ _5972_/X _5973_/X _5975_/X _5976_/X _5945_/X _5947_/X vssd1 vssd1 vccd1 vccd1
+ _5977_/X sky130_fd_sc_hd__mux4_2
XFILLER_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4928_ _4928_/A vssd1 vssd1 vccd1 vccd1 _7180_/D sky130_fd_sc_hd__clkbuf_1
X_7716_ _7716_/CLK _7716_/D vssd1 vssd1 vccd1 vccd1 _7716_/Q sky130_fd_sc_hd__dfxtp_1
X_7647_ _7647_/CLK _7647_/D vssd1 vssd1 vccd1 vccd1 _7647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4859_ _4820_/X _7255_/Q _4863_/S vssd1 vssd1 vccd1 vccd1 _4860_/A sky130_fd_sc_hd__mux2_1
X_7578_ _7578_/CLK _7578_/D vssd1 vssd1 vccd1 vccd1 _7578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6452__510 _6455__513/A vssd1 vssd1 vccd1 vccd1 _7575_/CLK sky130_fd_sc_hd__inv_2
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6741__130 _6743__132/A vssd1 vssd1 vccd1 vccd1 _7697_/CLK sky130_fd_sc_hd__inv_2
X_5900_ _7344_/Q _5073_/A _5902_/S vssd1 vssd1 vccd1 vccd1 _5901_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6880_ _7852_/Q _6880_/B vssd1 vssd1 vccd1 vccd1 _6882_/B sky130_fd_sc_hd__xnor2_1
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__2766_ clkbuf_0__2766_/X vssd1 vssd1 vccd1 vccd1 _5775__243/A sky130_fd_sc_hd__clkbuf_16
XFILLER_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_6_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7333_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4713_ _7473_/Q vssd1 vssd1 vccd1 vccd1 _4713_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7501_ _7501_/CLK _7501_/D vssd1 vssd1 vccd1 vccd1 _7501_/Q sky130_fd_sc_hd__dfxtp_1
X_5693_ _5693_/A vssd1 vssd1 vccd1 vccd1 _7208_/D sky130_fd_sc_hd__clkbuf_1
X_4644_ _3669_/X _7375_/Q _4648_/S vssd1 vssd1 vccd1 vccd1 _4645_/A sky130_fd_sc_hd__mux2_1
X_7432_ _7799_/CLK _7432_/D vssd1 vssd1 vccd1 vccd1 _7432_/Q sky130_fd_sc_hd__dfxtp_1
X_4575_ _4575_/A vssd1 vssd1 vccd1 vccd1 _7409_/D sky130_fd_sc_hd__clkbuf_1
X_7363_ _7363_/CLK _7363_/D vssd1 vssd1 vccd1 vccd1 _7363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3526_ _3927_/C vssd1 vssd1 vccd1 vccd1 _6325_/A sky130_fd_sc_hd__buf_2
X_6314_ _6314_/A vssd1 vssd1 vccd1 vccd1 _7470_/D sky130_fd_sc_hd__clkbuf_1
X_7294_ _7294_/CLK _7294_/D vssd1 vssd1 vccd1 vccd1 _7294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6245_ _6245_/A _6245_/B _6245_/C vssd1 vssd1 vccd1 vccd1 _6248_/B sky130_fd_sc_hd__nand3_2
XFILLER_69_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5127_ _7337_/Q _5131_/B vssd1 vssd1 vccd1 vccd1 _5128_/A sky130_fd_sc_hd__and2_1
XFILLER_29_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5058_ _5058_/A _5066_/B vssd1 vssd1 vccd1 vccd1 _5059_/A sky130_fd_sc_hd__or2_1
Xclkbuf_1_0_0__3311_ clkbuf_0__3311_/X vssd1 vssd1 vccd1 vccd1 _6831__29/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4009_ _4009_/A _4009_/B _3745_/A vssd1 vssd1 vccd1 vccd1 _4072_/B sky130_fd_sc_hd__or3b_2
XFILLER_38_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6487__58 _6488__59/A vssd1 vssd1 vccd1 vccd1 _7603_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6296__406 _6298__408/A vssd1 vssd1 vccd1 vccd1 _7459_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6376__452 _6376__452/A vssd1 vssd1 vccd1 vccd1 _7515_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4360_ _4360_/A vssd1 vssd1 vccd1 vccd1 _7501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _4291_/A vssd1 vssd1 vccd1 vccd1 _5433_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_98_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6030_ _6016_/A _6027_/X _6029_/X _5959_/A vssd1 vssd1 vccd1 vccd1 _6030_/X sky130_fd_sc_hd__o211a_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6932_ _6930_/Y _6931_/X _7014_/A vssd1 vssd1 vccd1 vccd1 _7799_/D sky130_fd_sc_hd__a21oi_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6863_ _6860_/Y _6861_/X _6862_/X _6250_/C _6250_/B vssd1 vssd1 vccd1 vccd1 _6867_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5814_ _5814_/A vssd1 vssd1 vccd1 vccd1 _5814_/X sky130_fd_sc_hd__buf_1
XFILLER_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6459__516 _6459__516/A vssd1 vssd1 vccd1 vccd1 _7581_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5676_ _7839_/Q _5676_/B vssd1 vssd1 vccd1 vccd1 _6326_/B sky130_fd_sc_hd__nand2_1
XFILLER_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7415_ _7415_/CLK _7415_/D vssd1 vssd1 vccd1 vccd1 _7415_/Q sky130_fd_sc_hd__dfxtp_1
X_4627_ _4627_/A vssd1 vssd1 vccd1 vccd1 _7383_/D sky130_fd_sc_hd__clkbuf_1
X_7346_ _7348_/CLK _7346_/D vssd1 vssd1 vccd1 vccd1 _7346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4558_ _4265_/X _7416_/Q _4558_/S vssd1 vssd1 vccd1 vccd1 _4559_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3509_ _4009_/A _3745_/A _4009_/B vssd1 vssd1 vccd1 vccd1 _4243_/A sky130_fd_sc_hd__or3b_1
X_6748__136 _6749__137/A vssd1 vssd1 vccd1 vccd1 _7703_/CLK sky130_fd_sc_hd__inv_2
X_4489_ _4393_/X _7448_/Q _4497_/S vssd1 vssd1 vccd1 vccd1 _4490_/A sky130_fd_sc_hd__mux2_1
X_7277_ _7277_/CLK _7277_/D vssd1 vssd1 vccd1 vccd1 _7277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6228_ _7799_/Q _6228_/B vssd1 vssd1 vccd1 vccd1 _6890_/B sky130_fd_sc_hd__xnor2_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5737__212 _5739__214/A vssd1 vssd1 vccd1 vccd1 _7229_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3087_ clkbuf_0__3087_/X vssd1 vssd1 vccd1 vccd1 _6292__403/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput95 _5108_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[11] sky130_fd_sc_hd__buf_2
XFILLER_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3860_ _3860_/A vssd1 vssd1 vccd1 vccd1 _7705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3791_ _3907_/B _3791_/B vssd1 vssd1 vccd1 vccd1 _4271_/A sky130_fd_sc_hd__and2_1
XFILLER_31_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5530_ _7296_/Q _7288_/Q _7264_/Q _7112_/Q _5502_/X _5416_/A vssd1 vssd1 vccd1 vccd1
+ _5530_/X sky130_fd_sc_hd__mux4_1
X_5461_ _5461_/A vssd1 vssd1 vccd1 vccd1 _5461_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7200_ _7407_/CLK _7200_/D vssd1 vssd1 vccd1 vccd1 _7200_/Q sky130_fd_sc_hd__dfxtp_1
X_4412_ _4411_/X _7480_/Q _4418_/S vssd1 vssd1 vccd1 vccd1 _4413_/A sky130_fd_sc_hd__mux2_1
X_5392_ _7204_/Q _5493_/A _5493_/B _5491_/A vssd1 vssd1 vccd1 vccd1 _5436_/A sky130_fd_sc_hd__or4_1
XFILLER_113_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7131_ _7372_/CLK _7131_/D vssd1 vssd1 vccd1 vccd1 _7131_/Q sky130_fd_sc_hd__dfxtp_1
X_4343_ _4155_/X _7508_/Q _4349_/S vssd1 vssd1 vccd1 vccd1 _4344_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7062_ _7106_/A _7062_/B vssd1 vssd1 vccd1 vccd1 _7063_/A sky130_fd_sc_hd__or2_1
X_4274_ _4987_/S vssd1 vssd1 vccd1 vccd1 _4979_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_113_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6013_ _7458_/Q vssd1 vssd1 vccd1 vccd1 _6013_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_86_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6915_ _6911_/A _6900_/Y _6914_/X vssd1 vssd1 vccd1 vccd1 _7795_/D sky130_fd_sc_hd__a21oi_1
X_6777_ _6783_/A vssd1 vssd1 vccd1 vccd1 _6777_/X sky130_fd_sc_hd__buf_1
XFILLER_23_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5728_ _7224_/Q _7339_/Q _6148_/S vssd1 vssd1 vccd1 vccd1 _5729_/A sky130_fd_sc_hd__mux2_1
X_3989_ _7635_/Q _3675_/X _3989_/S vssd1 vssd1 vccd1 vccd1 _3990_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5659_ _5667_/A _5659_/B vssd1 vssd1 vccd1 vccd1 _5660_/A sky130_fd_sc_hd__or2_1
XFILLER_117_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7329_ _7329_/CLK _7329_/D vssd1 vssd1 vccd1 vccd1 _7329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3139_ clkbuf_0__3139_/X vssd1 vssd1 vccd1 vccd1 _6512__79/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7685_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4961_ _4224_/X _7165_/Q _4965_/S vssd1 vssd1 vccd1 vccd1 _4962_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7680_ _7680_/CLK _7680_/D vssd1 vssd1 vccd1 vccd1 _7680_/Q sky130_fd_sc_hd__dfxtp_1
X_6700_ _6698_/Y _6699_/X _5970_/X vssd1 vssd1 vccd1 vccd1 _7679_/D sky130_fd_sc_hd__o21a_1
X_4892_ _4892_/A vssd1 vssd1 vccd1 vccd1 _7241_/D sky130_fd_sc_hd__clkbuf_1
X_3912_ _3816_/X _7667_/Q _3918_/S vssd1 vssd1 vccd1 vccd1 _3913_/A sky130_fd_sc_hd__mux2_1
X_6631_ _6668_/B _6631_/B _6630_/X vssd1 vssd1 vccd1 vccd1 _6634_/B sky130_fd_sc_hd__or3b_1
X_3843_ _4668_/A _4523_/B vssd1 vssd1 vccd1 vccd1 _3859_/S sky130_fd_sc_hd__nand2_2
X_6562_ _7680_/Q _7679_/Q _7678_/Q _7677_/Q vssd1 vssd1 vccd1 vccd1 _6617_/D sky130_fd_sc_hd__and4_1
X_3774_ _3774_/A vssd1 vssd1 vccd1 vccd1 _7725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5513_ _5521_/A vssd1 vssd1 vccd1 vccd1 _5513_/X sky130_fd_sc_hd__buf_2
Xclkbuf_0__3311_ _6826_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3311_/X sky130_fd_sc_hd__clkbuf_16
X_5444_ _7227_/Q vssd1 vssd1 vccd1 vccd1 _5679_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7114_ _7114_/CLK _7114_/D vssd1 vssd1 vccd1 vccd1 _7114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4326_ _4326_/A vssd1 vssd1 vccd1 vccd1 _7516_/D sky130_fd_sc_hd__clkbuf_1
X_4257_ _4256_/X _7534_/Q _4257_/S vssd1 vssd1 vccd1 vccd1 _4258_/A sky130_fd_sc_hd__mux2_1
X_7045_ _5049_/A _7839_/Q _7045_/S vssd1 vssd1 vccd1 vccd1 _7046_/B sky130_fd_sc_hd__mux2_1
X_6389__462 _6389__462/A vssd1 vssd1 vccd1 vccd1 _7525_/CLK sky130_fd_sc_hd__inv_2
X_4188_ _4063_/X _7557_/Q _4192_/S vssd1 vssd1 vccd1 vccd1 _4189_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2989_ clkbuf_0__2989_/X vssd1 vssd1 vccd1 vccd1 _6141__354/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5849__302 _5849__302/A vssd1 vssd1 vccd1 vccd1 _7319_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5160_ _5236_/B vssd1 vssd1 vccd1 vccd1 _5171_/C sky130_fd_sc_hd__clkbuf_1
X_5091_ _5091_/A vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__clkbuf_1
X_4111_ _4111_/A vssd1 vssd1 vccd1 vccd1 _4901_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_4042_ _3947_/X _7612_/Q _4044_/S vssd1 vssd1 vccd1 vccd1 _4043_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5993_ _5993_/A vssd1 vssd1 vccd1 vccd1 _5993_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7801_ _7802_/CLK _7801_/D vssd1 vssd1 vccd1 vccd1 _7801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__2774_ clkbuf_0__2774_/X vssd1 vssd1 vccd1 vccd1 _5818__278/A sky130_fd_sc_hd__clkbuf_4
X_7732_ _7732_/CLK _7732_/D vssd1 vssd1 vccd1 vccd1 _7732_/Q sky130_fd_sc_hd__dfxtp_1
X_4944_ _4944_/A vssd1 vssd1 vccd1 vccd1 _7173_/D sky130_fd_sc_hd__clkbuf_1
X_4875_ _7248_/Q _4408_/A _4875_/S vssd1 vssd1 vccd1 vccd1 _4876_/A sky130_fd_sc_hd__mux2_1
X_7663_ _7663_/CLK _7663_/D vssd1 vssd1 vccd1 vccd1 _7663_/Q sky130_fd_sc_hd__dfxtp_1
X_6614_ _7679_/Q _6621_/B _6621_/C _6621_/D _7680_/Q vssd1 vssd1 vccd1 vccd1 _6615_/B
+ sky130_fd_sc_hd__a41o_1
X_7594_ _7594_/CLK _7594_/D vssd1 vssd1 vccd1 vccd1 _7594_/Q sky130_fd_sc_hd__dfxtp_1
X_3826_ _3826_/A vssd1 vssd1 vccd1 vccd1 _7717_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__2990_ clkbuf_0__2990_/X vssd1 vssd1 vccd1 vccd1 _6153__359/A sky130_fd_sc_hd__clkbuf_4
X_6790__170 _6792__172/A vssd1 vssd1 vccd1 vccd1 _7737_/CLK sky130_fd_sc_hd__inv_2
X_3757_ _3757_/A vssd1 vssd1 vccd1 vccd1 _7732_/D sky130_fd_sc_hd__clkbuf_1
X_6545_ _6551_/A vssd1 vssd1 vccd1 vccd1 _6545_/X sky130_fd_sc_hd__buf_1
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5844__298 _5845__299/A vssd1 vssd1 vccd1 vccd1 _7315_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3688_ _3562_/X _7757_/Q _3690_/S vssd1 vssd1 vccd1 vccd1 _3689_/A sky130_fd_sc_hd__mux2_1
X_5427_ _5427_/A vssd1 vssd1 vccd1 vccd1 _5427_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_114_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5358_ _5358_/A vssd1 vssd1 vccd1 vccd1 _5358_/X sky130_fd_sc_hd__buf_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_3 _3824_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4309_ _5434_/A _4310_/B _4308_/Y vssd1 vssd1 vccd1 vccd1 _7522_/D sky130_fd_sc_hd__o21a_1
XFILLER_101_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5289_ _5287_/X _7330_/Q _5283_/X _5284_/X _7130_/Q vssd1 vssd1 vccd1 vccd1 _7130_/D
+ sky130_fd_sc_hd__o32a_1
X_7028_ _7028_/A _7030_/B vssd1 vssd1 vccd1 vccd1 _7029_/A sky130_fd_sc_hd__and2_1
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3087_ _6288_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3087_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_90_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6370__447 _6371__448/A vssd1 vssd1 vccd1 vccd1 _7510_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _4408_/X _7360_/Q _4660_/S vssd1 vssd1 vccd1 vccd1 _4661_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3611_ _3630_/D _4434_/A _4578_/A vssd1 vssd1 vccd1 vccd1 _4668_/A sky130_fd_sc_hd__and3b_4
X_4591_ _4591_/A vssd1 vssd1 vccd1 vccd1 _7399_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3111_ clkbuf_0__3111_/X vssd1 vssd1 vccd1 vccd1 _6371__448/A sky130_fd_sc_hd__clkbuf_4
X_6330_ _6348_/A vssd1 vssd1 vccd1 vccd1 _6330_/X sky130_fd_sc_hd__buf_1
X_3542_ _3927_/A _4447_/A _3541_/X vssd1 vssd1 vccd1 vccd1 _3542_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_115_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6261_ _7003_/A _6983_/A vssd1 vssd1 vccd1 vccd1 _6262_/A sky130_fd_sc_hd__and2_1
X_5212_ _7138_/Q _5199_/X _5204_/X _5211_/X vssd1 vssd1 vccd1 vccd1 _5212_/X sky130_fd_sc_hd__o22a_4
X_6192_ _6228_/B _6197_/A _6192_/C vssd1 vssd1 vccd1 vccd1 _6193_/B sky130_fd_sc_hd__and3_1
X_5143_ _5143_/A vssd1 vssd1 vccd1 vccd1 _5143_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5074_ _5074_/A vssd1 vssd1 vccd1 vccd1 _5074_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4025_ _4025_/A vssd1 vssd1 vccd1 vccd1 _7620_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5976_ _7572_/Q _7382_/Q _7730_/Q _7628_/Q _5942_/X _4465_/X vssd1 vssd1 vccd1 vccd1
+ _5976_/X sky130_fd_sc_hd__mux4_1
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4927_ _4227_/X _7180_/Q _4929_/S vssd1 vssd1 vccd1 vccd1 _4928_/A sky130_fd_sc_hd__mux2_1
X_7715_ _7715_/CLK _7715_/D vssd1 vssd1 vccd1 vccd1 _7715_/Q sky130_fd_sc_hd__dfxtp_1
X_7646_ _7646_/CLK _7646_/D vssd1 vssd1 vccd1 vccd1 _7646_/Q sky130_fd_sc_hd__dfxtp_1
X_4858_ _4858_/A vssd1 vssd1 vccd1 vccd1 _7256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3809_ _7527_/Q vssd1 vssd1 vccd1 vccd1 _4394_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3309_ clkbuf_0__3309_/X vssd1 vssd1 vccd1 vccd1 _6819__19/A sky130_fd_sc_hd__clkbuf_4
X_4789_ _4710_/X _7283_/Q _4795_/S vssd1 vssd1 vccd1 vccd1 _4790_/A sky130_fd_sc_hd__mux2_1
X_7577_ _7577_/CLK _7577_/D vssd1 vssd1 vccd1 vccd1 _7577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3139_ _6507_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3139_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6797__176 _6798__177/A vssd1 vssd1 vccd1 vccd1 _7743_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5786__252 _5788__254/A vssd1 vssd1 vccd1 vccd1 _7269_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7500_ _7500_/CLK _7500_/D vssd1 vssd1 vccd1 vccd1 _7500_/Q sky130_fd_sc_hd__dfxtp_1
X_4712_ _4712_/A vssd1 vssd1 vccd1 vccd1 _7315_/D sky130_fd_sc_hd__clkbuf_1
X_7431_ _7431_/CLK _7431_/D vssd1 vssd1 vccd1 vccd1 _7431_/Q sky130_fd_sc_hd__dfxtp_1
X_5692_ _7208_/Q _5096_/A _5692_/S vssd1 vssd1 vccd1 vccd1 _5693_/A sky130_fd_sc_hd__mux2_1
X_4643_ _4643_/A vssd1 vssd1 vccd1 vccd1 _7376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4574_ _4262_/X _7409_/Q _4576_/S vssd1 vssd1 vccd1 vccd1 _4575_/A sky130_fd_sc_hd__mux2_1
X_7362_ _7362_/CLK _7362_/D vssd1 vssd1 vccd1 vccd1 _7362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3525_ _3587_/A _3588_/A _3589_/A vssd1 vssd1 vccd1 vccd1 _3927_/C sky130_fd_sc_hd__a21o_1
X_6313_ _7816_/Q _6319_/B vssd1 vssd1 vccd1 vccd1 _6314_/A sky130_fd_sc_hd__and2_1
X_7293_ _7293_/CLK _7293_/D vssd1 vssd1 vccd1 vccd1 _7293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6244_ _7804_/Q vssd1 vssd1 vccd1 vccd1 _6244_/Y sky130_fd_sc_hd__inv_2
X_5126_ _5126_/A vssd1 vssd1 vccd1 vccd1 _5126_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5057_ _5068_/A vssd1 vssd1 vccd1 vccd1 _5066_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3310_ clkbuf_0__3310_/X vssd1 vssd1 vccd1 vccd1 _6822__21/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4008_ _4008_/A vssd1 vssd1 vccd1 vccd1 _7627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5959_ _5959_/A vssd1 vssd1 vccd1 vccd1 _5959_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7629_ _7629_/CLK _7629_/D vssd1 vssd1 vccd1 vccd1 _7629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6417__483 _6417__483/A vssd1 vssd1 vccd1 vccd1 _7548_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4290_ _5403_/A vssd1 vssd1 vccd1 vccd1 _4291_/A sky130_fd_sc_hd__buf_2
XFILLER_112_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2990_ _6142_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2990_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6931_ _6924_/X _6907_/X _6890_/B vssd1 vssd1 vccd1 vccd1 _6931_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6862_ _7848_/Q _6873_/B _6991_/B _6991_/A vssd1 vssd1 vccd1 vccd1 _6862_/X sky130_fd_sc_hd__o211a_1
XFILLER_50_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5675_ _7838_/Q vssd1 vssd1 vccd1 vccd1 _6901_/A sky130_fd_sc_hd__clkinv_4
X_7414_ _7414_/CLK _7414_/D vssd1 vssd1 vccd1 vccd1 _7414_/Q sky130_fd_sc_hd__dfxtp_1
X_4626_ _3669_/X _7383_/Q _4630_/S vssd1 vssd1 vccd1 vccd1 _4627_/A sky130_fd_sc_hd__mux2_1
X_7345_ _7348_/CLK _7345_/D vssd1 vssd1 vccd1 vccd1 _7345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4557_ _4557_/A vssd1 vssd1 vccd1 vccd1 _7417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3508_ _7465_/Q vssd1 vssd1 vccd1 vccd1 _4009_/B sky130_fd_sc_hd__clkbuf_1
X_7276_ _7276_/CLK _7276_/D vssd1 vssd1 vccd1 vccd1 _7276_/Q sky130_fd_sc_hd__dfxtp_1
X_4488_ _4503_/S vssd1 vssd1 vccd1 vccd1 _4497_/S sky130_fd_sc_hd__buf_2
X_6227_ _7852_/Q _6881_/B vssd1 vssd1 vccd1 vccd1 _6991_/C sky130_fd_sc_hd__xor2_1
XFILLER_106_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _5109_/A _5109_/B vssd1 vssd1 vccd1 vccd1 _5110_/A sky130_fd_sc_hd__and2_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _7760_/Q _7752_/Q _7744_/Q _7658_/Q _4465_/A _5954_/X vssd1 vssd1 vccd1 vccd1
+ _6089_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6492__62 _6492__62/A vssd1 vssd1 vccd1 vccd1 _7607_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7039__4 _7039__4/A vssd1 vssd1 vccd1 vccd1 _7837_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3086_ clkbuf_0__3086_/X vssd1 vssd1 vccd1 vccd1 _6286__398/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput96 _5110_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[12] sky130_fd_sc_hd__buf_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3790_ _7525_/Q _7524_/Q _7523_/Q vssd1 vssd1 vccd1 vccd1 _3791_/B sky130_fd_sc_hd__and3_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5460_ _7854_/Q _6326_/A _5457_/X _5459_/X vssd1 vssd1 vccd1 vccd1 _5460_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4411_ _4411_/A vssd1 vssd1 vccd1 vccd1 _4411_/X sky130_fd_sc_hd__clkbuf_2
X_5391_ _5679_/B _7227_/Q vssd1 vssd1 vccd1 vccd1 _5491_/A sky130_fd_sc_hd__or2b_1
XFILLER_98_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7130_ _7372_/CLK _7130_/D vssd1 vssd1 vccd1 vccd1 _7130_/Q sky130_fd_sc_hd__dfxtp_1
X_4342_ _4342_/A vssd1 vssd1 vccd1 vccd1 _7509_/D sky130_fd_sc_hd__clkbuf_1
X_5799__262 _5799__262/A vssd1 vssd1 vccd1 vccd1 _7279_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7061_ _5040_/A _6195_/A _7074_/S vssd1 vssd1 vccd1 vccd1 _7062_/B sky130_fd_sc_hd__mux2_1
X_4273_ _6310_/A _4284_/A _4829_/B vssd1 vssd1 vccd1 vccd1 _4987_/S sky130_fd_sc_hd__and3_4
X_6012_ _7410_/Q _7351_/Q _7418_/Q _7399_/Q _4446_/A _6011_/X vssd1 vssd1 vccd1 vccd1
+ _6012_/X sky130_fd_sc_hd__mux4_1
.ends

