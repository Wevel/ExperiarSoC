magic
tech sky130A
magscale 1 2
timestamp 1653063993
<< obsli1 >>
rect 1104 2159 68816 197489
<< obsm1 >>
rect 566 1708 69722 197520
<< metal2 >>
rect 294 199200 350 200000
rect 938 199200 994 200000
rect 1674 199200 1730 200000
rect 2410 199200 2466 200000
rect 3146 199200 3202 200000
rect 3790 199200 3846 200000
rect 4526 199200 4582 200000
rect 5262 199200 5318 200000
rect 5998 199200 6054 200000
rect 6642 199200 6698 200000
rect 7378 199200 7434 200000
rect 8114 199200 8170 200000
rect 8850 199200 8906 200000
rect 9494 199200 9550 200000
rect 10230 199200 10286 200000
rect 10966 199200 11022 200000
rect 11702 199200 11758 200000
rect 12438 199200 12494 200000
rect 13082 199200 13138 200000
rect 13818 199200 13874 200000
rect 14554 199200 14610 200000
rect 15290 199200 15346 200000
rect 15934 199200 15990 200000
rect 16670 199200 16726 200000
rect 17406 199200 17462 200000
rect 18142 199200 18198 200000
rect 18786 199200 18842 200000
rect 19522 199200 19578 200000
rect 20258 199200 20314 200000
rect 20994 199200 21050 200000
rect 21638 199200 21694 200000
rect 22374 199200 22430 200000
rect 23110 199200 23166 200000
rect 23846 199200 23902 200000
rect 24582 199200 24638 200000
rect 25226 199200 25282 200000
rect 25962 199200 26018 200000
rect 26698 199200 26754 200000
rect 27434 199200 27490 200000
rect 28078 199200 28134 200000
rect 28814 199200 28870 200000
rect 29550 199200 29606 200000
rect 30286 199200 30342 200000
rect 30930 199200 30986 200000
rect 31666 199200 31722 200000
rect 32402 199200 32458 200000
rect 33138 199200 33194 200000
rect 33782 199200 33838 200000
rect 34518 199200 34574 200000
rect 35254 199200 35310 200000
rect 35990 199200 36046 200000
rect 36726 199200 36782 200000
rect 37370 199200 37426 200000
rect 38106 199200 38162 200000
rect 38842 199200 38898 200000
rect 39578 199200 39634 200000
rect 40222 199200 40278 200000
rect 40958 199200 41014 200000
rect 41694 199200 41750 200000
rect 42430 199200 42486 200000
rect 43074 199200 43130 200000
rect 43810 199200 43866 200000
rect 44546 199200 44602 200000
rect 45282 199200 45338 200000
rect 45926 199200 45982 200000
rect 46662 199200 46718 200000
rect 47398 199200 47454 200000
rect 48134 199200 48190 200000
rect 48870 199200 48926 200000
rect 49514 199200 49570 200000
rect 50250 199200 50306 200000
rect 50986 199200 51042 200000
rect 51722 199200 51778 200000
rect 52366 199200 52422 200000
rect 53102 199200 53158 200000
rect 53838 199200 53894 200000
rect 54574 199200 54630 200000
rect 55218 199200 55274 200000
rect 55954 199200 56010 200000
rect 56690 199200 56746 200000
rect 57426 199200 57482 200000
rect 58070 199200 58126 200000
rect 58806 199200 58862 200000
rect 59542 199200 59598 200000
rect 60278 199200 60334 200000
rect 61014 199200 61070 200000
rect 61658 199200 61714 200000
rect 62394 199200 62450 200000
rect 63130 199200 63186 200000
rect 63866 199200 63922 200000
rect 64510 199200 64566 200000
rect 65246 199200 65302 200000
rect 65982 199200 66038 200000
rect 66718 199200 66774 200000
rect 67362 199200 67418 200000
rect 68098 199200 68154 200000
rect 68834 199200 68890 200000
rect 69570 199200 69626 200000
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 1950 0 2006 800
rect 2502 0 2558 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4710 0 4766 800
rect 5262 0 5318 800
rect 5814 0 5870 800
rect 6366 0 6422 800
rect 6918 0 6974 800
rect 7470 0 7526 800
rect 8022 0 8078 800
rect 8574 0 8630 800
rect 9126 0 9182 800
rect 9678 0 9734 800
rect 10230 0 10286 800
rect 10782 0 10838 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12438 0 12494 800
rect 12990 0 13046 800
rect 13542 0 13598 800
rect 14094 0 14150 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16394 0 16450 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
rect 23018 0 23074 800
rect 23570 0 23626 800
rect 24122 0 24178 800
rect 24674 0 24730 800
rect 25226 0 25282 800
rect 25778 0 25834 800
rect 26330 0 26386 800
rect 26882 0 26938 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28630 0 28686 800
rect 29182 0 29238 800
rect 29734 0 29790 800
rect 30286 0 30342 800
rect 30838 0 30894 800
rect 31390 0 31446 800
rect 31942 0 31998 800
rect 32494 0 32550 800
rect 33046 0 33102 800
rect 33598 0 33654 800
rect 34150 0 34206 800
rect 34702 0 34758 800
rect 35254 0 35310 800
rect 35806 0 35862 800
rect 36358 0 36414 800
rect 36910 0 36966 800
rect 37462 0 37518 800
rect 38014 0 38070 800
rect 38566 0 38622 800
rect 39118 0 39174 800
rect 39670 0 39726 800
rect 40222 0 40278 800
rect 40774 0 40830 800
rect 41326 0 41382 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43074 0 43130 800
rect 43626 0 43682 800
rect 44178 0 44234 800
rect 44730 0 44786 800
rect 45282 0 45338 800
rect 45834 0 45890 800
rect 46386 0 46442 800
rect 46938 0 46994 800
rect 47490 0 47546 800
rect 48042 0 48098 800
rect 48594 0 48650 800
rect 49146 0 49202 800
rect 49698 0 49754 800
rect 50250 0 50306 800
rect 50802 0 50858 800
rect 51354 0 51410 800
rect 51906 0 51962 800
rect 52458 0 52514 800
rect 53010 0 53066 800
rect 53562 0 53618 800
rect 54114 0 54170 800
rect 54666 0 54722 800
rect 55218 0 55274 800
rect 55770 0 55826 800
rect 56414 0 56470 800
rect 56966 0 57022 800
rect 57518 0 57574 800
rect 58070 0 58126 800
rect 58622 0 58678 800
rect 59174 0 59230 800
rect 59726 0 59782 800
rect 60278 0 60334 800
rect 60830 0 60886 800
rect 61382 0 61438 800
rect 61934 0 61990 800
rect 62486 0 62542 800
rect 63038 0 63094 800
rect 63590 0 63646 800
rect 64142 0 64198 800
rect 64694 0 64750 800
rect 65246 0 65302 800
rect 65798 0 65854 800
rect 66350 0 66406 800
rect 66902 0 66958 800
rect 67454 0 67510 800
rect 68006 0 68062 800
rect 68558 0 68614 800
rect 69110 0 69166 800
rect 69662 0 69718 800
<< obsm2 >>
rect 18 199144 238 199753
rect 406 199144 882 199753
rect 1050 199144 1618 199753
rect 1786 199144 2354 199753
rect 2522 199144 3090 199753
rect 3258 199144 3734 199753
rect 3902 199144 4470 199753
rect 4638 199144 5206 199753
rect 5374 199144 5942 199753
rect 6110 199144 6586 199753
rect 6754 199144 7322 199753
rect 7490 199144 8058 199753
rect 8226 199144 8794 199753
rect 8962 199144 9438 199753
rect 9606 199144 10174 199753
rect 10342 199144 10910 199753
rect 11078 199144 11646 199753
rect 11814 199144 12382 199753
rect 12550 199144 13026 199753
rect 13194 199144 13762 199753
rect 13930 199144 14498 199753
rect 14666 199144 15234 199753
rect 15402 199144 15878 199753
rect 16046 199144 16614 199753
rect 16782 199144 17350 199753
rect 17518 199144 18086 199753
rect 18254 199144 18730 199753
rect 18898 199144 19466 199753
rect 19634 199144 20202 199753
rect 20370 199144 20938 199753
rect 21106 199144 21582 199753
rect 21750 199144 22318 199753
rect 22486 199144 23054 199753
rect 23222 199144 23790 199753
rect 23958 199144 24526 199753
rect 24694 199144 25170 199753
rect 25338 199144 25906 199753
rect 26074 199144 26642 199753
rect 26810 199144 27378 199753
rect 27546 199144 28022 199753
rect 28190 199144 28758 199753
rect 28926 199144 29494 199753
rect 29662 199144 30230 199753
rect 30398 199144 30874 199753
rect 31042 199144 31610 199753
rect 31778 199144 32346 199753
rect 32514 199144 33082 199753
rect 33250 199144 33726 199753
rect 33894 199144 34462 199753
rect 34630 199144 35198 199753
rect 35366 199144 35934 199753
rect 36102 199144 36670 199753
rect 36838 199144 37314 199753
rect 37482 199144 38050 199753
rect 38218 199144 38786 199753
rect 38954 199144 39522 199753
rect 39690 199144 40166 199753
rect 40334 199144 40902 199753
rect 41070 199144 41638 199753
rect 41806 199144 42374 199753
rect 42542 199144 43018 199753
rect 43186 199144 43754 199753
rect 43922 199144 44490 199753
rect 44658 199144 45226 199753
rect 45394 199144 45870 199753
rect 46038 199144 46606 199753
rect 46774 199144 47342 199753
rect 47510 199144 48078 199753
rect 48246 199144 48814 199753
rect 48982 199144 49458 199753
rect 49626 199144 50194 199753
rect 50362 199144 50930 199753
rect 51098 199144 51666 199753
rect 51834 199144 52310 199753
rect 52478 199144 53046 199753
rect 53214 199144 53782 199753
rect 53950 199144 54518 199753
rect 54686 199144 55162 199753
rect 55330 199144 55898 199753
rect 56066 199144 56634 199753
rect 56802 199144 57370 199753
rect 57538 199144 58014 199753
rect 58182 199144 58750 199753
rect 58918 199144 59486 199753
rect 59654 199144 60222 199753
rect 60390 199144 60958 199753
rect 61126 199144 61602 199753
rect 61770 199144 62338 199753
rect 62506 199144 63074 199753
rect 63242 199144 63810 199753
rect 63978 199144 64454 199753
rect 64622 199144 65190 199753
rect 65358 199144 65926 199753
rect 66094 199144 66662 199753
rect 66830 199144 67306 199753
rect 67474 199144 68042 199753
rect 68210 199144 68778 199753
rect 68946 199144 69514 199753
rect 69682 199144 69716 199753
rect 18 856 69716 199144
rect 18 167 238 856
rect 406 167 790 856
rect 958 167 1342 856
rect 1510 167 1894 856
rect 2062 167 2446 856
rect 2614 167 2998 856
rect 3166 167 3550 856
rect 3718 167 4102 856
rect 4270 167 4654 856
rect 4822 167 5206 856
rect 5374 167 5758 856
rect 5926 167 6310 856
rect 6478 167 6862 856
rect 7030 167 7414 856
rect 7582 167 7966 856
rect 8134 167 8518 856
rect 8686 167 9070 856
rect 9238 167 9622 856
rect 9790 167 10174 856
rect 10342 167 10726 856
rect 10894 167 11278 856
rect 11446 167 11830 856
rect 11998 167 12382 856
rect 12550 167 12934 856
rect 13102 167 13486 856
rect 13654 167 14038 856
rect 14206 167 14682 856
rect 14850 167 15234 856
rect 15402 167 15786 856
rect 15954 167 16338 856
rect 16506 167 16890 856
rect 17058 167 17442 856
rect 17610 167 17994 856
rect 18162 167 18546 856
rect 18714 167 19098 856
rect 19266 167 19650 856
rect 19818 167 20202 856
rect 20370 167 20754 856
rect 20922 167 21306 856
rect 21474 167 21858 856
rect 22026 167 22410 856
rect 22578 167 22962 856
rect 23130 167 23514 856
rect 23682 167 24066 856
rect 24234 167 24618 856
rect 24786 167 25170 856
rect 25338 167 25722 856
rect 25890 167 26274 856
rect 26442 167 26826 856
rect 26994 167 27378 856
rect 27546 167 27930 856
rect 28098 167 28574 856
rect 28742 167 29126 856
rect 29294 167 29678 856
rect 29846 167 30230 856
rect 30398 167 30782 856
rect 30950 167 31334 856
rect 31502 167 31886 856
rect 32054 167 32438 856
rect 32606 167 32990 856
rect 33158 167 33542 856
rect 33710 167 34094 856
rect 34262 167 34646 856
rect 34814 167 35198 856
rect 35366 167 35750 856
rect 35918 167 36302 856
rect 36470 167 36854 856
rect 37022 167 37406 856
rect 37574 167 37958 856
rect 38126 167 38510 856
rect 38678 167 39062 856
rect 39230 167 39614 856
rect 39782 167 40166 856
rect 40334 167 40718 856
rect 40886 167 41270 856
rect 41438 167 41822 856
rect 41990 167 42466 856
rect 42634 167 43018 856
rect 43186 167 43570 856
rect 43738 167 44122 856
rect 44290 167 44674 856
rect 44842 167 45226 856
rect 45394 167 45778 856
rect 45946 167 46330 856
rect 46498 167 46882 856
rect 47050 167 47434 856
rect 47602 167 47986 856
rect 48154 167 48538 856
rect 48706 167 49090 856
rect 49258 167 49642 856
rect 49810 167 50194 856
rect 50362 167 50746 856
rect 50914 167 51298 856
rect 51466 167 51850 856
rect 52018 167 52402 856
rect 52570 167 52954 856
rect 53122 167 53506 856
rect 53674 167 54058 856
rect 54226 167 54610 856
rect 54778 167 55162 856
rect 55330 167 55714 856
rect 55882 167 56358 856
rect 56526 167 56910 856
rect 57078 167 57462 856
rect 57630 167 58014 856
rect 58182 167 58566 856
rect 58734 167 59118 856
rect 59286 167 59670 856
rect 59838 167 60222 856
rect 60390 167 60774 856
rect 60942 167 61326 856
rect 61494 167 61878 856
rect 62046 167 62430 856
rect 62598 167 62982 856
rect 63150 167 63534 856
rect 63702 167 64086 856
rect 64254 167 64638 856
rect 64806 167 65190 856
rect 65358 167 65742 856
rect 65910 167 66294 856
rect 66462 167 66846 856
rect 67014 167 67398 856
rect 67566 167 67950 856
rect 68118 167 68502 856
rect 68670 167 69054 856
rect 69222 167 69606 856
<< metal3 >>
rect 0 199656 800 199776
rect 69200 199384 70000 199504
rect 0 199112 800 199232
rect 0 198568 800 198688
rect 0 198160 800 198280
rect 69200 198296 70000 198416
rect 0 197616 800 197736
rect 69200 197344 70000 197464
rect 0 197072 800 197192
rect 0 196664 800 196784
rect 0 196120 800 196240
rect 69200 196256 70000 196376
rect 0 195576 800 195696
rect 0 195168 800 195288
rect 69200 195304 70000 195424
rect 0 194624 800 194744
rect 0 194080 800 194200
rect 69200 194216 70000 194336
rect 0 193672 800 193792
rect 0 193128 800 193248
rect 69200 193264 70000 193384
rect 0 192584 800 192704
rect 0 192176 800 192296
rect 69200 192176 70000 192296
rect 0 191632 800 191752
rect 0 191088 800 191208
rect 69200 191224 70000 191344
rect 0 190680 800 190800
rect 0 190136 800 190256
rect 69200 190136 70000 190256
rect 0 189592 800 189712
rect 0 189184 800 189304
rect 69200 189184 70000 189304
rect 0 188640 800 188760
rect 0 188096 800 188216
rect 69200 188096 70000 188216
rect 0 187688 800 187808
rect 0 187144 800 187264
rect 69200 187144 70000 187264
rect 0 186600 800 186720
rect 0 186192 800 186312
rect 69200 186056 70000 186176
rect 0 185648 800 185768
rect 0 185104 800 185224
rect 69200 185104 70000 185224
rect 0 184560 800 184680
rect 0 184152 800 184272
rect 69200 184016 70000 184136
rect 0 183608 800 183728
rect 0 183064 800 183184
rect 69200 183064 70000 183184
rect 0 182656 800 182776
rect 0 182112 800 182232
rect 69200 181976 70000 182096
rect 0 181568 800 181688
rect 0 181160 800 181280
rect 69200 181024 70000 181144
rect 0 180616 800 180736
rect 0 180072 800 180192
rect 69200 179936 70000 180056
rect 0 179664 800 179784
rect 0 179120 800 179240
rect 69200 178984 70000 179104
rect 0 178576 800 178696
rect 0 178168 800 178288
rect 69200 177896 70000 178016
rect 0 177624 800 177744
rect 0 177080 800 177200
rect 69200 176944 70000 177064
rect 0 176672 800 176792
rect 0 176128 800 176248
rect 69200 175856 70000 175976
rect 0 175584 800 175704
rect 0 175176 800 175296
rect 69200 174904 70000 175024
rect 0 174632 800 174752
rect 0 174088 800 174208
rect 0 173680 800 173800
rect 69200 173816 70000 173936
rect 0 173136 800 173256
rect 69200 172864 70000 172984
rect 0 172592 800 172712
rect 0 172184 800 172304
rect 0 171640 800 171760
rect 69200 171776 70000 171896
rect 0 171096 800 171216
rect 0 170688 800 170808
rect 69200 170824 70000 170944
rect 0 170144 800 170264
rect 0 169600 800 169720
rect 69200 169736 70000 169856
rect 0 169056 800 169176
rect 0 168648 800 168768
rect 69200 168784 70000 168904
rect 0 168104 800 168224
rect 0 167560 800 167680
rect 69200 167696 70000 167816
rect 0 167152 800 167272
rect 0 166608 800 166728
rect 69200 166744 70000 166864
rect 0 166064 800 166184
rect 0 165656 800 165776
rect 69200 165656 70000 165776
rect 0 165112 800 165232
rect 0 164568 800 164688
rect 69200 164704 70000 164824
rect 0 164160 800 164280
rect 0 163616 800 163736
rect 69200 163616 70000 163736
rect 0 163072 800 163192
rect 0 162664 800 162784
rect 69200 162664 70000 162784
rect 0 162120 800 162240
rect 0 161576 800 161696
rect 69200 161576 70000 161696
rect 0 161168 800 161288
rect 0 160624 800 160744
rect 69200 160624 70000 160744
rect 0 160080 800 160200
rect 0 159672 800 159792
rect 69200 159536 70000 159656
rect 0 159128 800 159248
rect 0 158584 800 158704
rect 69200 158584 70000 158704
rect 0 158176 800 158296
rect 0 157632 800 157752
rect 69200 157496 70000 157616
rect 0 157088 800 157208
rect 0 156680 800 156800
rect 69200 156544 70000 156664
rect 0 156136 800 156256
rect 0 155592 800 155712
rect 69200 155456 70000 155576
rect 0 155184 800 155304
rect 0 154640 800 154760
rect 69200 154504 70000 154624
rect 0 154096 800 154216
rect 0 153552 800 153672
rect 69200 153416 70000 153536
rect 0 153144 800 153264
rect 0 152600 800 152720
rect 69200 152464 70000 152584
rect 0 152056 800 152176
rect 0 151648 800 151768
rect 69200 151376 70000 151496
rect 0 151104 800 151224
rect 0 150560 800 150680
rect 69200 150424 70000 150544
rect 0 150152 800 150272
rect 0 149608 800 149728
rect 69200 149336 70000 149456
rect 0 149064 800 149184
rect 0 148656 800 148776
rect 69200 148384 70000 148504
rect 0 148112 800 148232
rect 0 147568 800 147688
rect 0 147160 800 147280
rect 69200 147296 70000 147416
rect 0 146616 800 146736
rect 69200 146344 70000 146464
rect 0 146072 800 146192
rect 0 145664 800 145784
rect 0 145120 800 145240
rect 69200 145256 70000 145376
rect 0 144576 800 144696
rect 0 144168 800 144288
rect 69200 144304 70000 144424
rect 0 143624 800 143744
rect 0 143080 800 143200
rect 69200 143216 70000 143336
rect 0 142672 800 142792
rect 0 142128 800 142248
rect 69200 142264 70000 142384
rect 0 141584 800 141704
rect 0 141176 800 141296
rect 69200 141176 70000 141296
rect 0 140632 800 140752
rect 0 140088 800 140208
rect 69200 140224 70000 140344
rect 0 139680 800 139800
rect 0 139136 800 139256
rect 69200 139136 70000 139256
rect 0 138592 800 138712
rect 0 138048 800 138168
rect 69200 138184 70000 138304
rect 0 137640 800 137760
rect 0 137096 800 137216
rect 69200 137096 70000 137216
rect 0 136552 800 136672
rect 0 136144 800 136264
rect 69200 136144 70000 136264
rect 0 135600 800 135720
rect 0 135056 800 135176
rect 69200 135056 70000 135176
rect 0 134648 800 134768
rect 0 134104 800 134224
rect 69200 134104 70000 134224
rect 0 133560 800 133680
rect 0 133152 800 133272
rect 69200 133016 70000 133136
rect 0 132608 800 132728
rect 0 132064 800 132184
rect 69200 132064 70000 132184
rect 0 131656 800 131776
rect 0 131112 800 131232
rect 69200 130976 70000 131096
rect 0 130568 800 130688
rect 0 130160 800 130280
rect 69200 130024 70000 130144
rect 0 129616 800 129736
rect 0 129072 800 129192
rect 69200 128936 70000 129056
rect 0 128664 800 128784
rect 0 128120 800 128240
rect 69200 127984 70000 128104
rect 0 127576 800 127696
rect 0 127168 800 127288
rect 69200 126896 70000 127016
rect 0 126624 800 126744
rect 0 126080 800 126200
rect 69200 125944 70000 126064
rect 0 125672 800 125792
rect 0 125128 800 125248
rect 69200 124856 70000 124976
rect 0 124584 800 124704
rect 0 124176 800 124296
rect 69200 123904 70000 124024
rect 0 123632 800 123752
rect 0 123088 800 123208
rect 69200 122816 70000 122936
rect 0 122544 800 122664
rect 0 122136 800 122256
rect 69200 121864 70000 121984
rect 0 121592 800 121712
rect 0 121048 800 121168
rect 0 120640 800 120760
rect 69200 120776 70000 120896
rect 0 120096 800 120216
rect 69200 119824 70000 119944
rect 0 119552 800 119672
rect 0 119144 800 119264
rect 0 118600 800 118720
rect 69200 118736 70000 118856
rect 0 118056 800 118176
rect 0 117648 800 117768
rect 69200 117784 70000 117904
rect 0 117104 800 117224
rect 0 116560 800 116680
rect 69200 116696 70000 116816
rect 0 116152 800 116272
rect 0 115608 800 115728
rect 69200 115744 70000 115864
rect 0 115064 800 115184
rect 0 114656 800 114776
rect 69200 114656 70000 114776
rect 0 114112 800 114232
rect 0 113568 800 113688
rect 69200 113704 70000 113824
rect 0 113160 800 113280
rect 0 112616 800 112736
rect 69200 112616 70000 112736
rect 0 112072 800 112192
rect 0 111664 800 111784
rect 69200 111664 70000 111784
rect 0 111120 800 111240
rect 0 110576 800 110696
rect 69200 110576 70000 110696
rect 0 110168 800 110288
rect 0 109624 800 109744
rect 69200 109624 70000 109744
rect 0 109080 800 109200
rect 0 108672 800 108792
rect 69200 108536 70000 108656
rect 0 108128 800 108248
rect 0 107584 800 107704
rect 69200 107584 70000 107704
rect 0 107040 800 107160
rect 0 106632 800 106752
rect 69200 106496 70000 106616
rect 0 106088 800 106208
rect 0 105544 800 105664
rect 69200 105544 70000 105664
rect 0 105136 800 105256
rect 0 104592 800 104712
rect 69200 104456 70000 104576
rect 0 104048 800 104168
rect 0 103640 800 103760
rect 69200 103504 70000 103624
rect 0 103096 800 103216
rect 0 102552 800 102672
rect 69200 102416 70000 102536
rect 0 102144 800 102264
rect 0 101600 800 101720
rect 69200 101464 70000 101584
rect 0 101056 800 101176
rect 0 100648 800 100768
rect 69200 100376 70000 100496
rect 0 100104 800 100224
rect 0 99560 800 99680
rect 0 99152 800 99272
rect 69200 99288 70000 99408
rect 0 98608 800 98728
rect 69200 98336 70000 98456
rect 0 98064 800 98184
rect 0 97656 800 97776
rect 0 97112 800 97232
rect 69200 97248 70000 97368
rect 0 96568 800 96688
rect 0 96160 800 96280
rect 69200 96296 70000 96416
rect 0 95616 800 95736
rect 0 95072 800 95192
rect 69200 95208 70000 95328
rect 0 94664 800 94784
rect 0 94120 800 94240
rect 69200 94256 70000 94376
rect 0 93576 800 93696
rect 0 93168 800 93288
rect 69200 93168 70000 93288
rect 0 92624 800 92744
rect 0 92080 800 92200
rect 69200 92216 70000 92336
rect 0 91536 800 91656
rect 0 91128 800 91248
rect 69200 91128 70000 91248
rect 0 90584 800 90704
rect 0 90040 800 90160
rect 69200 90176 70000 90296
rect 0 89632 800 89752
rect 0 89088 800 89208
rect 69200 89088 70000 89208
rect 0 88544 800 88664
rect 0 88136 800 88256
rect 69200 88136 70000 88256
rect 0 87592 800 87712
rect 0 87048 800 87168
rect 69200 87048 70000 87168
rect 0 86640 800 86760
rect 0 86096 800 86216
rect 69200 86096 70000 86216
rect 0 85552 800 85672
rect 0 85144 800 85264
rect 69200 85008 70000 85128
rect 0 84600 800 84720
rect 0 84056 800 84176
rect 69200 84056 70000 84176
rect 0 83648 800 83768
rect 0 83104 800 83224
rect 69200 82968 70000 83088
rect 0 82560 800 82680
rect 0 82152 800 82272
rect 69200 82016 70000 82136
rect 0 81608 800 81728
rect 0 81064 800 81184
rect 69200 80928 70000 81048
rect 0 80656 800 80776
rect 0 80112 800 80232
rect 69200 79976 70000 80096
rect 0 79568 800 79688
rect 0 79160 800 79280
rect 69200 78888 70000 79008
rect 0 78616 800 78736
rect 0 78072 800 78192
rect 69200 77936 70000 78056
rect 0 77664 800 77784
rect 0 77120 800 77240
rect 69200 76848 70000 76968
rect 0 76576 800 76696
rect 0 76032 800 76152
rect 69200 75896 70000 76016
rect 0 75624 800 75744
rect 0 75080 800 75200
rect 69200 74808 70000 74928
rect 0 74536 800 74656
rect 0 74128 800 74248
rect 69200 73856 70000 73976
rect 0 73584 800 73704
rect 0 73040 800 73160
rect 0 72632 800 72752
rect 69200 72768 70000 72888
rect 0 72088 800 72208
rect 69200 71816 70000 71936
rect 0 71544 800 71664
rect 0 71136 800 71256
rect 0 70592 800 70712
rect 69200 70728 70000 70848
rect 0 70048 800 70168
rect 0 69640 800 69760
rect 69200 69776 70000 69896
rect 0 69096 800 69216
rect 0 68552 800 68672
rect 69200 68688 70000 68808
rect 0 68144 800 68264
rect 0 67600 800 67720
rect 69200 67736 70000 67856
rect 0 67056 800 67176
rect 0 66648 800 66768
rect 69200 66648 70000 66768
rect 0 66104 800 66224
rect 0 65560 800 65680
rect 69200 65696 70000 65816
rect 0 65152 800 65272
rect 0 64608 800 64728
rect 69200 64608 70000 64728
rect 0 64064 800 64184
rect 0 63656 800 63776
rect 69200 63656 70000 63776
rect 0 63112 800 63232
rect 0 62568 800 62688
rect 69200 62568 70000 62688
rect 0 62160 800 62280
rect 0 61616 800 61736
rect 69200 61616 70000 61736
rect 0 61072 800 61192
rect 0 60528 800 60648
rect 69200 60528 70000 60648
rect 0 60120 800 60240
rect 0 59576 800 59696
rect 69200 59576 70000 59696
rect 0 59032 800 59152
rect 0 58624 800 58744
rect 69200 58488 70000 58608
rect 0 58080 800 58200
rect 0 57536 800 57656
rect 69200 57536 70000 57656
rect 0 57128 800 57248
rect 0 56584 800 56704
rect 69200 56448 70000 56568
rect 0 56040 800 56160
rect 0 55632 800 55752
rect 69200 55496 70000 55616
rect 0 55088 800 55208
rect 0 54544 800 54664
rect 69200 54408 70000 54528
rect 0 54136 800 54256
rect 0 53592 800 53712
rect 69200 53456 70000 53576
rect 0 53048 800 53168
rect 0 52640 800 52760
rect 69200 52368 70000 52488
rect 0 52096 800 52216
rect 0 51552 800 51672
rect 69200 51416 70000 51536
rect 0 51144 800 51264
rect 0 50600 800 50720
rect 69200 50328 70000 50448
rect 0 50056 800 50176
rect 0 49648 800 49768
rect 69200 49376 70000 49496
rect 0 49104 800 49224
rect 0 48560 800 48680
rect 0 48152 800 48272
rect 69200 48288 70000 48408
rect 0 47608 800 47728
rect 69200 47336 70000 47456
rect 0 47064 800 47184
rect 0 46656 800 46776
rect 0 46112 800 46232
rect 69200 46248 70000 46368
rect 0 45568 800 45688
rect 69200 45296 70000 45416
rect 0 45024 800 45144
rect 0 44616 800 44736
rect 0 44072 800 44192
rect 69200 44208 70000 44328
rect 0 43528 800 43648
rect 0 43120 800 43240
rect 69200 43256 70000 43376
rect 0 42576 800 42696
rect 0 42032 800 42152
rect 69200 42168 70000 42288
rect 0 41624 800 41744
rect 0 41080 800 41200
rect 69200 41216 70000 41336
rect 0 40536 800 40656
rect 0 40128 800 40248
rect 69200 40128 70000 40248
rect 0 39584 800 39704
rect 0 39040 800 39160
rect 69200 39176 70000 39296
rect 0 38632 800 38752
rect 0 38088 800 38208
rect 69200 38088 70000 38208
rect 0 37544 800 37664
rect 0 37136 800 37256
rect 69200 37136 70000 37256
rect 0 36592 800 36712
rect 0 36048 800 36168
rect 69200 36048 70000 36168
rect 0 35640 800 35760
rect 0 35096 800 35216
rect 69200 35096 70000 35216
rect 0 34552 800 34672
rect 0 34144 800 34264
rect 69200 34008 70000 34128
rect 0 33600 800 33720
rect 0 33056 800 33176
rect 69200 33056 70000 33176
rect 0 32648 800 32768
rect 0 32104 800 32224
rect 69200 31968 70000 32088
rect 0 31560 800 31680
rect 0 31152 800 31272
rect 69200 31016 70000 31136
rect 0 30608 800 30728
rect 0 30064 800 30184
rect 69200 29928 70000 30048
rect 0 29520 800 29640
rect 0 29112 800 29232
rect 69200 28976 70000 29096
rect 0 28568 800 28688
rect 0 28024 800 28144
rect 69200 27888 70000 28008
rect 0 27616 800 27736
rect 0 27072 800 27192
rect 69200 26936 70000 27056
rect 0 26528 800 26648
rect 0 26120 800 26240
rect 69200 25848 70000 25968
rect 0 25576 800 25696
rect 0 25032 800 25152
rect 69200 24896 70000 25016
rect 0 24624 800 24744
rect 0 24080 800 24200
rect 69200 23808 70000 23928
rect 0 23536 800 23656
rect 0 23128 800 23248
rect 69200 22856 70000 22976
rect 0 22584 800 22704
rect 0 22040 800 22160
rect 0 21632 800 21752
rect 69200 21768 70000 21888
rect 0 21088 800 21208
rect 69200 20816 70000 20936
rect 0 20544 800 20664
rect 0 20136 800 20256
rect 0 19592 800 19712
rect 69200 19728 70000 19848
rect 0 19048 800 19168
rect 0 18640 800 18760
rect 69200 18776 70000 18896
rect 0 18096 800 18216
rect 0 17552 800 17672
rect 69200 17688 70000 17808
rect 0 17144 800 17264
rect 0 16600 800 16720
rect 69200 16736 70000 16856
rect 0 16056 800 16176
rect 0 15648 800 15768
rect 69200 15648 70000 15768
rect 0 15104 800 15224
rect 0 14560 800 14680
rect 69200 14696 70000 14816
rect 0 14016 800 14136
rect 0 13608 800 13728
rect 69200 13608 70000 13728
rect 0 13064 800 13184
rect 0 12520 800 12640
rect 69200 12656 70000 12776
rect 0 12112 800 12232
rect 0 11568 800 11688
rect 69200 11568 70000 11688
rect 0 11024 800 11144
rect 0 10616 800 10736
rect 69200 10616 70000 10736
rect 0 10072 800 10192
rect 0 9528 800 9648
rect 69200 9528 70000 9648
rect 0 9120 800 9240
rect 0 8576 800 8696
rect 69200 8576 70000 8696
rect 0 8032 800 8152
rect 0 7624 800 7744
rect 69200 7488 70000 7608
rect 0 7080 800 7200
rect 0 6536 800 6656
rect 69200 6536 70000 6656
rect 0 6128 800 6248
rect 0 5584 800 5704
rect 69200 5448 70000 5568
rect 0 5040 800 5160
rect 0 4632 800 4752
rect 69200 4496 70000 4616
rect 0 4088 800 4208
rect 0 3544 800 3664
rect 69200 3408 70000 3528
rect 0 3136 800 3256
rect 0 2592 800 2712
rect 69200 2456 70000 2576
rect 0 2048 800 2168
rect 0 1640 800 1760
rect 69200 1368 70000 1488
rect 0 1096 800 1216
rect 0 552 800 672
rect 69200 416 70000 536
rect 0 144 800 264
<< obsm3 >>
rect 880 199584 69200 199749
rect 880 199576 69120 199584
rect 13 199312 69120 199576
rect 880 199304 69120 199312
rect 880 199032 69200 199304
rect 13 198768 69200 199032
rect 880 198496 69200 198768
rect 880 198488 69120 198496
rect 13 198360 69120 198488
rect 880 198216 69120 198360
rect 880 198080 69200 198216
rect 13 197816 69200 198080
rect 880 197544 69200 197816
rect 880 197536 69120 197544
rect 13 197272 69120 197536
rect 880 197264 69120 197272
rect 880 196992 69200 197264
rect 13 196864 69200 196992
rect 880 196584 69200 196864
rect 13 196456 69200 196584
rect 13 196320 69120 196456
rect 880 196176 69120 196320
rect 880 196040 69200 196176
rect 13 195776 69200 196040
rect 880 195504 69200 195776
rect 880 195496 69120 195504
rect 13 195368 69120 195496
rect 880 195224 69120 195368
rect 880 195088 69200 195224
rect 13 194824 69200 195088
rect 880 194544 69200 194824
rect 13 194416 69200 194544
rect 13 194280 69120 194416
rect 880 194136 69120 194280
rect 880 194000 69200 194136
rect 13 193872 69200 194000
rect 880 193592 69200 193872
rect 13 193464 69200 193592
rect 13 193328 69120 193464
rect 880 193184 69120 193328
rect 880 193048 69200 193184
rect 13 192784 69200 193048
rect 880 192504 69200 192784
rect 13 192376 69200 192504
rect 880 192096 69120 192376
rect 13 191832 69200 192096
rect 880 191552 69200 191832
rect 13 191424 69200 191552
rect 13 191288 69120 191424
rect 880 191144 69120 191288
rect 880 191008 69200 191144
rect 13 190880 69200 191008
rect 880 190600 69200 190880
rect 13 190336 69200 190600
rect 880 190056 69120 190336
rect 13 189792 69200 190056
rect 880 189512 69200 189792
rect 13 189384 69200 189512
rect 880 189104 69120 189384
rect 13 188840 69200 189104
rect 880 188560 69200 188840
rect 13 188296 69200 188560
rect 880 188016 69120 188296
rect 13 187888 69200 188016
rect 880 187608 69200 187888
rect 13 187344 69200 187608
rect 880 187064 69120 187344
rect 13 186800 69200 187064
rect 880 186520 69200 186800
rect 13 186392 69200 186520
rect 880 186256 69200 186392
rect 880 186112 69120 186256
rect 13 185976 69120 186112
rect 13 185848 69200 185976
rect 880 185568 69200 185848
rect 13 185304 69200 185568
rect 880 185024 69120 185304
rect 13 184760 69200 185024
rect 880 184480 69200 184760
rect 13 184352 69200 184480
rect 880 184216 69200 184352
rect 880 184072 69120 184216
rect 13 183936 69120 184072
rect 13 183808 69200 183936
rect 880 183528 69200 183808
rect 13 183264 69200 183528
rect 880 182984 69120 183264
rect 13 182856 69200 182984
rect 880 182576 69200 182856
rect 13 182312 69200 182576
rect 880 182176 69200 182312
rect 880 182032 69120 182176
rect 13 181896 69120 182032
rect 13 181768 69200 181896
rect 880 181488 69200 181768
rect 13 181360 69200 181488
rect 880 181224 69200 181360
rect 880 181080 69120 181224
rect 13 180944 69120 181080
rect 13 180816 69200 180944
rect 880 180536 69200 180816
rect 13 180272 69200 180536
rect 880 180136 69200 180272
rect 880 179992 69120 180136
rect 13 179864 69120 179992
rect 880 179856 69120 179864
rect 880 179584 69200 179856
rect 13 179320 69200 179584
rect 880 179184 69200 179320
rect 880 179040 69120 179184
rect 13 178904 69120 179040
rect 13 178776 69200 178904
rect 880 178496 69200 178776
rect 13 178368 69200 178496
rect 880 178096 69200 178368
rect 880 178088 69120 178096
rect 13 177824 69120 178088
rect 880 177816 69120 177824
rect 880 177544 69200 177816
rect 13 177280 69200 177544
rect 880 177144 69200 177280
rect 880 177000 69120 177144
rect 13 176872 69120 177000
rect 880 176864 69120 176872
rect 880 176592 69200 176864
rect 13 176328 69200 176592
rect 880 176056 69200 176328
rect 880 176048 69120 176056
rect 13 175784 69120 176048
rect 880 175776 69120 175784
rect 880 175504 69200 175776
rect 13 175376 69200 175504
rect 880 175104 69200 175376
rect 880 175096 69120 175104
rect 13 174832 69120 175096
rect 880 174824 69120 174832
rect 880 174552 69200 174824
rect 13 174288 69200 174552
rect 880 174016 69200 174288
rect 880 174008 69120 174016
rect 13 173880 69120 174008
rect 880 173736 69120 173880
rect 880 173600 69200 173736
rect 13 173336 69200 173600
rect 880 173064 69200 173336
rect 880 173056 69120 173064
rect 13 172792 69120 173056
rect 880 172784 69120 172792
rect 880 172512 69200 172784
rect 13 172384 69200 172512
rect 880 172104 69200 172384
rect 13 171976 69200 172104
rect 13 171840 69120 171976
rect 880 171696 69120 171840
rect 880 171560 69200 171696
rect 13 171296 69200 171560
rect 880 171024 69200 171296
rect 880 171016 69120 171024
rect 13 170888 69120 171016
rect 880 170744 69120 170888
rect 880 170608 69200 170744
rect 13 170344 69200 170608
rect 880 170064 69200 170344
rect 13 169936 69200 170064
rect 13 169800 69120 169936
rect 880 169656 69120 169800
rect 880 169520 69200 169656
rect 13 169256 69200 169520
rect 880 168984 69200 169256
rect 880 168976 69120 168984
rect 13 168848 69120 168976
rect 880 168704 69120 168848
rect 880 168568 69200 168704
rect 13 168304 69200 168568
rect 880 168024 69200 168304
rect 13 167896 69200 168024
rect 13 167760 69120 167896
rect 880 167616 69120 167760
rect 880 167480 69200 167616
rect 13 167352 69200 167480
rect 880 167072 69200 167352
rect 13 166944 69200 167072
rect 13 166808 69120 166944
rect 880 166664 69120 166808
rect 880 166528 69200 166664
rect 13 166264 69200 166528
rect 880 165984 69200 166264
rect 13 165856 69200 165984
rect 880 165576 69120 165856
rect 13 165312 69200 165576
rect 880 165032 69200 165312
rect 13 164904 69200 165032
rect 13 164768 69120 164904
rect 880 164624 69120 164768
rect 880 164488 69200 164624
rect 13 164360 69200 164488
rect 880 164080 69200 164360
rect 13 163816 69200 164080
rect 880 163536 69120 163816
rect 13 163272 69200 163536
rect 880 162992 69200 163272
rect 13 162864 69200 162992
rect 880 162584 69120 162864
rect 13 162320 69200 162584
rect 880 162040 69200 162320
rect 13 161776 69200 162040
rect 880 161496 69120 161776
rect 13 161368 69200 161496
rect 880 161088 69200 161368
rect 13 160824 69200 161088
rect 880 160544 69120 160824
rect 13 160280 69200 160544
rect 880 160000 69200 160280
rect 13 159872 69200 160000
rect 880 159736 69200 159872
rect 880 159592 69120 159736
rect 13 159456 69120 159592
rect 13 159328 69200 159456
rect 880 159048 69200 159328
rect 13 158784 69200 159048
rect 880 158504 69120 158784
rect 13 158376 69200 158504
rect 880 158096 69200 158376
rect 13 157832 69200 158096
rect 880 157696 69200 157832
rect 880 157552 69120 157696
rect 13 157416 69120 157552
rect 13 157288 69200 157416
rect 880 157008 69200 157288
rect 13 156880 69200 157008
rect 880 156744 69200 156880
rect 880 156600 69120 156744
rect 13 156464 69120 156600
rect 13 156336 69200 156464
rect 880 156056 69200 156336
rect 13 155792 69200 156056
rect 880 155656 69200 155792
rect 880 155512 69120 155656
rect 13 155384 69120 155512
rect 880 155376 69120 155384
rect 880 155104 69200 155376
rect 13 154840 69200 155104
rect 880 154704 69200 154840
rect 880 154560 69120 154704
rect 13 154424 69120 154560
rect 13 154296 69200 154424
rect 880 154016 69200 154296
rect 13 153752 69200 154016
rect 880 153616 69200 153752
rect 880 153472 69120 153616
rect 13 153344 69120 153472
rect 880 153336 69120 153344
rect 880 153064 69200 153336
rect 13 152800 69200 153064
rect 880 152664 69200 152800
rect 880 152520 69120 152664
rect 13 152384 69120 152520
rect 13 152256 69200 152384
rect 880 151976 69200 152256
rect 13 151848 69200 151976
rect 880 151576 69200 151848
rect 880 151568 69120 151576
rect 13 151304 69120 151568
rect 880 151296 69120 151304
rect 880 151024 69200 151296
rect 13 150760 69200 151024
rect 880 150624 69200 150760
rect 880 150480 69120 150624
rect 13 150352 69120 150480
rect 880 150344 69120 150352
rect 880 150072 69200 150344
rect 13 149808 69200 150072
rect 880 149536 69200 149808
rect 880 149528 69120 149536
rect 13 149264 69120 149528
rect 880 149256 69120 149264
rect 880 148984 69200 149256
rect 13 148856 69200 148984
rect 880 148584 69200 148856
rect 880 148576 69120 148584
rect 13 148312 69120 148576
rect 880 148304 69120 148312
rect 880 148032 69200 148304
rect 13 147768 69200 148032
rect 880 147496 69200 147768
rect 880 147488 69120 147496
rect 13 147360 69120 147488
rect 880 147216 69120 147360
rect 880 147080 69200 147216
rect 13 146816 69200 147080
rect 880 146544 69200 146816
rect 880 146536 69120 146544
rect 13 146272 69120 146536
rect 880 146264 69120 146272
rect 880 145992 69200 146264
rect 13 145864 69200 145992
rect 880 145584 69200 145864
rect 13 145456 69200 145584
rect 13 145320 69120 145456
rect 880 145176 69120 145320
rect 880 145040 69200 145176
rect 13 144776 69200 145040
rect 880 144504 69200 144776
rect 880 144496 69120 144504
rect 13 144368 69120 144496
rect 880 144224 69120 144368
rect 880 144088 69200 144224
rect 13 143824 69200 144088
rect 880 143544 69200 143824
rect 13 143416 69200 143544
rect 13 143280 69120 143416
rect 880 143136 69120 143280
rect 880 143000 69200 143136
rect 13 142872 69200 143000
rect 880 142592 69200 142872
rect 13 142464 69200 142592
rect 13 142328 69120 142464
rect 880 142184 69120 142328
rect 880 142048 69200 142184
rect 13 141784 69200 142048
rect 880 141504 69200 141784
rect 13 141376 69200 141504
rect 880 141096 69120 141376
rect 13 140832 69200 141096
rect 880 140552 69200 140832
rect 13 140424 69200 140552
rect 13 140288 69120 140424
rect 880 140144 69120 140288
rect 880 140008 69200 140144
rect 13 139880 69200 140008
rect 880 139600 69200 139880
rect 13 139336 69200 139600
rect 880 139056 69120 139336
rect 13 138792 69200 139056
rect 880 138512 69200 138792
rect 13 138384 69200 138512
rect 13 138248 69120 138384
rect 880 138104 69120 138248
rect 880 137968 69200 138104
rect 13 137840 69200 137968
rect 880 137560 69200 137840
rect 13 137296 69200 137560
rect 880 137016 69120 137296
rect 13 136752 69200 137016
rect 880 136472 69200 136752
rect 13 136344 69200 136472
rect 880 136064 69120 136344
rect 13 135800 69200 136064
rect 880 135520 69200 135800
rect 13 135256 69200 135520
rect 880 134976 69120 135256
rect 13 134848 69200 134976
rect 880 134568 69200 134848
rect 13 134304 69200 134568
rect 880 134024 69120 134304
rect 13 133760 69200 134024
rect 880 133480 69200 133760
rect 13 133352 69200 133480
rect 880 133216 69200 133352
rect 880 133072 69120 133216
rect 13 132936 69120 133072
rect 13 132808 69200 132936
rect 880 132528 69200 132808
rect 13 132264 69200 132528
rect 880 131984 69120 132264
rect 13 131856 69200 131984
rect 880 131576 69200 131856
rect 13 131312 69200 131576
rect 880 131176 69200 131312
rect 880 131032 69120 131176
rect 13 130896 69120 131032
rect 13 130768 69200 130896
rect 880 130488 69200 130768
rect 13 130360 69200 130488
rect 880 130224 69200 130360
rect 880 130080 69120 130224
rect 13 129944 69120 130080
rect 13 129816 69200 129944
rect 880 129536 69200 129816
rect 13 129272 69200 129536
rect 880 129136 69200 129272
rect 880 128992 69120 129136
rect 13 128864 69120 128992
rect 880 128856 69120 128864
rect 880 128584 69200 128856
rect 13 128320 69200 128584
rect 880 128184 69200 128320
rect 880 128040 69120 128184
rect 13 127904 69120 128040
rect 13 127776 69200 127904
rect 880 127496 69200 127776
rect 13 127368 69200 127496
rect 880 127096 69200 127368
rect 880 127088 69120 127096
rect 13 126824 69120 127088
rect 880 126816 69120 126824
rect 880 126544 69200 126816
rect 13 126280 69200 126544
rect 880 126144 69200 126280
rect 880 126000 69120 126144
rect 13 125872 69120 126000
rect 880 125864 69120 125872
rect 880 125592 69200 125864
rect 13 125328 69200 125592
rect 880 125056 69200 125328
rect 880 125048 69120 125056
rect 13 124784 69120 125048
rect 880 124776 69120 124784
rect 880 124504 69200 124776
rect 13 124376 69200 124504
rect 880 124104 69200 124376
rect 880 124096 69120 124104
rect 13 123832 69120 124096
rect 880 123824 69120 123832
rect 880 123552 69200 123824
rect 13 123288 69200 123552
rect 880 123016 69200 123288
rect 880 123008 69120 123016
rect 13 122744 69120 123008
rect 880 122736 69120 122744
rect 880 122464 69200 122736
rect 13 122336 69200 122464
rect 880 122064 69200 122336
rect 880 122056 69120 122064
rect 13 121792 69120 122056
rect 880 121784 69120 121792
rect 880 121512 69200 121784
rect 13 121248 69200 121512
rect 880 120976 69200 121248
rect 880 120968 69120 120976
rect 13 120840 69120 120968
rect 880 120696 69120 120840
rect 880 120560 69200 120696
rect 13 120296 69200 120560
rect 880 120024 69200 120296
rect 880 120016 69120 120024
rect 13 119752 69120 120016
rect 880 119744 69120 119752
rect 880 119472 69200 119744
rect 13 119344 69200 119472
rect 880 119064 69200 119344
rect 13 118936 69200 119064
rect 13 118800 69120 118936
rect 880 118656 69120 118800
rect 880 118520 69200 118656
rect 13 118256 69200 118520
rect 880 117984 69200 118256
rect 880 117976 69120 117984
rect 13 117848 69120 117976
rect 880 117704 69120 117848
rect 880 117568 69200 117704
rect 13 117304 69200 117568
rect 880 117024 69200 117304
rect 13 116896 69200 117024
rect 13 116760 69120 116896
rect 880 116616 69120 116760
rect 880 116480 69200 116616
rect 13 116352 69200 116480
rect 880 116072 69200 116352
rect 13 115944 69200 116072
rect 13 115808 69120 115944
rect 880 115664 69120 115808
rect 880 115528 69200 115664
rect 13 115264 69200 115528
rect 880 114984 69200 115264
rect 13 114856 69200 114984
rect 880 114576 69120 114856
rect 13 114312 69200 114576
rect 880 114032 69200 114312
rect 13 113904 69200 114032
rect 13 113768 69120 113904
rect 880 113624 69120 113768
rect 880 113488 69200 113624
rect 13 113360 69200 113488
rect 880 113080 69200 113360
rect 13 112816 69200 113080
rect 880 112536 69120 112816
rect 13 112272 69200 112536
rect 880 111992 69200 112272
rect 13 111864 69200 111992
rect 880 111584 69120 111864
rect 13 111320 69200 111584
rect 880 111040 69200 111320
rect 13 110776 69200 111040
rect 880 110496 69120 110776
rect 13 110368 69200 110496
rect 880 110088 69200 110368
rect 13 109824 69200 110088
rect 880 109544 69120 109824
rect 13 109280 69200 109544
rect 880 109000 69200 109280
rect 13 108872 69200 109000
rect 880 108736 69200 108872
rect 880 108592 69120 108736
rect 13 108456 69120 108592
rect 13 108328 69200 108456
rect 880 108048 69200 108328
rect 13 107784 69200 108048
rect 880 107504 69120 107784
rect 13 107240 69200 107504
rect 880 106960 69200 107240
rect 13 106832 69200 106960
rect 880 106696 69200 106832
rect 880 106552 69120 106696
rect 13 106416 69120 106552
rect 13 106288 69200 106416
rect 880 106008 69200 106288
rect 13 105744 69200 106008
rect 880 105464 69120 105744
rect 13 105336 69200 105464
rect 880 105056 69200 105336
rect 13 104792 69200 105056
rect 880 104656 69200 104792
rect 880 104512 69120 104656
rect 13 104376 69120 104512
rect 13 104248 69200 104376
rect 880 103968 69200 104248
rect 13 103840 69200 103968
rect 880 103704 69200 103840
rect 880 103560 69120 103704
rect 13 103424 69120 103560
rect 13 103296 69200 103424
rect 880 103016 69200 103296
rect 13 102752 69200 103016
rect 880 102616 69200 102752
rect 880 102472 69120 102616
rect 13 102344 69120 102472
rect 880 102336 69120 102344
rect 880 102064 69200 102336
rect 13 101800 69200 102064
rect 880 101664 69200 101800
rect 880 101520 69120 101664
rect 13 101384 69120 101520
rect 13 101256 69200 101384
rect 880 100976 69200 101256
rect 13 100848 69200 100976
rect 880 100576 69200 100848
rect 880 100568 69120 100576
rect 13 100304 69120 100568
rect 880 100296 69120 100304
rect 880 100024 69200 100296
rect 13 99760 69200 100024
rect 880 99488 69200 99760
rect 880 99480 69120 99488
rect 13 99352 69120 99480
rect 880 99208 69120 99352
rect 880 99072 69200 99208
rect 13 98808 69200 99072
rect 880 98536 69200 98808
rect 880 98528 69120 98536
rect 13 98264 69120 98528
rect 880 98256 69120 98264
rect 880 97984 69200 98256
rect 13 97856 69200 97984
rect 880 97576 69200 97856
rect 13 97448 69200 97576
rect 13 97312 69120 97448
rect 880 97168 69120 97312
rect 880 97032 69200 97168
rect 13 96768 69200 97032
rect 880 96496 69200 96768
rect 880 96488 69120 96496
rect 13 96360 69120 96488
rect 880 96216 69120 96360
rect 880 96080 69200 96216
rect 13 95816 69200 96080
rect 880 95536 69200 95816
rect 13 95408 69200 95536
rect 13 95272 69120 95408
rect 880 95128 69120 95272
rect 880 94992 69200 95128
rect 13 94864 69200 94992
rect 880 94584 69200 94864
rect 13 94456 69200 94584
rect 13 94320 69120 94456
rect 880 94176 69120 94320
rect 880 94040 69200 94176
rect 13 93776 69200 94040
rect 880 93496 69200 93776
rect 13 93368 69200 93496
rect 880 93088 69120 93368
rect 13 92824 69200 93088
rect 880 92544 69200 92824
rect 13 92416 69200 92544
rect 13 92280 69120 92416
rect 880 92136 69120 92280
rect 880 92000 69200 92136
rect 13 91736 69200 92000
rect 880 91456 69200 91736
rect 13 91328 69200 91456
rect 880 91048 69120 91328
rect 13 90784 69200 91048
rect 880 90504 69200 90784
rect 13 90376 69200 90504
rect 13 90240 69120 90376
rect 880 90096 69120 90240
rect 880 89960 69200 90096
rect 13 89832 69200 89960
rect 880 89552 69200 89832
rect 13 89288 69200 89552
rect 880 89008 69120 89288
rect 13 88744 69200 89008
rect 880 88464 69200 88744
rect 13 88336 69200 88464
rect 880 88056 69120 88336
rect 13 87792 69200 88056
rect 880 87512 69200 87792
rect 13 87248 69200 87512
rect 880 86968 69120 87248
rect 13 86840 69200 86968
rect 880 86560 69200 86840
rect 13 86296 69200 86560
rect 880 86016 69120 86296
rect 13 85752 69200 86016
rect 880 85472 69200 85752
rect 13 85344 69200 85472
rect 880 85208 69200 85344
rect 880 85064 69120 85208
rect 13 84928 69120 85064
rect 13 84800 69200 84928
rect 880 84520 69200 84800
rect 13 84256 69200 84520
rect 880 83976 69120 84256
rect 13 83848 69200 83976
rect 880 83568 69200 83848
rect 13 83304 69200 83568
rect 880 83168 69200 83304
rect 880 83024 69120 83168
rect 13 82888 69120 83024
rect 13 82760 69200 82888
rect 880 82480 69200 82760
rect 13 82352 69200 82480
rect 880 82216 69200 82352
rect 880 82072 69120 82216
rect 13 81936 69120 82072
rect 13 81808 69200 81936
rect 880 81528 69200 81808
rect 13 81264 69200 81528
rect 880 81128 69200 81264
rect 880 80984 69120 81128
rect 13 80856 69120 80984
rect 880 80848 69120 80856
rect 880 80576 69200 80848
rect 13 80312 69200 80576
rect 880 80176 69200 80312
rect 880 80032 69120 80176
rect 13 79896 69120 80032
rect 13 79768 69200 79896
rect 880 79488 69200 79768
rect 13 79360 69200 79488
rect 880 79088 69200 79360
rect 880 79080 69120 79088
rect 13 78816 69120 79080
rect 880 78808 69120 78816
rect 880 78536 69200 78808
rect 13 78272 69200 78536
rect 880 78136 69200 78272
rect 880 77992 69120 78136
rect 13 77864 69120 77992
rect 880 77856 69120 77864
rect 880 77584 69200 77856
rect 13 77320 69200 77584
rect 880 77048 69200 77320
rect 880 77040 69120 77048
rect 13 76776 69120 77040
rect 880 76768 69120 76776
rect 880 76496 69200 76768
rect 13 76232 69200 76496
rect 880 76096 69200 76232
rect 880 75952 69120 76096
rect 13 75824 69120 75952
rect 880 75816 69120 75824
rect 880 75544 69200 75816
rect 13 75280 69200 75544
rect 880 75008 69200 75280
rect 880 75000 69120 75008
rect 13 74736 69120 75000
rect 880 74728 69120 74736
rect 880 74456 69200 74728
rect 13 74328 69200 74456
rect 880 74056 69200 74328
rect 880 74048 69120 74056
rect 13 73784 69120 74048
rect 880 73776 69120 73784
rect 880 73504 69200 73776
rect 13 73240 69200 73504
rect 880 72968 69200 73240
rect 880 72960 69120 72968
rect 13 72832 69120 72960
rect 880 72688 69120 72832
rect 880 72552 69200 72688
rect 13 72288 69200 72552
rect 880 72016 69200 72288
rect 880 72008 69120 72016
rect 13 71744 69120 72008
rect 880 71736 69120 71744
rect 880 71464 69200 71736
rect 13 71336 69200 71464
rect 880 71056 69200 71336
rect 13 70928 69200 71056
rect 13 70792 69120 70928
rect 880 70648 69120 70792
rect 880 70512 69200 70648
rect 13 70248 69200 70512
rect 880 69976 69200 70248
rect 880 69968 69120 69976
rect 13 69840 69120 69968
rect 880 69696 69120 69840
rect 880 69560 69200 69696
rect 13 69296 69200 69560
rect 880 69016 69200 69296
rect 13 68888 69200 69016
rect 13 68752 69120 68888
rect 880 68608 69120 68752
rect 880 68472 69200 68608
rect 13 68344 69200 68472
rect 880 68064 69200 68344
rect 13 67936 69200 68064
rect 13 67800 69120 67936
rect 880 67656 69120 67800
rect 880 67520 69200 67656
rect 13 67256 69200 67520
rect 880 66976 69200 67256
rect 13 66848 69200 66976
rect 880 66568 69120 66848
rect 13 66304 69200 66568
rect 880 66024 69200 66304
rect 13 65896 69200 66024
rect 13 65760 69120 65896
rect 880 65616 69120 65760
rect 880 65480 69200 65616
rect 13 65352 69200 65480
rect 880 65072 69200 65352
rect 13 64808 69200 65072
rect 880 64528 69120 64808
rect 13 64264 69200 64528
rect 880 63984 69200 64264
rect 13 63856 69200 63984
rect 880 63576 69120 63856
rect 13 63312 69200 63576
rect 880 63032 69200 63312
rect 13 62768 69200 63032
rect 880 62488 69120 62768
rect 13 62360 69200 62488
rect 880 62080 69200 62360
rect 13 61816 69200 62080
rect 880 61536 69120 61816
rect 13 61272 69200 61536
rect 880 60992 69200 61272
rect 13 60728 69200 60992
rect 880 60448 69120 60728
rect 13 60320 69200 60448
rect 880 60040 69200 60320
rect 13 59776 69200 60040
rect 880 59496 69120 59776
rect 13 59232 69200 59496
rect 880 58952 69200 59232
rect 13 58824 69200 58952
rect 880 58688 69200 58824
rect 880 58544 69120 58688
rect 13 58408 69120 58544
rect 13 58280 69200 58408
rect 880 58000 69200 58280
rect 13 57736 69200 58000
rect 880 57456 69120 57736
rect 13 57328 69200 57456
rect 880 57048 69200 57328
rect 13 56784 69200 57048
rect 880 56648 69200 56784
rect 880 56504 69120 56648
rect 13 56368 69120 56504
rect 13 56240 69200 56368
rect 880 55960 69200 56240
rect 13 55832 69200 55960
rect 880 55696 69200 55832
rect 880 55552 69120 55696
rect 13 55416 69120 55552
rect 13 55288 69200 55416
rect 880 55008 69200 55288
rect 13 54744 69200 55008
rect 880 54608 69200 54744
rect 880 54464 69120 54608
rect 13 54336 69120 54464
rect 880 54328 69120 54336
rect 880 54056 69200 54328
rect 13 53792 69200 54056
rect 880 53656 69200 53792
rect 880 53512 69120 53656
rect 13 53376 69120 53512
rect 13 53248 69200 53376
rect 880 52968 69200 53248
rect 13 52840 69200 52968
rect 880 52568 69200 52840
rect 880 52560 69120 52568
rect 13 52296 69120 52560
rect 880 52288 69120 52296
rect 880 52016 69200 52288
rect 13 51752 69200 52016
rect 880 51616 69200 51752
rect 880 51472 69120 51616
rect 13 51344 69120 51472
rect 880 51336 69120 51344
rect 880 51064 69200 51336
rect 13 50800 69200 51064
rect 880 50528 69200 50800
rect 880 50520 69120 50528
rect 13 50256 69120 50520
rect 880 50248 69120 50256
rect 880 49976 69200 50248
rect 13 49848 69200 49976
rect 880 49576 69200 49848
rect 880 49568 69120 49576
rect 13 49304 69120 49568
rect 880 49296 69120 49304
rect 880 49024 69200 49296
rect 13 48760 69200 49024
rect 880 48488 69200 48760
rect 880 48480 69120 48488
rect 13 48352 69120 48480
rect 880 48208 69120 48352
rect 880 48072 69200 48208
rect 13 47808 69200 48072
rect 880 47536 69200 47808
rect 880 47528 69120 47536
rect 13 47264 69120 47528
rect 880 47256 69120 47264
rect 880 46984 69200 47256
rect 13 46856 69200 46984
rect 880 46576 69200 46856
rect 13 46448 69200 46576
rect 13 46312 69120 46448
rect 880 46168 69120 46312
rect 880 46032 69200 46168
rect 13 45768 69200 46032
rect 880 45496 69200 45768
rect 880 45488 69120 45496
rect 13 45224 69120 45488
rect 880 45216 69120 45224
rect 880 44944 69200 45216
rect 13 44816 69200 44944
rect 880 44536 69200 44816
rect 13 44408 69200 44536
rect 13 44272 69120 44408
rect 880 44128 69120 44272
rect 880 43992 69200 44128
rect 13 43728 69200 43992
rect 880 43456 69200 43728
rect 880 43448 69120 43456
rect 13 43320 69120 43448
rect 880 43176 69120 43320
rect 880 43040 69200 43176
rect 13 42776 69200 43040
rect 880 42496 69200 42776
rect 13 42368 69200 42496
rect 13 42232 69120 42368
rect 880 42088 69120 42232
rect 880 41952 69200 42088
rect 13 41824 69200 41952
rect 880 41544 69200 41824
rect 13 41416 69200 41544
rect 13 41280 69120 41416
rect 880 41136 69120 41280
rect 880 41000 69200 41136
rect 13 40736 69200 41000
rect 880 40456 69200 40736
rect 13 40328 69200 40456
rect 880 40048 69120 40328
rect 13 39784 69200 40048
rect 880 39504 69200 39784
rect 13 39376 69200 39504
rect 13 39240 69120 39376
rect 880 39096 69120 39240
rect 880 38960 69200 39096
rect 13 38832 69200 38960
rect 880 38552 69200 38832
rect 13 38288 69200 38552
rect 880 38008 69120 38288
rect 13 37744 69200 38008
rect 880 37464 69200 37744
rect 13 37336 69200 37464
rect 880 37056 69120 37336
rect 13 36792 69200 37056
rect 880 36512 69200 36792
rect 13 36248 69200 36512
rect 880 35968 69120 36248
rect 13 35840 69200 35968
rect 880 35560 69200 35840
rect 13 35296 69200 35560
rect 880 35016 69120 35296
rect 13 34752 69200 35016
rect 880 34472 69200 34752
rect 13 34344 69200 34472
rect 880 34208 69200 34344
rect 880 34064 69120 34208
rect 13 33928 69120 34064
rect 13 33800 69200 33928
rect 880 33520 69200 33800
rect 13 33256 69200 33520
rect 880 32976 69120 33256
rect 13 32848 69200 32976
rect 880 32568 69200 32848
rect 13 32304 69200 32568
rect 880 32168 69200 32304
rect 880 32024 69120 32168
rect 13 31888 69120 32024
rect 13 31760 69200 31888
rect 880 31480 69200 31760
rect 13 31352 69200 31480
rect 880 31216 69200 31352
rect 880 31072 69120 31216
rect 13 30936 69120 31072
rect 13 30808 69200 30936
rect 880 30528 69200 30808
rect 13 30264 69200 30528
rect 880 30128 69200 30264
rect 880 29984 69120 30128
rect 13 29848 69120 29984
rect 13 29720 69200 29848
rect 880 29440 69200 29720
rect 13 29312 69200 29440
rect 880 29176 69200 29312
rect 880 29032 69120 29176
rect 13 28896 69120 29032
rect 13 28768 69200 28896
rect 880 28488 69200 28768
rect 13 28224 69200 28488
rect 880 28088 69200 28224
rect 880 27944 69120 28088
rect 13 27816 69120 27944
rect 880 27808 69120 27816
rect 880 27536 69200 27808
rect 13 27272 69200 27536
rect 880 27136 69200 27272
rect 880 26992 69120 27136
rect 13 26856 69120 26992
rect 13 26728 69200 26856
rect 880 26448 69200 26728
rect 13 26320 69200 26448
rect 880 26048 69200 26320
rect 880 26040 69120 26048
rect 13 25776 69120 26040
rect 880 25768 69120 25776
rect 880 25496 69200 25768
rect 13 25232 69200 25496
rect 880 25096 69200 25232
rect 880 24952 69120 25096
rect 13 24824 69120 24952
rect 880 24816 69120 24824
rect 880 24544 69200 24816
rect 13 24280 69200 24544
rect 880 24008 69200 24280
rect 880 24000 69120 24008
rect 13 23736 69120 24000
rect 880 23728 69120 23736
rect 880 23456 69200 23728
rect 13 23328 69200 23456
rect 880 23056 69200 23328
rect 880 23048 69120 23056
rect 13 22784 69120 23048
rect 880 22776 69120 22784
rect 880 22504 69200 22776
rect 13 22240 69200 22504
rect 880 21968 69200 22240
rect 880 21960 69120 21968
rect 13 21832 69120 21960
rect 880 21688 69120 21832
rect 880 21552 69200 21688
rect 13 21288 69200 21552
rect 880 21016 69200 21288
rect 880 21008 69120 21016
rect 13 20744 69120 21008
rect 880 20736 69120 20744
rect 880 20464 69200 20736
rect 13 20336 69200 20464
rect 880 20056 69200 20336
rect 13 19928 69200 20056
rect 13 19792 69120 19928
rect 880 19648 69120 19792
rect 880 19512 69200 19648
rect 13 19248 69200 19512
rect 880 18976 69200 19248
rect 880 18968 69120 18976
rect 13 18840 69120 18968
rect 880 18696 69120 18840
rect 880 18560 69200 18696
rect 13 18296 69200 18560
rect 880 18016 69200 18296
rect 13 17888 69200 18016
rect 13 17752 69120 17888
rect 880 17608 69120 17752
rect 880 17472 69200 17608
rect 13 17344 69200 17472
rect 880 17064 69200 17344
rect 13 16936 69200 17064
rect 13 16800 69120 16936
rect 880 16656 69120 16800
rect 880 16520 69200 16656
rect 13 16256 69200 16520
rect 880 15976 69200 16256
rect 13 15848 69200 15976
rect 880 15568 69120 15848
rect 13 15304 69200 15568
rect 880 15024 69200 15304
rect 13 14896 69200 15024
rect 13 14760 69120 14896
rect 880 14616 69120 14760
rect 880 14480 69200 14616
rect 13 14216 69200 14480
rect 880 13936 69200 14216
rect 13 13808 69200 13936
rect 880 13528 69120 13808
rect 13 13264 69200 13528
rect 880 12984 69200 13264
rect 13 12856 69200 12984
rect 13 12720 69120 12856
rect 880 12576 69120 12720
rect 880 12440 69200 12576
rect 13 12312 69200 12440
rect 880 12032 69200 12312
rect 13 11768 69200 12032
rect 880 11488 69120 11768
rect 13 11224 69200 11488
rect 880 10944 69200 11224
rect 13 10816 69200 10944
rect 880 10536 69120 10816
rect 13 10272 69200 10536
rect 880 9992 69200 10272
rect 13 9728 69200 9992
rect 880 9448 69120 9728
rect 13 9320 69200 9448
rect 880 9040 69200 9320
rect 13 8776 69200 9040
rect 880 8496 69120 8776
rect 13 8232 69200 8496
rect 880 7952 69200 8232
rect 13 7824 69200 7952
rect 880 7688 69200 7824
rect 880 7544 69120 7688
rect 13 7408 69120 7544
rect 13 7280 69200 7408
rect 880 7000 69200 7280
rect 13 6736 69200 7000
rect 880 6456 69120 6736
rect 13 6328 69200 6456
rect 880 6048 69200 6328
rect 13 5784 69200 6048
rect 880 5648 69200 5784
rect 880 5504 69120 5648
rect 13 5368 69120 5504
rect 13 5240 69200 5368
rect 880 4960 69200 5240
rect 13 4832 69200 4960
rect 880 4696 69200 4832
rect 880 4552 69120 4696
rect 13 4416 69120 4552
rect 13 4288 69200 4416
rect 880 4008 69200 4288
rect 13 3744 69200 4008
rect 880 3608 69200 3744
rect 880 3464 69120 3608
rect 13 3336 69120 3464
rect 880 3328 69120 3336
rect 880 3056 69200 3328
rect 13 2792 69200 3056
rect 880 2656 69200 2792
rect 880 2512 69120 2656
rect 13 2376 69120 2512
rect 13 2248 69200 2376
rect 880 1968 69200 2248
rect 13 1840 69200 1968
rect 880 1568 69200 1840
rect 880 1560 69120 1568
rect 13 1296 69120 1560
rect 880 1288 69120 1296
rect 880 1016 69200 1288
rect 13 752 69200 1016
rect 880 616 69200 752
rect 880 472 69120 616
rect 13 344 69120 472
rect 880 336 69120 344
rect 880 171 69200 336
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
<< obsm4 >>
rect 427 2619 4128 197165
rect 4608 2619 19488 197165
rect 19968 2619 34848 197165
rect 35328 2619 47229 197165
<< labels >>
rlabel metal2 s 13542 0 13598 800 6 master0_wb_ack_i
port 1 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 master0_wb_adr_o[0]
port 2 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 master0_wb_adr_o[10]
port 3 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 master0_wb_adr_o[11]
port 4 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 master0_wb_adr_o[12]
port 5 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 master0_wb_adr_o[13]
port 6 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 master0_wb_adr_o[14]
port 7 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 master0_wb_adr_o[15]
port 8 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 master0_wb_adr_o[16]
port 9 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 master0_wb_adr_o[17]
port 10 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 master0_wb_adr_o[18]
port 11 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 master0_wb_adr_o[19]
port 12 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 master0_wb_adr_o[1]
port 13 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 master0_wb_adr_o[20]
port 14 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 master0_wb_adr_o[21]
port 15 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 master0_wb_adr_o[22]
port 16 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 master0_wb_adr_o[23]
port 17 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 master0_wb_adr_o[24]
port 18 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 master0_wb_adr_o[25]
port 19 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 master0_wb_adr_o[26]
port 20 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 master0_wb_adr_o[27]
port 21 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 master0_wb_adr_o[2]
port 22 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 master0_wb_adr_o[3]
port 23 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 master0_wb_adr_o[4]
port 24 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 master0_wb_adr_o[5]
port 25 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 master0_wb_adr_o[6]
port 26 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 master0_wb_adr_o[7]
port 27 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 master0_wb_adr_o[8]
port 28 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 master0_wb_adr_o[9]
port 29 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 master0_wb_cyc_o
port 30 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 master0_wb_data_i[0]
port 31 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 master0_wb_data_i[10]
port 32 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 master0_wb_data_i[11]
port 33 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 master0_wb_data_i[12]
port 34 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 master0_wb_data_i[13]
port 35 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 master0_wb_data_i[14]
port 36 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 master0_wb_data_i[15]
port 37 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 master0_wb_data_i[16]
port 38 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 master0_wb_data_i[17]
port 39 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 master0_wb_data_i[18]
port 40 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 master0_wb_data_i[19]
port 41 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 master0_wb_data_i[1]
port 42 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 master0_wb_data_i[20]
port 43 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 master0_wb_data_i[21]
port 44 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 master0_wb_data_i[22]
port 45 nsew signal output
rlabel metal2 s 58070 0 58126 800 6 master0_wb_data_i[23]
port 46 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 master0_wb_data_i[24]
port 47 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 master0_wb_data_i[25]
port 48 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 master0_wb_data_i[26]
port 49 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 master0_wb_data_i[27]
port 50 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 master0_wb_data_i[28]
port 51 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 master0_wb_data_i[29]
port 52 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 master0_wb_data_i[2]
port 53 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 master0_wb_data_i[30]
port 54 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 master0_wb_data_i[31]
port 55 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 master0_wb_data_i[3]
port 56 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 master0_wb_data_i[4]
port 57 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 master0_wb_data_i[5]
port 58 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 master0_wb_data_i[6]
port 59 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 master0_wb_data_i[7]
port 60 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 master0_wb_data_i[8]
port 61 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 master0_wb_data_i[9]
port 62 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 master0_wb_data_o[0]
port 63 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 master0_wb_data_o[10]
port 64 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 master0_wb_data_o[11]
port 65 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 master0_wb_data_o[12]
port 66 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 master0_wb_data_o[13]
port 67 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 master0_wb_data_o[14]
port 68 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 master0_wb_data_o[15]
port 69 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 master0_wb_data_o[16]
port 70 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 master0_wb_data_o[17]
port 71 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 master0_wb_data_o[18]
port 72 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 master0_wb_data_o[19]
port 73 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 master0_wb_data_o[1]
port 74 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 master0_wb_data_o[20]
port 75 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 master0_wb_data_o[21]
port 76 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 master0_wb_data_o[22]
port 77 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 master0_wb_data_o[23]
port 78 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 master0_wb_data_o[24]
port 79 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 master0_wb_data_o[25]
port 80 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 master0_wb_data_o[26]
port 81 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 master0_wb_data_o[27]
port 82 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 master0_wb_data_o[28]
port 83 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 master0_wb_data_o[29]
port 84 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 master0_wb_data_o[2]
port 85 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 master0_wb_data_o[30]
port 86 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 master0_wb_data_o[31]
port 87 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 master0_wb_data_o[3]
port 88 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 master0_wb_data_o[4]
port 89 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 master0_wb_data_o[5]
port 90 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 master0_wb_data_o[6]
port 91 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 master0_wb_data_o[7]
port 92 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 master0_wb_data_o[8]
port 93 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 master0_wb_data_o[9]
port 94 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 master0_wb_error_i
port 95 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 master0_wb_sel_o[0]
port 96 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 master0_wb_sel_o[1]
port 97 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 master0_wb_sel_o[2]
port 98 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 master0_wb_sel_o[3]
port 99 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 master0_wb_stall_i
port 100 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 master0_wb_stb_o
port 101 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 master0_wb_we_o
port 102 nsew signal input
rlabel metal3 s 0 100104 800 100224 6 master1_wb_ack_i
port 103 nsew signal output
rlabel metal3 s 0 103096 800 103216 6 master1_wb_adr_o[0]
port 104 nsew signal input
rlabel metal3 s 0 120096 800 120216 6 master1_wb_adr_o[10]
port 105 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 master1_wb_adr_o[11]
port 106 nsew signal input
rlabel metal3 s 0 123088 800 123208 6 master1_wb_adr_o[12]
port 107 nsew signal input
rlabel metal3 s 0 124584 800 124704 6 master1_wb_adr_o[13]
port 108 nsew signal input
rlabel metal3 s 0 126080 800 126200 6 master1_wb_adr_o[14]
port 109 nsew signal input
rlabel metal3 s 0 127576 800 127696 6 master1_wb_adr_o[15]
port 110 nsew signal input
rlabel metal3 s 0 129072 800 129192 6 master1_wb_adr_o[16]
port 111 nsew signal input
rlabel metal3 s 0 130568 800 130688 6 master1_wb_adr_o[17]
port 112 nsew signal input
rlabel metal3 s 0 132064 800 132184 6 master1_wb_adr_o[18]
port 113 nsew signal input
rlabel metal3 s 0 133560 800 133680 6 master1_wb_adr_o[19]
port 114 nsew signal input
rlabel metal3 s 0 105136 800 105256 6 master1_wb_adr_o[1]
port 115 nsew signal input
rlabel metal3 s 0 135056 800 135176 6 master1_wb_adr_o[20]
port 116 nsew signal input
rlabel metal3 s 0 136552 800 136672 6 master1_wb_adr_o[21]
port 117 nsew signal input
rlabel metal3 s 0 138048 800 138168 6 master1_wb_adr_o[22]
port 118 nsew signal input
rlabel metal3 s 0 139680 800 139800 6 master1_wb_adr_o[23]
port 119 nsew signal input
rlabel metal3 s 0 141176 800 141296 6 master1_wb_adr_o[24]
port 120 nsew signal input
rlabel metal3 s 0 142672 800 142792 6 master1_wb_adr_o[25]
port 121 nsew signal input
rlabel metal3 s 0 144168 800 144288 6 master1_wb_adr_o[26]
port 122 nsew signal input
rlabel metal3 s 0 145664 800 145784 6 master1_wb_adr_o[27]
port 123 nsew signal input
rlabel metal3 s 0 107040 800 107160 6 master1_wb_adr_o[2]
port 124 nsew signal input
rlabel metal3 s 0 109080 800 109200 6 master1_wb_adr_o[3]
port 125 nsew signal input
rlabel metal3 s 0 111120 800 111240 6 master1_wb_adr_o[4]
port 126 nsew signal input
rlabel metal3 s 0 112616 800 112736 6 master1_wb_adr_o[5]
port 127 nsew signal input
rlabel metal3 s 0 114112 800 114232 6 master1_wb_adr_o[6]
port 128 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 master1_wb_adr_o[7]
port 129 nsew signal input
rlabel metal3 s 0 117104 800 117224 6 master1_wb_adr_o[8]
port 130 nsew signal input
rlabel metal3 s 0 118600 800 118720 6 master1_wb_adr_o[9]
port 131 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 master1_wb_cyc_o
port 132 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 master1_wb_data_i[0]
port 133 nsew signal output
rlabel metal3 s 0 120640 800 120760 6 master1_wb_data_i[10]
port 134 nsew signal output
rlabel metal3 s 0 122136 800 122256 6 master1_wb_data_i[11]
port 135 nsew signal output
rlabel metal3 s 0 123632 800 123752 6 master1_wb_data_i[12]
port 136 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 master1_wb_data_i[13]
port 137 nsew signal output
rlabel metal3 s 0 126624 800 126744 6 master1_wb_data_i[14]
port 138 nsew signal output
rlabel metal3 s 0 128120 800 128240 6 master1_wb_data_i[15]
port 139 nsew signal output
rlabel metal3 s 0 129616 800 129736 6 master1_wb_data_i[16]
port 140 nsew signal output
rlabel metal3 s 0 131112 800 131232 6 master1_wb_data_i[17]
port 141 nsew signal output
rlabel metal3 s 0 132608 800 132728 6 master1_wb_data_i[18]
port 142 nsew signal output
rlabel metal3 s 0 134104 800 134224 6 master1_wb_data_i[19]
port 143 nsew signal output
rlabel metal3 s 0 105544 800 105664 6 master1_wb_data_i[1]
port 144 nsew signal output
rlabel metal3 s 0 135600 800 135720 6 master1_wb_data_i[20]
port 145 nsew signal output
rlabel metal3 s 0 137096 800 137216 6 master1_wb_data_i[21]
port 146 nsew signal output
rlabel metal3 s 0 138592 800 138712 6 master1_wb_data_i[22]
port 147 nsew signal output
rlabel metal3 s 0 140088 800 140208 6 master1_wb_data_i[23]
port 148 nsew signal output
rlabel metal3 s 0 141584 800 141704 6 master1_wb_data_i[24]
port 149 nsew signal output
rlabel metal3 s 0 143080 800 143200 6 master1_wb_data_i[25]
port 150 nsew signal output
rlabel metal3 s 0 144576 800 144696 6 master1_wb_data_i[26]
port 151 nsew signal output
rlabel metal3 s 0 146072 800 146192 6 master1_wb_data_i[27]
port 152 nsew signal output
rlabel metal3 s 0 147160 800 147280 6 master1_wb_data_i[28]
port 153 nsew signal output
rlabel metal3 s 0 148112 800 148232 6 master1_wb_data_i[29]
port 154 nsew signal output
rlabel metal3 s 0 107584 800 107704 6 master1_wb_data_i[2]
port 155 nsew signal output
rlabel metal3 s 0 149064 800 149184 6 master1_wb_data_i[30]
port 156 nsew signal output
rlabel metal3 s 0 150152 800 150272 6 master1_wb_data_i[31]
port 157 nsew signal output
rlabel metal3 s 0 109624 800 109744 6 master1_wb_data_i[3]
port 158 nsew signal output
rlabel metal3 s 0 111664 800 111784 6 master1_wb_data_i[4]
port 159 nsew signal output
rlabel metal3 s 0 113160 800 113280 6 master1_wb_data_i[5]
port 160 nsew signal output
rlabel metal3 s 0 114656 800 114776 6 master1_wb_data_i[6]
port 161 nsew signal output
rlabel metal3 s 0 116152 800 116272 6 master1_wb_data_i[7]
port 162 nsew signal output
rlabel metal3 s 0 117648 800 117768 6 master1_wb_data_i[8]
port 163 nsew signal output
rlabel metal3 s 0 119144 800 119264 6 master1_wb_data_i[9]
port 164 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 master1_wb_data_o[0]
port 165 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 master1_wb_data_o[10]
port 166 nsew signal input
rlabel metal3 s 0 122544 800 122664 6 master1_wb_data_o[11]
port 167 nsew signal input
rlabel metal3 s 0 124176 800 124296 6 master1_wb_data_o[12]
port 168 nsew signal input
rlabel metal3 s 0 125672 800 125792 6 master1_wb_data_o[13]
port 169 nsew signal input
rlabel metal3 s 0 127168 800 127288 6 master1_wb_data_o[14]
port 170 nsew signal input
rlabel metal3 s 0 128664 800 128784 6 master1_wb_data_o[15]
port 171 nsew signal input
rlabel metal3 s 0 130160 800 130280 6 master1_wb_data_o[16]
port 172 nsew signal input
rlabel metal3 s 0 131656 800 131776 6 master1_wb_data_o[17]
port 173 nsew signal input
rlabel metal3 s 0 133152 800 133272 6 master1_wb_data_o[18]
port 174 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 master1_wb_data_o[19]
port 175 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 master1_wb_data_o[1]
port 176 nsew signal input
rlabel metal3 s 0 136144 800 136264 6 master1_wb_data_o[20]
port 177 nsew signal input
rlabel metal3 s 0 137640 800 137760 6 master1_wb_data_o[21]
port 178 nsew signal input
rlabel metal3 s 0 139136 800 139256 6 master1_wb_data_o[22]
port 179 nsew signal input
rlabel metal3 s 0 140632 800 140752 6 master1_wb_data_o[23]
port 180 nsew signal input
rlabel metal3 s 0 142128 800 142248 6 master1_wb_data_o[24]
port 181 nsew signal input
rlabel metal3 s 0 143624 800 143744 6 master1_wb_data_o[25]
port 182 nsew signal input
rlabel metal3 s 0 145120 800 145240 6 master1_wb_data_o[26]
port 183 nsew signal input
rlabel metal3 s 0 146616 800 146736 6 master1_wb_data_o[27]
port 184 nsew signal input
rlabel metal3 s 0 147568 800 147688 6 master1_wb_data_o[28]
port 185 nsew signal input
rlabel metal3 s 0 148656 800 148776 6 master1_wb_data_o[29]
port 186 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 master1_wb_data_o[2]
port 187 nsew signal input
rlabel metal3 s 0 149608 800 149728 6 master1_wb_data_o[30]
port 188 nsew signal input
rlabel metal3 s 0 150560 800 150680 6 master1_wb_data_o[31]
port 189 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 master1_wb_data_o[3]
port 190 nsew signal input
rlabel metal3 s 0 112072 800 112192 6 master1_wb_data_o[4]
port 191 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 master1_wb_data_o[5]
port 192 nsew signal input
rlabel metal3 s 0 115064 800 115184 6 master1_wb_data_o[6]
port 193 nsew signal input
rlabel metal3 s 0 116560 800 116680 6 master1_wb_data_o[7]
port 194 nsew signal input
rlabel metal3 s 0 118056 800 118176 6 master1_wb_data_o[8]
port 195 nsew signal input
rlabel metal3 s 0 119552 800 119672 6 master1_wb_data_o[9]
port 196 nsew signal input
rlabel metal3 s 0 101056 800 101176 6 master1_wb_error_i
port 197 nsew signal output
rlabel metal3 s 0 104592 800 104712 6 master1_wb_sel_o[0]
port 198 nsew signal input
rlabel metal3 s 0 106632 800 106752 6 master1_wb_sel_o[1]
port 199 nsew signal input
rlabel metal3 s 0 108672 800 108792 6 master1_wb_sel_o[2]
port 200 nsew signal input
rlabel metal3 s 0 110576 800 110696 6 master1_wb_sel_o[3]
port 201 nsew signal input
rlabel metal3 s 0 101600 800 101720 6 master1_wb_stall_i
port 202 nsew signal output
rlabel metal3 s 0 102144 800 102264 6 master1_wb_stb_o
port 203 nsew signal input
rlabel metal3 s 0 102552 800 102672 6 master1_wb_we_o
port 204 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 master2_wb_ack_i
port 205 nsew signal output
rlabel metal3 s 0 52096 800 52216 6 master2_wb_adr_o[0]
port 206 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 master2_wb_adr_o[10]
port 207 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 master2_wb_adr_o[11]
port 208 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 master2_wb_adr_o[12]
port 209 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 master2_wb_adr_o[13]
port 210 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 master2_wb_adr_o[14]
port 211 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 master2_wb_adr_o[15]
port 212 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 master2_wb_adr_o[16]
port 213 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 master2_wb_adr_o[17]
port 214 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 master2_wb_adr_o[18]
port 215 nsew signal input
rlabel metal3 s 0 82560 800 82680 6 master2_wb_adr_o[19]
port 216 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 master2_wb_adr_o[1]
port 217 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 master2_wb_adr_o[20]
port 218 nsew signal input
rlabel metal3 s 0 85552 800 85672 6 master2_wb_adr_o[21]
port 219 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 master2_wb_adr_o[22]
port 220 nsew signal input
rlabel metal3 s 0 88544 800 88664 6 master2_wb_adr_o[23]
port 221 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 master2_wb_adr_o[24]
port 222 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 master2_wb_adr_o[25]
port 223 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 master2_wb_adr_o[26]
port 224 nsew signal input
rlabel metal3 s 0 94664 800 94784 6 master2_wb_adr_o[27]
port 225 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 master2_wb_adr_o[2]
port 226 nsew signal input
rlabel metal3 s 0 58080 800 58200 6 master2_wb_adr_o[3]
port 227 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 master2_wb_adr_o[4]
port 228 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 master2_wb_adr_o[5]
port 229 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 master2_wb_adr_o[6]
port 230 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 master2_wb_adr_o[7]
port 231 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 master2_wb_adr_o[8]
port 232 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 master2_wb_adr_o[9]
port 233 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 master2_wb_cyc_o
port 234 nsew signal input
rlabel metal3 s 0 52640 800 52760 6 master2_wb_data_i[0]
port 235 nsew signal output
rlabel metal3 s 0 69640 800 69760 6 master2_wb_data_i[10]
port 236 nsew signal output
rlabel metal3 s 0 71136 800 71256 6 master2_wb_data_i[11]
port 237 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 master2_wb_data_i[12]
port 238 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 master2_wb_data_i[13]
port 239 nsew signal output
rlabel metal3 s 0 75624 800 75744 6 master2_wb_data_i[14]
port 240 nsew signal output
rlabel metal3 s 0 77120 800 77240 6 master2_wb_data_i[15]
port 241 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 master2_wb_data_i[16]
port 242 nsew signal output
rlabel metal3 s 0 80112 800 80232 6 master2_wb_data_i[17]
port 243 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 master2_wb_data_i[18]
port 244 nsew signal output
rlabel metal3 s 0 83104 800 83224 6 master2_wb_data_i[19]
port 245 nsew signal output
rlabel metal3 s 0 54544 800 54664 6 master2_wb_data_i[1]
port 246 nsew signal output
rlabel metal3 s 0 84600 800 84720 6 master2_wb_data_i[20]
port 247 nsew signal output
rlabel metal3 s 0 86096 800 86216 6 master2_wb_data_i[21]
port 248 nsew signal output
rlabel metal3 s 0 87592 800 87712 6 master2_wb_data_i[22]
port 249 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 master2_wb_data_i[23]
port 250 nsew signal output
rlabel metal3 s 0 90584 800 90704 6 master2_wb_data_i[24]
port 251 nsew signal output
rlabel metal3 s 0 92080 800 92200 6 master2_wb_data_i[25]
port 252 nsew signal output
rlabel metal3 s 0 93576 800 93696 6 master2_wb_data_i[26]
port 253 nsew signal output
rlabel metal3 s 0 95072 800 95192 6 master2_wb_data_i[27]
port 254 nsew signal output
rlabel metal3 s 0 96160 800 96280 6 master2_wb_data_i[28]
port 255 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 master2_wb_data_i[29]
port 256 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 master2_wb_data_i[2]
port 257 nsew signal output
rlabel metal3 s 0 98064 800 98184 6 master2_wb_data_i[30]
port 258 nsew signal output
rlabel metal3 s 0 99152 800 99272 6 master2_wb_data_i[31]
port 259 nsew signal output
rlabel metal3 s 0 58624 800 58744 6 master2_wb_data_i[3]
port 260 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 master2_wb_data_i[4]
port 261 nsew signal output
rlabel metal3 s 0 62160 800 62280 6 master2_wb_data_i[5]
port 262 nsew signal output
rlabel metal3 s 0 63656 800 63776 6 master2_wb_data_i[6]
port 263 nsew signal output
rlabel metal3 s 0 65152 800 65272 6 master2_wb_data_i[7]
port 264 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 master2_wb_data_i[8]
port 265 nsew signal output
rlabel metal3 s 0 68144 800 68264 6 master2_wb_data_i[9]
port 266 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 master2_wb_data_o[0]
port 267 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 master2_wb_data_o[10]
port 268 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 master2_wb_data_o[11]
port 269 nsew signal input
rlabel metal3 s 0 73040 800 73160 6 master2_wb_data_o[12]
port 270 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 master2_wb_data_o[13]
port 271 nsew signal input
rlabel metal3 s 0 76032 800 76152 6 master2_wb_data_o[14]
port 272 nsew signal input
rlabel metal3 s 0 77664 800 77784 6 master2_wb_data_o[15]
port 273 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 master2_wb_data_o[16]
port 274 nsew signal input
rlabel metal3 s 0 80656 800 80776 6 master2_wb_data_o[17]
port 275 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 master2_wb_data_o[18]
port 276 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 master2_wb_data_o[19]
port 277 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 master2_wb_data_o[1]
port 278 nsew signal input
rlabel metal3 s 0 85144 800 85264 6 master2_wb_data_o[20]
port 279 nsew signal input
rlabel metal3 s 0 86640 800 86760 6 master2_wb_data_o[21]
port 280 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 master2_wb_data_o[22]
port 281 nsew signal input
rlabel metal3 s 0 89632 800 89752 6 master2_wb_data_o[23]
port 282 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 master2_wb_data_o[24]
port 283 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 master2_wb_data_o[25]
port 284 nsew signal input
rlabel metal3 s 0 94120 800 94240 6 master2_wb_data_o[26]
port 285 nsew signal input
rlabel metal3 s 0 95616 800 95736 6 master2_wb_data_o[27]
port 286 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 master2_wb_data_o[28]
port 287 nsew signal input
rlabel metal3 s 0 97656 800 97776 6 master2_wb_data_o[29]
port 288 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 master2_wb_data_o[2]
port 289 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 master2_wb_data_o[30]
port 290 nsew signal input
rlabel metal3 s 0 99560 800 99680 6 master2_wb_data_o[31]
port 291 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 master2_wb_data_o[3]
port 292 nsew signal input
rlabel metal3 s 0 61072 800 61192 6 master2_wb_data_o[4]
port 293 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 master2_wb_data_o[5]
port 294 nsew signal input
rlabel metal3 s 0 64064 800 64184 6 master2_wb_data_o[6]
port 295 nsew signal input
rlabel metal3 s 0 65560 800 65680 6 master2_wb_data_o[7]
port 296 nsew signal input
rlabel metal3 s 0 67056 800 67176 6 master2_wb_data_o[8]
port 297 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 master2_wb_data_o[9]
port 298 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 master2_wb_error_i
port 299 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 master2_wb_sel_o[0]
port 300 nsew signal input
rlabel metal3 s 0 55632 800 55752 6 master2_wb_sel_o[1]
port 301 nsew signal input
rlabel metal3 s 0 57536 800 57656 6 master2_wb_sel_o[2]
port 302 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 master2_wb_sel_o[3]
port 303 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 master2_wb_stall_i
port 304 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 master2_wb_stb_o
port 305 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 master2_wb_we_o
port 306 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 probe_master0_currentSlave[0]
port 307 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 probe_master0_currentSlave[1]
port 308 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 probe_master0_currentSlave[2]
port 309 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 probe_master1_currentSlave[0]
port 310 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 probe_master1_currentSlave[1]
port 311 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 probe_master1_currentSlave[2]
port 312 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 probe_master2_currentSlave[0]
port 313 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 probe_master2_currentSlave[1]
port 314 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 probe_master2_currentSlave[2]
port 315 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 probe_master3_currentSlave[0]
port 316 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 probe_master3_currentSlave[1]
port 317 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 probe_master3_currentSlave[2]
port 318 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 probe_slave0_currentMaster[0]
port 319 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 probe_slave0_currentMaster[1]
port 320 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 probe_slave1_currentMaster[0]
port 321 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 probe_slave1_currentMaster[1]
port 322 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 probe_slave2_currentMaster[0]
port 323 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 probe_slave2_currentMaster[1]
port 324 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 probe_slave3_currentMaster[0]
port 325 nsew signal output
rlabel metal2 s 10230 0 10286 800 6 probe_slave3_currentMaster[1]
port 326 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 probe_slave4_currentMaster[0]
port 327 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 probe_slave4_currentMaster[1]
port 328 nsew signal output
rlabel metal3 s 0 151104 800 151224 6 slave0_wb_ack_o
port 329 nsew signal input
rlabel metal3 s 0 154096 800 154216 6 slave0_wb_adr_i[0]
port 330 nsew signal output
rlabel metal3 s 0 171096 800 171216 6 slave0_wb_adr_i[10]
port 331 nsew signal output
rlabel metal3 s 0 172592 800 172712 6 slave0_wb_adr_i[11]
port 332 nsew signal output
rlabel metal3 s 0 174088 800 174208 6 slave0_wb_adr_i[12]
port 333 nsew signal output
rlabel metal3 s 0 175584 800 175704 6 slave0_wb_adr_i[13]
port 334 nsew signal output
rlabel metal3 s 0 177080 800 177200 6 slave0_wb_adr_i[14]
port 335 nsew signal output
rlabel metal3 s 0 178576 800 178696 6 slave0_wb_adr_i[15]
port 336 nsew signal output
rlabel metal3 s 0 180072 800 180192 6 slave0_wb_adr_i[16]
port 337 nsew signal output
rlabel metal3 s 0 181568 800 181688 6 slave0_wb_adr_i[17]
port 338 nsew signal output
rlabel metal3 s 0 183064 800 183184 6 slave0_wb_adr_i[18]
port 339 nsew signal output
rlabel metal3 s 0 184560 800 184680 6 slave0_wb_adr_i[19]
port 340 nsew signal output
rlabel metal3 s 0 156136 800 156256 6 slave0_wb_adr_i[1]
port 341 nsew signal output
rlabel metal3 s 0 186192 800 186312 6 slave0_wb_adr_i[20]
port 342 nsew signal output
rlabel metal3 s 0 187688 800 187808 6 slave0_wb_adr_i[21]
port 343 nsew signal output
rlabel metal3 s 0 189184 800 189304 6 slave0_wb_adr_i[22]
port 344 nsew signal output
rlabel metal3 s 0 190680 800 190800 6 slave0_wb_adr_i[23]
port 345 nsew signal output
rlabel metal3 s 0 158176 800 158296 6 slave0_wb_adr_i[2]
port 346 nsew signal output
rlabel metal3 s 0 160080 800 160200 6 slave0_wb_adr_i[3]
port 347 nsew signal output
rlabel metal3 s 0 162120 800 162240 6 slave0_wb_adr_i[4]
port 348 nsew signal output
rlabel metal3 s 0 163616 800 163736 6 slave0_wb_adr_i[5]
port 349 nsew signal output
rlabel metal3 s 0 165112 800 165232 6 slave0_wb_adr_i[6]
port 350 nsew signal output
rlabel metal3 s 0 166608 800 166728 6 slave0_wb_adr_i[7]
port 351 nsew signal output
rlabel metal3 s 0 168104 800 168224 6 slave0_wb_adr_i[8]
port 352 nsew signal output
rlabel metal3 s 0 169600 800 169720 6 slave0_wb_adr_i[9]
port 353 nsew signal output
rlabel metal3 s 0 151648 800 151768 6 slave0_wb_cyc_i
port 354 nsew signal output
rlabel metal3 s 0 154640 800 154760 6 slave0_wb_data_i[0]
port 355 nsew signal output
rlabel metal3 s 0 171640 800 171760 6 slave0_wb_data_i[10]
port 356 nsew signal output
rlabel metal3 s 0 173136 800 173256 6 slave0_wb_data_i[11]
port 357 nsew signal output
rlabel metal3 s 0 174632 800 174752 6 slave0_wb_data_i[12]
port 358 nsew signal output
rlabel metal3 s 0 176128 800 176248 6 slave0_wb_data_i[13]
port 359 nsew signal output
rlabel metal3 s 0 177624 800 177744 6 slave0_wb_data_i[14]
port 360 nsew signal output
rlabel metal3 s 0 179120 800 179240 6 slave0_wb_data_i[15]
port 361 nsew signal output
rlabel metal3 s 0 180616 800 180736 6 slave0_wb_data_i[16]
port 362 nsew signal output
rlabel metal3 s 0 182112 800 182232 6 slave0_wb_data_i[17]
port 363 nsew signal output
rlabel metal3 s 0 183608 800 183728 6 slave0_wb_data_i[18]
port 364 nsew signal output
rlabel metal3 s 0 185104 800 185224 6 slave0_wb_data_i[19]
port 365 nsew signal output
rlabel metal3 s 0 156680 800 156800 6 slave0_wb_data_i[1]
port 366 nsew signal output
rlabel metal3 s 0 186600 800 186720 6 slave0_wb_data_i[20]
port 367 nsew signal output
rlabel metal3 s 0 188096 800 188216 6 slave0_wb_data_i[21]
port 368 nsew signal output
rlabel metal3 s 0 189592 800 189712 6 slave0_wb_data_i[22]
port 369 nsew signal output
rlabel metal3 s 0 191088 800 191208 6 slave0_wb_data_i[23]
port 370 nsew signal output
rlabel metal3 s 0 192176 800 192296 6 slave0_wb_data_i[24]
port 371 nsew signal output
rlabel metal3 s 0 193128 800 193248 6 slave0_wb_data_i[25]
port 372 nsew signal output
rlabel metal3 s 0 194080 800 194200 6 slave0_wb_data_i[26]
port 373 nsew signal output
rlabel metal3 s 0 195168 800 195288 6 slave0_wb_data_i[27]
port 374 nsew signal output
rlabel metal3 s 0 196120 800 196240 6 slave0_wb_data_i[28]
port 375 nsew signal output
rlabel metal3 s 0 197072 800 197192 6 slave0_wb_data_i[29]
port 376 nsew signal output
rlabel metal3 s 0 158584 800 158704 6 slave0_wb_data_i[2]
port 377 nsew signal output
rlabel metal3 s 0 198160 800 198280 6 slave0_wb_data_i[30]
port 378 nsew signal output
rlabel metal3 s 0 199112 800 199232 6 slave0_wb_data_i[31]
port 379 nsew signal output
rlabel metal3 s 0 160624 800 160744 6 slave0_wb_data_i[3]
port 380 nsew signal output
rlabel metal3 s 0 162664 800 162784 6 slave0_wb_data_i[4]
port 381 nsew signal output
rlabel metal3 s 0 164160 800 164280 6 slave0_wb_data_i[5]
port 382 nsew signal output
rlabel metal3 s 0 165656 800 165776 6 slave0_wb_data_i[6]
port 383 nsew signal output
rlabel metal3 s 0 167152 800 167272 6 slave0_wb_data_i[7]
port 384 nsew signal output
rlabel metal3 s 0 168648 800 168768 6 slave0_wb_data_i[8]
port 385 nsew signal output
rlabel metal3 s 0 170144 800 170264 6 slave0_wb_data_i[9]
port 386 nsew signal output
rlabel metal3 s 0 155184 800 155304 6 slave0_wb_data_o[0]
port 387 nsew signal input
rlabel metal3 s 0 172184 800 172304 6 slave0_wb_data_o[10]
port 388 nsew signal input
rlabel metal3 s 0 173680 800 173800 6 slave0_wb_data_o[11]
port 389 nsew signal input
rlabel metal3 s 0 175176 800 175296 6 slave0_wb_data_o[12]
port 390 nsew signal input
rlabel metal3 s 0 176672 800 176792 6 slave0_wb_data_o[13]
port 391 nsew signal input
rlabel metal3 s 0 178168 800 178288 6 slave0_wb_data_o[14]
port 392 nsew signal input
rlabel metal3 s 0 179664 800 179784 6 slave0_wb_data_o[15]
port 393 nsew signal input
rlabel metal3 s 0 181160 800 181280 6 slave0_wb_data_o[16]
port 394 nsew signal input
rlabel metal3 s 0 182656 800 182776 6 slave0_wb_data_o[17]
port 395 nsew signal input
rlabel metal3 s 0 184152 800 184272 6 slave0_wb_data_o[18]
port 396 nsew signal input
rlabel metal3 s 0 185648 800 185768 6 slave0_wb_data_o[19]
port 397 nsew signal input
rlabel metal3 s 0 157088 800 157208 6 slave0_wb_data_o[1]
port 398 nsew signal input
rlabel metal3 s 0 187144 800 187264 6 slave0_wb_data_o[20]
port 399 nsew signal input
rlabel metal3 s 0 188640 800 188760 6 slave0_wb_data_o[21]
port 400 nsew signal input
rlabel metal3 s 0 190136 800 190256 6 slave0_wb_data_o[22]
port 401 nsew signal input
rlabel metal3 s 0 191632 800 191752 6 slave0_wb_data_o[23]
port 402 nsew signal input
rlabel metal3 s 0 192584 800 192704 6 slave0_wb_data_o[24]
port 403 nsew signal input
rlabel metal3 s 0 193672 800 193792 6 slave0_wb_data_o[25]
port 404 nsew signal input
rlabel metal3 s 0 194624 800 194744 6 slave0_wb_data_o[26]
port 405 nsew signal input
rlabel metal3 s 0 195576 800 195696 6 slave0_wb_data_o[27]
port 406 nsew signal input
rlabel metal3 s 0 196664 800 196784 6 slave0_wb_data_o[28]
port 407 nsew signal input
rlabel metal3 s 0 197616 800 197736 6 slave0_wb_data_o[29]
port 408 nsew signal input
rlabel metal3 s 0 159128 800 159248 6 slave0_wb_data_o[2]
port 409 nsew signal input
rlabel metal3 s 0 198568 800 198688 6 slave0_wb_data_o[30]
port 410 nsew signal input
rlabel metal3 s 0 199656 800 199776 6 slave0_wb_data_o[31]
port 411 nsew signal input
rlabel metal3 s 0 161168 800 161288 6 slave0_wb_data_o[3]
port 412 nsew signal input
rlabel metal3 s 0 163072 800 163192 6 slave0_wb_data_o[4]
port 413 nsew signal input
rlabel metal3 s 0 164568 800 164688 6 slave0_wb_data_o[5]
port 414 nsew signal input
rlabel metal3 s 0 166064 800 166184 6 slave0_wb_data_o[6]
port 415 nsew signal input
rlabel metal3 s 0 167560 800 167680 6 slave0_wb_data_o[7]
port 416 nsew signal input
rlabel metal3 s 0 169056 800 169176 6 slave0_wb_data_o[8]
port 417 nsew signal input
rlabel metal3 s 0 170688 800 170808 6 slave0_wb_data_o[9]
port 418 nsew signal input
rlabel metal3 s 0 152056 800 152176 6 slave0_wb_error_o
port 419 nsew signal input
rlabel metal3 s 0 155592 800 155712 6 slave0_wb_sel_i[0]
port 420 nsew signal output
rlabel metal3 s 0 157632 800 157752 6 slave0_wb_sel_i[1]
port 421 nsew signal output
rlabel metal3 s 0 159672 800 159792 6 slave0_wb_sel_i[2]
port 422 nsew signal output
rlabel metal3 s 0 161576 800 161696 6 slave0_wb_sel_i[3]
port 423 nsew signal output
rlabel metal3 s 0 152600 800 152720 6 slave0_wb_stall_o
port 424 nsew signal input
rlabel metal3 s 0 153144 800 153264 6 slave0_wb_stb_i
port 425 nsew signal output
rlabel metal3 s 0 153552 800 153672 6 slave0_wb_we_i
port 426 nsew signal output
rlabel metal3 s 0 144 800 264 6 slave1_wb_ack_o
port 427 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 slave1_wb_adr_i[0]
port 428 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 slave1_wb_adr_i[10]
port 429 nsew signal output
rlabel metal3 s 0 21632 800 21752 6 slave1_wb_adr_i[11]
port 430 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 slave1_wb_adr_i[12]
port 431 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 slave1_wb_adr_i[13]
port 432 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 slave1_wb_adr_i[14]
port 433 nsew signal output
rlabel metal3 s 0 27616 800 27736 6 slave1_wb_adr_i[15]
port 434 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 slave1_wb_adr_i[16]
port 435 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 slave1_wb_adr_i[17]
port 436 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 slave1_wb_adr_i[18]
port 437 nsew signal output
rlabel metal3 s 0 33600 800 33720 6 slave1_wb_adr_i[19]
port 438 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 slave1_wb_adr_i[1]
port 439 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 slave1_wb_adr_i[20]
port 440 nsew signal output
rlabel metal3 s 0 36592 800 36712 6 slave1_wb_adr_i[21]
port 441 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 slave1_wb_adr_i[22]
port 442 nsew signal output
rlabel metal3 s 0 39584 800 39704 6 slave1_wb_adr_i[23]
port 443 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 slave1_wb_adr_i[2]
port 444 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 slave1_wb_adr_i[3]
port 445 nsew signal output
rlabel metal3 s 0 11024 800 11144 6 slave1_wb_adr_i[4]
port 446 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 slave1_wb_adr_i[5]
port 447 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 slave1_wb_adr_i[6]
port 448 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 slave1_wb_adr_i[7]
port 449 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 slave1_wb_adr_i[8]
port 450 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 slave1_wb_adr_i[9]
port 451 nsew signal output
rlabel metal3 s 0 552 800 672 6 slave1_wb_cyc_i
port 452 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 slave1_wb_data_i[0]
port 453 nsew signal output
rlabel metal3 s 0 20544 800 20664 6 slave1_wb_data_i[10]
port 454 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 slave1_wb_data_i[11]
port 455 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 slave1_wb_data_i[12]
port 456 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 slave1_wb_data_i[13]
port 457 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 slave1_wb_data_i[14]
port 458 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 slave1_wb_data_i[15]
port 459 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 slave1_wb_data_i[16]
port 460 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 slave1_wb_data_i[17]
port 461 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 slave1_wb_data_i[18]
port 462 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 slave1_wb_data_i[19]
port 463 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 slave1_wb_data_i[1]
port 464 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 slave1_wb_data_i[20]
port 465 nsew signal output
rlabel metal3 s 0 37136 800 37256 6 slave1_wb_data_i[21]
port 466 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 slave1_wb_data_i[22]
port 467 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 slave1_wb_data_i[23]
port 468 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 slave1_wb_data_i[24]
port 469 nsew signal output
rlabel metal3 s 0 42032 800 42152 6 slave1_wb_data_i[25]
port 470 nsew signal output
rlabel metal3 s 0 43120 800 43240 6 slave1_wb_data_i[26]
port 471 nsew signal output
rlabel metal3 s 0 44072 800 44192 6 slave1_wb_data_i[27]
port 472 nsew signal output
rlabel metal3 s 0 45024 800 45144 6 slave1_wb_data_i[28]
port 473 nsew signal output
rlabel metal3 s 0 46112 800 46232 6 slave1_wb_data_i[29]
port 474 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 slave1_wb_data_i[2]
port 475 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 slave1_wb_data_i[30]
port 476 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 slave1_wb_data_i[31]
port 477 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 slave1_wb_data_i[3]
port 478 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 slave1_wb_data_i[4]
port 479 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 slave1_wb_data_i[5]
port 480 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 slave1_wb_data_i[6]
port 481 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 slave1_wb_data_i[7]
port 482 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 slave1_wb_data_i[8]
port 483 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 slave1_wb_data_i[9]
port 484 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 slave1_wb_data_o[0]
port 485 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 slave1_wb_data_o[10]
port 486 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 slave1_wb_data_o[11]
port 487 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 slave1_wb_data_o[12]
port 488 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 slave1_wb_data_o[13]
port 489 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 slave1_wb_data_o[14]
port 490 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 slave1_wb_data_o[15]
port 491 nsew signal input
rlabel metal3 s 0 30064 800 30184 6 slave1_wb_data_o[16]
port 492 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 slave1_wb_data_o[17]
port 493 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 slave1_wb_data_o[18]
port 494 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 slave1_wb_data_o[19]
port 495 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 slave1_wb_data_o[1]
port 496 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 slave1_wb_data_o[20]
port 497 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 slave1_wb_data_o[21]
port 498 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 slave1_wb_data_o[22]
port 499 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 slave1_wb_data_o[23]
port 500 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 slave1_wb_data_o[24]
port 501 nsew signal input
rlabel metal3 s 0 42576 800 42696 6 slave1_wb_data_o[25]
port 502 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 slave1_wb_data_o[26]
port 503 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 slave1_wb_data_o[27]
port 504 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 slave1_wb_data_o[28]
port 505 nsew signal input
rlabel metal3 s 0 46656 800 46776 6 slave1_wb_data_o[29]
port 506 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 slave1_wb_data_o[2]
port 507 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 slave1_wb_data_o[30]
port 508 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 slave1_wb_data_o[31]
port 509 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 slave1_wb_data_o[3]
port 510 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 slave1_wb_data_o[4]
port 511 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 slave1_wb_data_o[5]
port 512 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 slave1_wb_data_o[6]
port 513 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 slave1_wb_data_o[7]
port 514 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 slave1_wb_data_o[8]
port 515 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 slave1_wb_data_o[9]
port 516 nsew signal input
rlabel metal3 s 0 1096 800 1216 6 slave1_wb_error_o
port 517 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 slave1_wb_sel_i[0]
port 518 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 slave1_wb_sel_i[1]
port 519 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 slave1_wb_sel_i[2]
port 520 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 slave1_wb_sel_i[3]
port 521 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 slave1_wb_stall_o
port 522 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 slave1_wb_stb_i
port 523 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 slave1_wb_we_i
port 524 nsew signal output
rlabel metal2 s 294 199200 350 200000 6 slave2_wb_ack_o
port 525 nsew signal input
rlabel metal2 s 4526 199200 4582 200000 6 slave2_wb_adr_i[0]
port 526 nsew signal output
rlabel metal2 s 28814 199200 28870 200000 6 slave2_wb_adr_i[10]
port 527 nsew signal output
rlabel metal2 s 30930 199200 30986 200000 6 slave2_wb_adr_i[11]
port 528 nsew signal output
rlabel metal2 s 33138 199200 33194 200000 6 slave2_wb_adr_i[12]
port 529 nsew signal output
rlabel metal2 s 35254 199200 35310 200000 6 slave2_wb_adr_i[13]
port 530 nsew signal output
rlabel metal2 s 37370 199200 37426 200000 6 slave2_wb_adr_i[14]
port 531 nsew signal output
rlabel metal2 s 39578 199200 39634 200000 6 slave2_wb_adr_i[15]
port 532 nsew signal output
rlabel metal2 s 41694 199200 41750 200000 6 slave2_wb_adr_i[16]
port 533 nsew signal output
rlabel metal2 s 43810 199200 43866 200000 6 slave2_wb_adr_i[17]
port 534 nsew signal output
rlabel metal2 s 45926 199200 45982 200000 6 slave2_wb_adr_i[18]
port 535 nsew signal output
rlabel metal2 s 48134 199200 48190 200000 6 slave2_wb_adr_i[19]
port 536 nsew signal output
rlabel metal2 s 7378 199200 7434 200000 6 slave2_wb_adr_i[1]
port 537 nsew signal output
rlabel metal2 s 50250 199200 50306 200000 6 slave2_wb_adr_i[20]
port 538 nsew signal output
rlabel metal2 s 52366 199200 52422 200000 6 slave2_wb_adr_i[21]
port 539 nsew signal output
rlabel metal2 s 54574 199200 54630 200000 6 slave2_wb_adr_i[22]
port 540 nsew signal output
rlabel metal2 s 56690 199200 56746 200000 6 slave2_wb_adr_i[23]
port 541 nsew signal output
rlabel metal2 s 10230 199200 10286 200000 6 slave2_wb_adr_i[2]
port 542 nsew signal output
rlabel metal2 s 13082 199200 13138 200000 6 slave2_wb_adr_i[3]
port 543 nsew signal output
rlabel metal2 s 15934 199200 15990 200000 6 slave2_wb_adr_i[4]
port 544 nsew signal output
rlabel metal2 s 18142 199200 18198 200000 6 slave2_wb_adr_i[5]
port 545 nsew signal output
rlabel metal2 s 20258 199200 20314 200000 6 slave2_wb_adr_i[6]
port 546 nsew signal output
rlabel metal2 s 22374 199200 22430 200000 6 slave2_wb_adr_i[7]
port 547 nsew signal output
rlabel metal2 s 24582 199200 24638 200000 6 slave2_wb_adr_i[8]
port 548 nsew signal output
rlabel metal2 s 26698 199200 26754 200000 6 slave2_wb_adr_i[9]
port 549 nsew signal output
rlabel metal2 s 938 199200 994 200000 6 slave2_wb_cyc_i
port 550 nsew signal output
rlabel metal2 s 5262 199200 5318 200000 6 slave2_wb_data_i[0]
port 551 nsew signal output
rlabel metal2 s 29550 199200 29606 200000 6 slave2_wb_data_i[10]
port 552 nsew signal output
rlabel metal2 s 31666 199200 31722 200000 6 slave2_wb_data_i[11]
port 553 nsew signal output
rlabel metal2 s 33782 199200 33838 200000 6 slave2_wb_data_i[12]
port 554 nsew signal output
rlabel metal2 s 35990 199200 36046 200000 6 slave2_wb_data_i[13]
port 555 nsew signal output
rlabel metal2 s 38106 199200 38162 200000 6 slave2_wb_data_i[14]
port 556 nsew signal output
rlabel metal2 s 40222 199200 40278 200000 6 slave2_wb_data_i[15]
port 557 nsew signal output
rlabel metal2 s 42430 199200 42486 200000 6 slave2_wb_data_i[16]
port 558 nsew signal output
rlabel metal2 s 44546 199200 44602 200000 6 slave2_wb_data_i[17]
port 559 nsew signal output
rlabel metal2 s 46662 199200 46718 200000 6 slave2_wb_data_i[18]
port 560 nsew signal output
rlabel metal2 s 48870 199200 48926 200000 6 slave2_wb_data_i[19]
port 561 nsew signal output
rlabel metal2 s 8114 199200 8170 200000 6 slave2_wb_data_i[1]
port 562 nsew signal output
rlabel metal2 s 50986 199200 51042 200000 6 slave2_wb_data_i[20]
port 563 nsew signal output
rlabel metal2 s 53102 199200 53158 200000 6 slave2_wb_data_i[21]
port 564 nsew signal output
rlabel metal2 s 55218 199200 55274 200000 6 slave2_wb_data_i[22]
port 565 nsew signal output
rlabel metal2 s 57426 199200 57482 200000 6 slave2_wb_data_i[23]
port 566 nsew signal output
rlabel metal2 s 58806 199200 58862 200000 6 slave2_wb_data_i[24]
port 567 nsew signal output
rlabel metal2 s 60278 199200 60334 200000 6 slave2_wb_data_i[25]
port 568 nsew signal output
rlabel metal2 s 61658 199200 61714 200000 6 slave2_wb_data_i[26]
port 569 nsew signal output
rlabel metal2 s 63130 199200 63186 200000 6 slave2_wb_data_i[27]
port 570 nsew signal output
rlabel metal2 s 64510 199200 64566 200000 6 slave2_wb_data_i[28]
port 571 nsew signal output
rlabel metal2 s 65982 199200 66038 200000 6 slave2_wb_data_i[29]
port 572 nsew signal output
rlabel metal2 s 10966 199200 11022 200000 6 slave2_wb_data_i[2]
port 573 nsew signal output
rlabel metal2 s 67362 199200 67418 200000 6 slave2_wb_data_i[30]
port 574 nsew signal output
rlabel metal2 s 68834 199200 68890 200000 6 slave2_wb_data_i[31]
port 575 nsew signal output
rlabel metal2 s 13818 199200 13874 200000 6 slave2_wb_data_i[3]
port 576 nsew signal output
rlabel metal2 s 16670 199200 16726 200000 6 slave2_wb_data_i[4]
port 577 nsew signal output
rlabel metal2 s 18786 199200 18842 200000 6 slave2_wb_data_i[5]
port 578 nsew signal output
rlabel metal2 s 20994 199200 21050 200000 6 slave2_wb_data_i[6]
port 579 nsew signal output
rlabel metal2 s 23110 199200 23166 200000 6 slave2_wb_data_i[7]
port 580 nsew signal output
rlabel metal2 s 25226 199200 25282 200000 6 slave2_wb_data_i[8]
port 581 nsew signal output
rlabel metal2 s 27434 199200 27490 200000 6 slave2_wb_data_i[9]
port 582 nsew signal output
rlabel metal2 s 5998 199200 6054 200000 6 slave2_wb_data_o[0]
port 583 nsew signal input
rlabel metal2 s 30286 199200 30342 200000 6 slave2_wb_data_o[10]
port 584 nsew signal input
rlabel metal2 s 32402 199200 32458 200000 6 slave2_wb_data_o[11]
port 585 nsew signal input
rlabel metal2 s 34518 199200 34574 200000 6 slave2_wb_data_o[12]
port 586 nsew signal input
rlabel metal2 s 36726 199200 36782 200000 6 slave2_wb_data_o[13]
port 587 nsew signal input
rlabel metal2 s 38842 199200 38898 200000 6 slave2_wb_data_o[14]
port 588 nsew signal input
rlabel metal2 s 40958 199200 41014 200000 6 slave2_wb_data_o[15]
port 589 nsew signal input
rlabel metal2 s 43074 199200 43130 200000 6 slave2_wb_data_o[16]
port 590 nsew signal input
rlabel metal2 s 45282 199200 45338 200000 6 slave2_wb_data_o[17]
port 591 nsew signal input
rlabel metal2 s 47398 199200 47454 200000 6 slave2_wb_data_o[18]
port 592 nsew signal input
rlabel metal2 s 49514 199200 49570 200000 6 slave2_wb_data_o[19]
port 593 nsew signal input
rlabel metal2 s 8850 199200 8906 200000 6 slave2_wb_data_o[1]
port 594 nsew signal input
rlabel metal2 s 51722 199200 51778 200000 6 slave2_wb_data_o[20]
port 595 nsew signal input
rlabel metal2 s 53838 199200 53894 200000 6 slave2_wb_data_o[21]
port 596 nsew signal input
rlabel metal2 s 55954 199200 56010 200000 6 slave2_wb_data_o[22]
port 597 nsew signal input
rlabel metal2 s 58070 199200 58126 200000 6 slave2_wb_data_o[23]
port 598 nsew signal input
rlabel metal2 s 59542 199200 59598 200000 6 slave2_wb_data_o[24]
port 599 nsew signal input
rlabel metal2 s 61014 199200 61070 200000 6 slave2_wb_data_o[25]
port 600 nsew signal input
rlabel metal2 s 62394 199200 62450 200000 6 slave2_wb_data_o[26]
port 601 nsew signal input
rlabel metal2 s 63866 199200 63922 200000 6 slave2_wb_data_o[27]
port 602 nsew signal input
rlabel metal2 s 65246 199200 65302 200000 6 slave2_wb_data_o[28]
port 603 nsew signal input
rlabel metal2 s 66718 199200 66774 200000 6 slave2_wb_data_o[29]
port 604 nsew signal input
rlabel metal2 s 11702 199200 11758 200000 6 slave2_wb_data_o[2]
port 605 nsew signal input
rlabel metal2 s 68098 199200 68154 200000 6 slave2_wb_data_o[30]
port 606 nsew signal input
rlabel metal2 s 69570 199200 69626 200000 6 slave2_wb_data_o[31]
port 607 nsew signal input
rlabel metal2 s 14554 199200 14610 200000 6 slave2_wb_data_o[3]
port 608 nsew signal input
rlabel metal2 s 17406 199200 17462 200000 6 slave2_wb_data_o[4]
port 609 nsew signal input
rlabel metal2 s 19522 199200 19578 200000 6 slave2_wb_data_o[5]
port 610 nsew signal input
rlabel metal2 s 21638 199200 21694 200000 6 slave2_wb_data_o[6]
port 611 nsew signal input
rlabel metal2 s 23846 199200 23902 200000 6 slave2_wb_data_o[7]
port 612 nsew signal input
rlabel metal2 s 25962 199200 26018 200000 6 slave2_wb_data_o[8]
port 613 nsew signal input
rlabel metal2 s 28078 199200 28134 200000 6 slave2_wb_data_o[9]
port 614 nsew signal input
rlabel metal2 s 1674 199200 1730 200000 6 slave2_wb_error_o
port 615 nsew signal input
rlabel metal2 s 6642 199200 6698 200000 6 slave2_wb_sel_i[0]
port 616 nsew signal output
rlabel metal2 s 9494 199200 9550 200000 6 slave2_wb_sel_i[1]
port 617 nsew signal output
rlabel metal2 s 12438 199200 12494 200000 6 slave2_wb_sel_i[2]
port 618 nsew signal output
rlabel metal2 s 15290 199200 15346 200000 6 slave2_wb_sel_i[3]
port 619 nsew signal output
rlabel metal2 s 2410 199200 2466 200000 6 slave2_wb_stall_o
port 620 nsew signal input
rlabel metal2 s 3146 199200 3202 200000 6 slave2_wb_stb_i
port 621 nsew signal output
rlabel metal2 s 3790 199200 3846 200000 6 slave2_wb_we_i
port 622 nsew signal output
rlabel metal3 s 69200 100376 70000 100496 6 slave3_wb_ack_o
port 623 nsew signal input
rlabel metal3 s 69200 106496 70000 106616 6 slave3_wb_adr_i[0]
port 624 nsew signal output
rlabel metal3 s 69200 141176 70000 141296 6 slave3_wb_adr_i[10]
port 625 nsew signal output
rlabel metal3 s 69200 144304 70000 144424 6 slave3_wb_adr_i[11]
port 626 nsew signal output
rlabel metal3 s 69200 147296 70000 147416 6 slave3_wb_adr_i[12]
port 627 nsew signal output
rlabel metal3 s 69200 150424 70000 150544 6 slave3_wb_adr_i[13]
port 628 nsew signal output
rlabel metal3 s 69200 153416 70000 153536 6 slave3_wb_adr_i[14]
port 629 nsew signal output
rlabel metal3 s 69200 156544 70000 156664 6 slave3_wb_adr_i[15]
port 630 nsew signal output
rlabel metal3 s 69200 159536 70000 159656 6 slave3_wb_adr_i[16]
port 631 nsew signal output
rlabel metal3 s 69200 162664 70000 162784 6 slave3_wb_adr_i[17]
port 632 nsew signal output
rlabel metal3 s 69200 165656 70000 165776 6 slave3_wb_adr_i[18]
port 633 nsew signal output
rlabel metal3 s 69200 168784 70000 168904 6 slave3_wb_adr_i[19]
port 634 nsew signal output
rlabel metal3 s 69200 110576 70000 110696 6 slave3_wb_adr_i[1]
port 635 nsew signal output
rlabel metal3 s 69200 171776 70000 171896 6 slave3_wb_adr_i[20]
port 636 nsew signal output
rlabel metal3 s 69200 174904 70000 175024 6 slave3_wb_adr_i[21]
port 637 nsew signal output
rlabel metal3 s 69200 177896 70000 178016 6 slave3_wb_adr_i[22]
port 638 nsew signal output
rlabel metal3 s 69200 181024 70000 181144 6 slave3_wb_adr_i[23]
port 639 nsew signal output
rlabel metal3 s 69200 114656 70000 114776 6 slave3_wb_adr_i[2]
port 640 nsew signal output
rlabel metal3 s 69200 118736 70000 118856 6 slave3_wb_adr_i[3]
port 641 nsew signal output
rlabel metal3 s 69200 122816 70000 122936 6 slave3_wb_adr_i[4]
port 642 nsew signal output
rlabel metal3 s 69200 125944 70000 126064 6 slave3_wb_adr_i[5]
port 643 nsew signal output
rlabel metal3 s 69200 128936 70000 129056 6 slave3_wb_adr_i[6]
port 644 nsew signal output
rlabel metal3 s 69200 132064 70000 132184 6 slave3_wb_adr_i[7]
port 645 nsew signal output
rlabel metal3 s 69200 135056 70000 135176 6 slave3_wb_adr_i[8]
port 646 nsew signal output
rlabel metal3 s 69200 138184 70000 138304 6 slave3_wb_adr_i[9]
port 647 nsew signal output
rlabel metal3 s 69200 101464 70000 101584 6 slave3_wb_cyc_i
port 648 nsew signal output
rlabel metal3 s 69200 107584 70000 107704 6 slave3_wb_data_i[0]
port 649 nsew signal output
rlabel metal3 s 69200 142264 70000 142384 6 slave3_wb_data_i[10]
port 650 nsew signal output
rlabel metal3 s 69200 145256 70000 145376 6 slave3_wb_data_i[11]
port 651 nsew signal output
rlabel metal3 s 69200 148384 70000 148504 6 slave3_wb_data_i[12]
port 652 nsew signal output
rlabel metal3 s 69200 151376 70000 151496 6 slave3_wb_data_i[13]
port 653 nsew signal output
rlabel metal3 s 69200 154504 70000 154624 6 slave3_wb_data_i[14]
port 654 nsew signal output
rlabel metal3 s 69200 157496 70000 157616 6 slave3_wb_data_i[15]
port 655 nsew signal output
rlabel metal3 s 69200 160624 70000 160744 6 slave3_wb_data_i[16]
port 656 nsew signal output
rlabel metal3 s 69200 163616 70000 163736 6 slave3_wb_data_i[17]
port 657 nsew signal output
rlabel metal3 s 69200 166744 70000 166864 6 slave3_wb_data_i[18]
port 658 nsew signal output
rlabel metal3 s 69200 169736 70000 169856 6 slave3_wb_data_i[19]
port 659 nsew signal output
rlabel metal3 s 69200 111664 70000 111784 6 slave3_wb_data_i[1]
port 660 nsew signal output
rlabel metal3 s 69200 172864 70000 172984 6 slave3_wb_data_i[20]
port 661 nsew signal output
rlabel metal3 s 69200 175856 70000 175976 6 slave3_wb_data_i[21]
port 662 nsew signal output
rlabel metal3 s 69200 178984 70000 179104 6 slave3_wb_data_i[22]
port 663 nsew signal output
rlabel metal3 s 69200 181976 70000 182096 6 slave3_wb_data_i[23]
port 664 nsew signal output
rlabel metal3 s 69200 184016 70000 184136 6 slave3_wb_data_i[24]
port 665 nsew signal output
rlabel metal3 s 69200 186056 70000 186176 6 slave3_wb_data_i[25]
port 666 nsew signal output
rlabel metal3 s 69200 188096 70000 188216 6 slave3_wb_data_i[26]
port 667 nsew signal output
rlabel metal3 s 69200 190136 70000 190256 6 slave3_wb_data_i[27]
port 668 nsew signal output
rlabel metal3 s 69200 192176 70000 192296 6 slave3_wb_data_i[28]
port 669 nsew signal output
rlabel metal3 s 69200 194216 70000 194336 6 slave3_wb_data_i[29]
port 670 nsew signal output
rlabel metal3 s 69200 115744 70000 115864 6 slave3_wb_data_i[2]
port 671 nsew signal output
rlabel metal3 s 69200 196256 70000 196376 6 slave3_wb_data_i[30]
port 672 nsew signal output
rlabel metal3 s 69200 198296 70000 198416 6 slave3_wb_data_i[31]
port 673 nsew signal output
rlabel metal3 s 69200 119824 70000 119944 6 slave3_wb_data_i[3]
port 674 nsew signal output
rlabel metal3 s 69200 123904 70000 124024 6 slave3_wb_data_i[4]
port 675 nsew signal output
rlabel metal3 s 69200 126896 70000 127016 6 slave3_wb_data_i[5]
port 676 nsew signal output
rlabel metal3 s 69200 130024 70000 130144 6 slave3_wb_data_i[6]
port 677 nsew signal output
rlabel metal3 s 69200 133016 70000 133136 6 slave3_wb_data_i[7]
port 678 nsew signal output
rlabel metal3 s 69200 136144 70000 136264 6 slave3_wb_data_i[8]
port 679 nsew signal output
rlabel metal3 s 69200 139136 70000 139256 6 slave3_wb_data_i[9]
port 680 nsew signal output
rlabel metal3 s 69200 108536 70000 108656 6 slave3_wb_data_o[0]
port 681 nsew signal input
rlabel metal3 s 69200 143216 70000 143336 6 slave3_wb_data_o[10]
port 682 nsew signal input
rlabel metal3 s 69200 146344 70000 146464 6 slave3_wb_data_o[11]
port 683 nsew signal input
rlabel metal3 s 69200 149336 70000 149456 6 slave3_wb_data_o[12]
port 684 nsew signal input
rlabel metal3 s 69200 152464 70000 152584 6 slave3_wb_data_o[13]
port 685 nsew signal input
rlabel metal3 s 69200 155456 70000 155576 6 slave3_wb_data_o[14]
port 686 nsew signal input
rlabel metal3 s 69200 158584 70000 158704 6 slave3_wb_data_o[15]
port 687 nsew signal input
rlabel metal3 s 69200 161576 70000 161696 6 slave3_wb_data_o[16]
port 688 nsew signal input
rlabel metal3 s 69200 164704 70000 164824 6 slave3_wb_data_o[17]
port 689 nsew signal input
rlabel metal3 s 69200 167696 70000 167816 6 slave3_wb_data_o[18]
port 690 nsew signal input
rlabel metal3 s 69200 170824 70000 170944 6 slave3_wb_data_o[19]
port 691 nsew signal input
rlabel metal3 s 69200 112616 70000 112736 6 slave3_wb_data_o[1]
port 692 nsew signal input
rlabel metal3 s 69200 173816 70000 173936 6 slave3_wb_data_o[20]
port 693 nsew signal input
rlabel metal3 s 69200 176944 70000 177064 6 slave3_wb_data_o[21]
port 694 nsew signal input
rlabel metal3 s 69200 179936 70000 180056 6 slave3_wb_data_o[22]
port 695 nsew signal input
rlabel metal3 s 69200 183064 70000 183184 6 slave3_wb_data_o[23]
port 696 nsew signal input
rlabel metal3 s 69200 185104 70000 185224 6 slave3_wb_data_o[24]
port 697 nsew signal input
rlabel metal3 s 69200 187144 70000 187264 6 slave3_wb_data_o[25]
port 698 nsew signal input
rlabel metal3 s 69200 189184 70000 189304 6 slave3_wb_data_o[26]
port 699 nsew signal input
rlabel metal3 s 69200 191224 70000 191344 6 slave3_wb_data_o[27]
port 700 nsew signal input
rlabel metal3 s 69200 193264 70000 193384 6 slave3_wb_data_o[28]
port 701 nsew signal input
rlabel metal3 s 69200 195304 70000 195424 6 slave3_wb_data_o[29]
port 702 nsew signal input
rlabel metal3 s 69200 116696 70000 116816 6 slave3_wb_data_o[2]
port 703 nsew signal input
rlabel metal3 s 69200 197344 70000 197464 6 slave3_wb_data_o[30]
port 704 nsew signal input
rlabel metal3 s 69200 199384 70000 199504 6 slave3_wb_data_o[31]
port 705 nsew signal input
rlabel metal3 s 69200 120776 70000 120896 6 slave3_wb_data_o[3]
port 706 nsew signal input
rlabel metal3 s 69200 124856 70000 124976 6 slave3_wb_data_o[4]
port 707 nsew signal input
rlabel metal3 s 69200 127984 70000 128104 6 slave3_wb_data_o[5]
port 708 nsew signal input
rlabel metal3 s 69200 130976 70000 131096 6 slave3_wb_data_o[6]
port 709 nsew signal input
rlabel metal3 s 69200 134104 70000 134224 6 slave3_wb_data_o[7]
port 710 nsew signal input
rlabel metal3 s 69200 137096 70000 137216 6 slave3_wb_data_o[8]
port 711 nsew signal input
rlabel metal3 s 69200 140224 70000 140344 6 slave3_wb_data_o[9]
port 712 nsew signal input
rlabel metal3 s 69200 102416 70000 102536 6 slave3_wb_error_o
port 713 nsew signal input
rlabel metal3 s 69200 109624 70000 109744 6 slave3_wb_sel_i[0]
port 714 nsew signal output
rlabel metal3 s 69200 113704 70000 113824 6 slave3_wb_sel_i[1]
port 715 nsew signal output
rlabel metal3 s 69200 117784 70000 117904 6 slave3_wb_sel_i[2]
port 716 nsew signal output
rlabel metal3 s 69200 121864 70000 121984 6 slave3_wb_sel_i[3]
port 717 nsew signal output
rlabel metal3 s 69200 103504 70000 103624 6 slave3_wb_stall_o
port 718 nsew signal input
rlabel metal3 s 69200 104456 70000 104576 6 slave3_wb_stb_i
port 719 nsew signal output
rlabel metal3 s 69200 105544 70000 105664 6 slave3_wb_we_i
port 720 nsew signal output
rlabel metal3 s 69200 416 70000 536 6 slave4_wb_ack_o
port 721 nsew signal input
rlabel metal3 s 69200 6536 70000 6656 6 slave4_wb_adr_i[0]
port 722 nsew signal output
rlabel metal3 s 69200 41216 70000 41336 6 slave4_wb_adr_i[10]
port 723 nsew signal output
rlabel metal3 s 69200 44208 70000 44328 6 slave4_wb_adr_i[11]
port 724 nsew signal output
rlabel metal3 s 69200 47336 70000 47456 6 slave4_wb_adr_i[12]
port 725 nsew signal output
rlabel metal3 s 69200 50328 70000 50448 6 slave4_wb_adr_i[13]
port 726 nsew signal output
rlabel metal3 s 69200 53456 70000 53576 6 slave4_wb_adr_i[14]
port 727 nsew signal output
rlabel metal3 s 69200 56448 70000 56568 6 slave4_wb_adr_i[15]
port 728 nsew signal output
rlabel metal3 s 69200 59576 70000 59696 6 slave4_wb_adr_i[16]
port 729 nsew signal output
rlabel metal3 s 69200 62568 70000 62688 6 slave4_wb_adr_i[17]
port 730 nsew signal output
rlabel metal3 s 69200 65696 70000 65816 6 slave4_wb_adr_i[18]
port 731 nsew signal output
rlabel metal3 s 69200 68688 70000 68808 6 slave4_wb_adr_i[19]
port 732 nsew signal output
rlabel metal3 s 69200 10616 70000 10736 6 slave4_wb_adr_i[1]
port 733 nsew signal output
rlabel metal3 s 69200 71816 70000 71936 6 slave4_wb_adr_i[20]
port 734 nsew signal output
rlabel metal3 s 69200 74808 70000 74928 6 slave4_wb_adr_i[21]
port 735 nsew signal output
rlabel metal3 s 69200 77936 70000 78056 6 slave4_wb_adr_i[22]
port 736 nsew signal output
rlabel metal3 s 69200 80928 70000 81048 6 slave4_wb_adr_i[23]
port 737 nsew signal output
rlabel metal3 s 69200 14696 70000 14816 6 slave4_wb_adr_i[2]
port 738 nsew signal output
rlabel metal3 s 69200 18776 70000 18896 6 slave4_wb_adr_i[3]
port 739 nsew signal output
rlabel metal3 s 69200 22856 70000 22976 6 slave4_wb_adr_i[4]
port 740 nsew signal output
rlabel metal3 s 69200 25848 70000 25968 6 slave4_wb_adr_i[5]
port 741 nsew signal output
rlabel metal3 s 69200 28976 70000 29096 6 slave4_wb_adr_i[6]
port 742 nsew signal output
rlabel metal3 s 69200 31968 70000 32088 6 slave4_wb_adr_i[7]
port 743 nsew signal output
rlabel metal3 s 69200 35096 70000 35216 6 slave4_wb_adr_i[8]
port 744 nsew signal output
rlabel metal3 s 69200 38088 70000 38208 6 slave4_wb_adr_i[9]
port 745 nsew signal output
rlabel metal3 s 69200 1368 70000 1488 6 slave4_wb_cyc_i
port 746 nsew signal output
rlabel metal3 s 69200 7488 70000 7608 6 slave4_wb_data_i[0]
port 747 nsew signal output
rlabel metal3 s 69200 42168 70000 42288 6 slave4_wb_data_i[10]
port 748 nsew signal output
rlabel metal3 s 69200 45296 70000 45416 6 slave4_wb_data_i[11]
port 749 nsew signal output
rlabel metal3 s 69200 48288 70000 48408 6 slave4_wb_data_i[12]
port 750 nsew signal output
rlabel metal3 s 69200 51416 70000 51536 6 slave4_wb_data_i[13]
port 751 nsew signal output
rlabel metal3 s 69200 54408 70000 54528 6 slave4_wb_data_i[14]
port 752 nsew signal output
rlabel metal3 s 69200 57536 70000 57656 6 slave4_wb_data_i[15]
port 753 nsew signal output
rlabel metal3 s 69200 60528 70000 60648 6 slave4_wb_data_i[16]
port 754 nsew signal output
rlabel metal3 s 69200 63656 70000 63776 6 slave4_wb_data_i[17]
port 755 nsew signal output
rlabel metal3 s 69200 66648 70000 66768 6 slave4_wb_data_i[18]
port 756 nsew signal output
rlabel metal3 s 69200 69776 70000 69896 6 slave4_wb_data_i[19]
port 757 nsew signal output
rlabel metal3 s 69200 11568 70000 11688 6 slave4_wb_data_i[1]
port 758 nsew signal output
rlabel metal3 s 69200 72768 70000 72888 6 slave4_wb_data_i[20]
port 759 nsew signal output
rlabel metal3 s 69200 75896 70000 76016 6 slave4_wb_data_i[21]
port 760 nsew signal output
rlabel metal3 s 69200 78888 70000 79008 6 slave4_wb_data_i[22]
port 761 nsew signal output
rlabel metal3 s 69200 82016 70000 82136 6 slave4_wb_data_i[23]
port 762 nsew signal output
rlabel metal3 s 69200 84056 70000 84176 6 slave4_wb_data_i[24]
port 763 nsew signal output
rlabel metal3 s 69200 86096 70000 86216 6 slave4_wb_data_i[25]
port 764 nsew signal output
rlabel metal3 s 69200 88136 70000 88256 6 slave4_wb_data_i[26]
port 765 nsew signal output
rlabel metal3 s 69200 90176 70000 90296 6 slave4_wb_data_i[27]
port 766 nsew signal output
rlabel metal3 s 69200 92216 70000 92336 6 slave4_wb_data_i[28]
port 767 nsew signal output
rlabel metal3 s 69200 94256 70000 94376 6 slave4_wb_data_i[29]
port 768 nsew signal output
rlabel metal3 s 69200 15648 70000 15768 6 slave4_wb_data_i[2]
port 769 nsew signal output
rlabel metal3 s 69200 96296 70000 96416 6 slave4_wb_data_i[30]
port 770 nsew signal output
rlabel metal3 s 69200 98336 70000 98456 6 slave4_wb_data_i[31]
port 771 nsew signal output
rlabel metal3 s 69200 19728 70000 19848 6 slave4_wb_data_i[3]
port 772 nsew signal output
rlabel metal3 s 69200 23808 70000 23928 6 slave4_wb_data_i[4]
port 773 nsew signal output
rlabel metal3 s 69200 26936 70000 27056 6 slave4_wb_data_i[5]
port 774 nsew signal output
rlabel metal3 s 69200 29928 70000 30048 6 slave4_wb_data_i[6]
port 775 nsew signal output
rlabel metal3 s 69200 33056 70000 33176 6 slave4_wb_data_i[7]
port 776 nsew signal output
rlabel metal3 s 69200 36048 70000 36168 6 slave4_wb_data_i[8]
port 777 nsew signal output
rlabel metal3 s 69200 39176 70000 39296 6 slave4_wb_data_i[9]
port 778 nsew signal output
rlabel metal3 s 69200 8576 70000 8696 6 slave4_wb_data_o[0]
port 779 nsew signal input
rlabel metal3 s 69200 43256 70000 43376 6 slave4_wb_data_o[10]
port 780 nsew signal input
rlabel metal3 s 69200 46248 70000 46368 6 slave4_wb_data_o[11]
port 781 nsew signal input
rlabel metal3 s 69200 49376 70000 49496 6 slave4_wb_data_o[12]
port 782 nsew signal input
rlabel metal3 s 69200 52368 70000 52488 6 slave4_wb_data_o[13]
port 783 nsew signal input
rlabel metal3 s 69200 55496 70000 55616 6 slave4_wb_data_o[14]
port 784 nsew signal input
rlabel metal3 s 69200 58488 70000 58608 6 slave4_wb_data_o[15]
port 785 nsew signal input
rlabel metal3 s 69200 61616 70000 61736 6 slave4_wb_data_o[16]
port 786 nsew signal input
rlabel metal3 s 69200 64608 70000 64728 6 slave4_wb_data_o[17]
port 787 nsew signal input
rlabel metal3 s 69200 67736 70000 67856 6 slave4_wb_data_o[18]
port 788 nsew signal input
rlabel metal3 s 69200 70728 70000 70848 6 slave4_wb_data_o[19]
port 789 nsew signal input
rlabel metal3 s 69200 12656 70000 12776 6 slave4_wb_data_o[1]
port 790 nsew signal input
rlabel metal3 s 69200 73856 70000 73976 6 slave4_wb_data_o[20]
port 791 nsew signal input
rlabel metal3 s 69200 76848 70000 76968 6 slave4_wb_data_o[21]
port 792 nsew signal input
rlabel metal3 s 69200 79976 70000 80096 6 slave4_wb_data_o[22]
port 793 nsew signal input
rlabel metal3 s 69200 82968 70000 83088 6 slave4_wb_data_o[23]
port 794 nsew signal input
rlabel metal3 s 69200 85008 70000 85128 6 slave4_wb_data_o[24]
port 795 nsew signal input
rlabel metal3 s 69200 87048 70000 87168 6 slave4_wb_data_o[25]
port 796 nsew signal input
rlabel metal3 s 69200 89088 70000 89208 6 slave4_wb_data_o[26]
port 797 nsew signal input
rlabel metal3 s 69200 91128 70000 91248 6 slave4_wb_data_o[27]
port 798 nsew signal input
rlabel metal3 s 69200 93168 70000 93288 6 slave4_wb_data_o[28]
port 799 nsew signal input
rlabel metal3 s 69200 95208 70000 95328 6 slave4_wb_data_o[29]
port 800 nsew signal input
rlabel metal3 s 69200 16736 70000 16856 6 slave4_wb_data_o[2]
port 801 nsew signal input
rlabel metal3 s 69200 97248 70000 97368 6 slave4_wb_data_o[30]
port 802 nsew signal input
rlabel metal3 s 69200 99288 70000 99408 6 slave4_wb_data_o[31]
port 803 nsew signal input
rlabel metal3 s 69200 20816 70000 20936 6 slave4_wb_data_o[3]
port 804 nsew signal input
rlabel metal3 s 69200 24896 70000 25016 6 slave4_wb_data_o[4]
port 805 nsew signal input
rlabel metal3 s 69200 27888 70000 28008 6 slave4_wb_data_o[5]
port 806 nsew signal input
rlabel metal3 s 69200 31016 70000 31136 6 slave4_wb_data_o[6]
port 807 nsew signal input
rlabel metal3 s 69200 34008 70000 34128 6 slave4_wb_data_o[7]
port 808 nsew signal input
rlabel metal3 s 69200 37136 70000 37256 6 slave4_wb_data_o[8]
port 809 nsew signal input
rlabel metal3 s 69200 40128 70000 40248 6 slave4_wb_data_o[9]
port 810 nsew signal input
rlabel metal3 s 69200 2456 70000 2576 6 slave4_wb_error_o
port 811 nsew signal input
rlabel metal3 s 69200 9528 70000 9648 6 slave4_wb_sel_i[0]
port 812 nsew signal output
rlabel metal3 s 69200 13608 70000 13728 6 slave4_wb_sel_i[1]
port 813 nsew signal output
rlabel metal3 s 69200 17688 70000 17808 6 slave4_wb_sel_i[2]
port 814 nsew signal output
rlabel metal3 s 69200 21768 70000 21888 6 slave4_wb_sel_i[3]
port 815 nsew signal output
rlabel metal3 s 69200 3408 70000 3528 6 slave4_wb_stall_o
port 816 nsew signal input
rlabel metal3 s 69200 4496 70000 4616 6 slave4_wb_stb_i
port 817 nsew signal output
rlabel metal3 s 69200 5448 70000 5568 6 slave4_wb_we_i
port 818 nsew signal output
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 819 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 819 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 819 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 820 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 820 nsew ground bidirectional
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 821 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 822 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12571144
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/WishboneInterconnect/runs/WishboneInterconnect/results/signoff/WishboneInterconnect.magic.gds
string GDS_START 600892
<< end >>

