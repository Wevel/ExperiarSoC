VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Peripherals
  CLASS BLOCK ;
  FOREIGN Peripherals ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 950.000 ;
  PIN flash_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END flash_csb
  PIN flash_io0_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END flash_io0_read
  PIN flash_io0_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END flash_io0_we
  PIN flash_io0_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END flash_io0_write
  PIN flash_io1_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END flash_io1_read
  PIN flash_io1_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END flash_io1_we
  PIN flash_io1_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END flash_io1_write
  PIN flash_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END flash_sck
  PIN internal_uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END internal_uart_rx
  PIN internal_uart_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END internal_uart_tx
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 946.000 6.810 950.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 946.000 85.010 950.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 946.000 92.830 950.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 946.000 100.650 950.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 946.000 108.470 950.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 946.000 116.290 950.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 946.000 124.110 950.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 946.000 131.930 950.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 946.000 139.750 950.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 946.000 147.570 950.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 946.000 155.390 950.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 946.000 14.630 950.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 946.000 163.210 950.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 946.000 171.030 950.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 946.000 178.850 950.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 946.000 186.670 950.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 946.000 194.490 950.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 946.000 202.310 950.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 946.000 210.130 950.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 946.000 217.950 950.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 946.000 225.770 950.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 946.000 233.590 950.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 946.000 22.450 950.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 946.000 241.410 950.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 946.000 249.230 950.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 946.000 257.050 950.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 946.000 264.870 950.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 946.000 272.690 950.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 946.000 280.510 950.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 946.000 288.330 950.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 946.000 296.150 950.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 946.000 30.270 950.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 946.000 38.090 950.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 946.000 45.910 950.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 946.000 53.730 950.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 946.000 61.550 950.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 946.000 69.370 950.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 946.000 77.190 950.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 946.000 303.970 950.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 946.000 382.170 950.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 946.000 389.990 950.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 946.000 397.810 950.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 946.000 405.630 950.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 946.000 413.450 950.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 946.000 421.270 950.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 946.000 429.090 950.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 946.000 436.910 950.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 946.000 444.730 950.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 946.000 452.550 950.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 946.000 311.790 950.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 946.000 460.370 950.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 946.000 468.190 950.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 946.000 476.010 950.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 946.000 483.830 950.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 946.000 491.650 950.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 946.000 499.470 950.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 946.000 507.290 950.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 946.000 515.110 950.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 946.000 522.930 950.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 946.000 530.750 950.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 946.000 319.610 950.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 946.000 538.570 950.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 946.000 546.390 950.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 946.000 554.210 950.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 946.000 562.030 950.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 946.000 569.850 950.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 946.000 577.670 950.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 946.000 585.490 950.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 946.000 593.310 950.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 946.000 327.430 950.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 946.000 335.250 950.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 946.000 343.070 950.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 946.000 350.890 950.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 946.000 358.710 950.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 946.000 366.530 950.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 946.000 374.350 950.000 ;
    END
  END io_out[9]
  PIN jtag_tck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 395.800 600.000 396.400 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 553.560 600.000 554.160 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 711.320 600.000 711.920 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 869.080 600.000 869.680 ;
    END
  END jtag_tms
  PIN peripheral_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END peripheral_irq[0]
  PIN peripheral_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END peripheral_irq[1]
  PIN peripheral_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END peripheral_irq[2]
  PIN peripheral_irq[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END peripheral_irq[3]
  PIN peripheral_irq[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END peripheral_irq[4]
  PIN peripheral_irq[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END peripheral_irq[5]
  PIN peripheral_irq[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END peripheral_irq[6]
  PIN peripheral_irq[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END peripheral_irq[7]
  PIN peripheral_irq[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END peripheral_irq[8]
  PIN peripheral_irq[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END peripheral_irq[9]
  PIN probe_blink[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 80.280 600.000 80.880 ;
    END
  END probe_blink[0]
  PIN probe_blink[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 238.040 600.000 238.640 ;
    END
  END probe_blink[1]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 938.640 ;
    END
  END vccd1
  PIN vga_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END vga_b[0]
  PIN vga_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END vga_b[1]
  PIN vga_g[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 0.000 549.150 4.000 ;
    END
  END vga_g[0]
  PIN vga_g[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END vga_g[1]
  PIN vga_hsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END vga_hsync
  PIN vga_r[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END vga_r[0]
  PIN vga_r[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END vga_r[1]
  PIN vga_vsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END vga_vsync
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 938.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 938.640 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 434.560 4.000 435.160 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 487.600 4.000 488.200 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.680 4.000 594.280 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.760 4.000 700.360 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.280 4.000 726.880 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.800 4.000 753.400 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END wb_cyc_i
  PIN wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END wb_data_i[0]
  PIN wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.880 4.000 417.480 ;
    END
  END wb_data_i[10]
  PIN wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END wb_data_i[11]
  PIN wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.920 4.000 470.520 ;
    END
  END wb_data_i[12]
  PIN wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END wb_data_i[13]
  PIN wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.960 4.000 523.560 ;
    END
  END wb_data_i[14]
  PIN wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END wb_data_i[15]
  PIN wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.000 4.000 576.600 ;
    END
  END wb_data_i[16]
  PIN wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END wb_data_i[17]
  PIN wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END wb_data_i[18]
  PIN wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END wb_data_i[19]
  PIN wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END wb_data_i[1]
  PIN wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.080 4.000 682.680 ;
    END
  END wb_data_i[20]
  PIN wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 4.000 709.200 ;
    END
  END wb_data_i[21]
  PIN wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.120 4.000 735.720 ;
    END
  END wb_data_i[22]
  PIN wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END wb_data_i[23]
  PIN wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 4.000 779.920 ;
    END
  END wb_data_i[24]
  PIN wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END wb_data_i[25]
  PIN wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.680 4.000 815.280 ;
    END
  END wb_data_i[26]
  PIN wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END wb_data_i[27]
  PIN wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END wb_data_i[28]
  PIN wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.720 4.000 868.320 ;
    END
  END wb_data_i[29]
  PIN wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END wb_data_i[2]
  PIN wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 885.400 4.000 886.000 ;
    END
  END wb_data_i[30]
  PIN wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 903.080 4.000 903.680 ;
    END
  END wb_data_i[31]
  PIN wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END wb_data_i[3]
  PIN wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END wb_data_i[4]
  PIN wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END wb_data_i[5]
  PIN wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END wb_data_i[6]
  PIN wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END wb_data_i[7]
  PIN wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END wb_data_i[8]
  PIN wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END wb_data_i[9]
  PIN wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END wb_data_o[0]
  PIN wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END wb_data_o[10]
  PIN wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END wb_data_o[11]
  PIN wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END wb_data_o[12]
  PIN wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.280 4.000 505.880 ;
    END
  END wb_data_o[13]
  PIN wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END wb_data_o[14]
  PIN wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 558.320 4.000 558.920 ;
    END
  END wb_data_o[15]
  PIN wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END wb_data_o[16]
  PIN wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 611.360 4.000 611.960 ;
    END
  END wb_data_o[17]
  PIN wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END wb_data_o[18]
  PIN wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 664.400 4.000 665.000 ;
    END
  END wb_data_o[19]
  PIN wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END wb_data_o[1]
  PIN wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END wb_data_o[20]
  PIN wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END wb_data_o[21]
  PIN wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END wb_data_o[22]
  PIN wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 770.480 4.000 771.080 ;
    END
  END wb_data_o[23]
  PIN wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.160 4.000 788.760 ;
    END
  END wb_data_o[24]
  PIN wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END wb_data_o[25]
  PIN wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 823.520 4.000 824.120 ;
    END
  END wb_data_o[26]
  PIN wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 841.200 4.000 841.800 ;
    END
  END wb_data_o[27]
  PIN wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 858.880 4.000 859.480 ;
    END
  END wb_data_o[28]
  PIN wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 876.560 4.000 877.160 ;
    END
  END wb_data_o[29]
  PIN wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END wb_data_o[2]
  PIN wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END wb_data_o[30]
  PIN wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.920 4.000 912.520 ;
    END
  END wb_data_o[31]
  PIN wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END wb_data_o[3]
  PIN wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END wb_data_o[4]
  PIN wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END wb_data_o[5]
  PIN wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END wb_data_o[6]
  PIN wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END wb_data_o[7]
  PIN wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END wb_data_o[8]
  PIN wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.200 4.000 399.800 ;
    END
  END wb_data_o[9]
  PIN wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END wb_error_o
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.360 4.000 169.960 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END wb_sel_i[3]
  PIN wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END wb_stall_o
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 938.485 ;
      LAYER met1 ;
        RECT 4.670 4.460 595.630 945.500 ;
      LAYER met2 ;
        RECT 4.690 945.720 6.250 946.000 ;
        RECT 7.090 945.720 14.070 946.000 ;
        RECT 14.910 945.720 21.890 946.000 ;
        RECT 22.730 945.720 29.710 946.000 ;
        RECT 30.550 945.720 37.530 946.000 ;
        RECT 38.370 945.720 45.350 946.000 ;
        RECT 46.190 945.720 53.170 946.000 ;
        RECT 54.010 945.720 60.990 946.000 ;
        RECT 61.830 945.720 68.810 946.000 ;
        RECT 69.650 945.720 76.630 946.000 ;
        RECT 77.470 945.720 84.450 946.000 ;
        RECT 85.290 945.720 92.270 946.000 ;
        RECT 93.110 945.720 100.090 946.000 ;
        RECT 100.930 945.720 107.910 946.000 ;
        RECT 108.750 945.720 115.730 946.000 ;
        RECT 116.570 945.720 123.550 946.000 ;
        RECT 124.390 945.720 131.370 946.000 ;
        RECT 132.210 945.720 139.190 946.000 ;
        RECT 140.030 945.720 147.010 946.000 ;
        RECT 147.850 945.720 154.830 946.000 ;
        RECT 155.670 945.720 162.650 946.000 ;
        RECT 163.490 945.720 170.470 946.000 ;
        RECT 171.310 945.720 178.290 946.000 ;
        RECT 179.130 945.720 186.110 946.000 ;
        RECT 186.950 945.720 193.930 946.000 ;
        RECT 194.770 945.720 201.750 946.000 ;
        RECT 202.590 945.720 209.570 946.000 ;
        RECT 210.410 945.720 217.390 946.000 ;
        RECT 218.230 945.720 225.210 946.000 ;
        RECT 226.050 945.720 233.030 946.000 ;
        RECT 233.870 945.720 240.850 946.000 ;
        RECT 241.690 945.720 248.670 946.000 ;
        RECT 249.510 945.720 256.490 946.000 ;
        RECT 257.330 945.720 264.310 946.000 ;
        RECT 265.150 945.720 272.130 946.000 ;
        RECT 272.970 945.720 279.950 946.000 ;
        RECT 280.790 945.720 287.770 946.000 ;
        RECT 288.610 945.720 295.590 946.000 ;
        RECT 296.430 945.720 303.410 946.000 ;
        RECT 304.250 945.720 311.230 946.000 ;
        RECT 312.070 945.720 319.050 946.000 ;
        RECT 319.890 945.720 326.870 946.000 ;
        RECT 327.710 945.720 334.690 946.000 ;
        RECT 335.530 945.720 342.510 946.000 ;
        RECT 343.350 945.720 350.330 946.000 ;
        RECT 351.170 945.720 358.150 946.000 ;
        RECT 358.990 945.720 365.970 946.000 ;
        RECT 366.810 945.720 373.790 946.000 ;
        RECT 374.630 945.720 381.610 946.000 ;
        RECT 382.450 945.720 389.430 946.000 ;
        RECT 390.270 945.720 397.250 946.000 ;
        RECT 398.090 945.720 405.070 946.000 ;
        RECT 405.910 945.720 412.890 946.000 ;
        RECT 413.730 945.720 420.710 946.000 ;
        RECT 421.550 945.720 428.530 946.000 ;
        RECT 429.370 945.720 436.350 946.000 ;
        RECT 437.190 945.720 444.170 946.000 ;
        RECT 445.010 945.720 451.990 946.000 ;
        RECT 452.830 945.720 459.810 946.000 ;
        RECT 460.650 945.720 467.630 946.000 ;
        RECT 468.470 945.720 475.450 946.000 ;
        RECT 476.290 945.720 483.270 946.000 ;
        RECT 484.110 945.720 491.090 946.000 ;
        RECT 491.930 945.720 498.910 946.000 ;
        RECT 499.750 945.720 506.730 946.000 ;
        RECT 507.570 945.720 514.550 946.000 ;
        RECT 515.390 945.720 522.370 946.000 ;
        RECT 523.210 945.720 530.190 946.000 ;
        RECT 531.030 945.720 538.010 946.000 ;
        RECT 538.850 945.720 545.830 946.000 ;
        RECT 546.670 945.720 553.650 946.000 ;
        RECT 554.490 945.720 561.470 946.000 ;
        RECT 562.310 945.720 569.290 946.000 ;
        RECT 570.130 945.720 577.110 946.000 ;
        RECT 577.950 945.720 584.930 946.000 ;
        RECT 585.770 945.720 592.750 946.000 ;
        RECT 593.590 945.720 595.610 946.000 ;
        RECT 4.690 4.280 595.610 945.720 ;
        RECT 4.690 3.670 15.450 4.280 ;
        RECT 16.290 3.670 24.190 4.280 ;
        RECT 25.030 3.670 32.930 4.280 ;
        RECT 33.770 3.670 41.670 4.280 ;
        RECT 42.510 3.670 50.410 4.280 ;
        RECT 51.250 3.670 59.150 4.280 ;
        RECT 59.990 3.670 67.890 4.280 ;
        RECT 68.730 3.670 76.630 4.280 ;
        RECT 77.470 3.670 85.370 4.280 ;
        RECT 86.210 3.670 94.110 4.280 ;
        RECT 94.950 3.670 102.850 4.280 ;
        RECT 103.690 3.670 111.590 4.280 ;
        RECT 112.430 3.670 120.330 4.280 ;
        RECT 121.170 3.670 129.070 4.280 ;
        RECT 129.910 3.670 137.810 4.280 ;
        RECT 138.650 3.670 146.550 4.280 ;
        RECT 147.390 3.670 155.290 4.280 ;
        RECT 156.130 3.670 164.030 4.280 ;
        RECT 164.870 3.670 172.770 4.280 ;
        RECT 173.610 3.670 181.510 4.280 ;
        RECT 182.350 3.670 190.250 4.280 ;
        RECT 191.090 3.670 198.990 4.280 ;
        RECT 199.830 3.670 207.730 4.280 ;
        RECT 208.570 3.670 216.470 4.280 ;
        RECT 217.310 3.670 225.210 4.280 ;
        RECT 226.050 3.670 233.950 4.280 ;
        RECT 234.790 3.670 242.690 4.280 ;
        RECT 243.530 3.670 251.430 4.280 ;
        RECT 252.270 3.670 260.170 4.280 ;
        RECT 261.010 3.670 268.910 4.280 ;
        RECT 269.750 3.670 277.650 4.280 ;
        RECT 278.490 3.670 286.390 4.280 ;
        RECT 287.230 3.670 295.130 4.280 ;
        RECT 295.970 3.670 303.870 4.280 ;
        RECT 304.710 3.670 312.610 4.280 ;
        RECT 313.450 3.670 321.350 4.280 ;
        RECT 322.190 3.670 330.090 4.280 ;
        RECT 330.930 3.670 338.830 4.280 ;
        RECT 339.670 3.670 347.570 4.280 ;
        RECT 348.410 3.670 356.310 4.280 ;
        RECT 357.150 3.670 365.050 4.280 ;
        RECT 365.890 3.670 373.790 4.280 ;
        RECT 374.630 3.670 382.530 4.280 ;
        RECT 383.370 3.670 391.270 4.280 ;
        RECT 392.110 3.670 400.010 4.280 ;
        RECT 400.850 3.670 408.750 4.280 ;
        RECT 409.590 3.670 417.490 4.280 ;
        RECT 418.330 3.670 426.230 4.280 ;
        RECT 427.070 3.670 434.970 4.280 ;
        RECT 435.810 3.670 443.710 4.280 ;
        RECT 444.550 3.670 452.450 4.280 ;
        RECT 453.290 3.670 461.190 4.280 ;
        RECT 462.030 3.670 469.930 4.280 ;
        RECT 470.770 3.670 478.670 4.280 ;
        RECT 479.510 3.670 487.410 4.280 ;
        RECT 488.250 3.670 496.150 4.280 ;
        RECT 496.990 3.670 504.890 4.280 ;
        RECT 505.730 3.670 513.630 4.280 ;
        RECT 514.470 3.670 522.370 4.280 ;
        RECT 523.210 3.670 531.110 4.280 ;
        RECT 531.950 3.670 539.850 4.280 ;
        RECT 540.690 3.670 548.590 4.280 ;
        RECT 549.430 3.670 557.330 4.280 ;
        RECT 558.170 3.670 566.070 4.280 ;
        RECT 566.910 3.670 574.810 4.280 ;
        RECT 575.650 3.670 583.550 4.280 ;
        RECT 584.390 3.670 595.610 4.280 ;
      LAYER met3 ;
        RECT 4.000 912.920 596.000 938.565 ;
        RECT 4.400 911.520 596.000 912.920 ;
        RECT 4.000 904.080 596.000 911.520 ;
        RECT 4.400 902.680 596.000 904.080 ;
        RECT 4.000 895.240 596.000 902.680 ;
        RECT 4.400 893.840 596.000 895.240 ;
        RECT 4.000 886.400 596.000 893.840 ;
        RECT 4.400 885.000 596.000 886.400 ;
        RECT 4.000 877.560 596.000 885.000 ;
        RECT 4.400 876.160 596.000 877.560 ;
        RECT 4.000 870.080 596.000 876.160 ;
        RECT 4.000 868.720 595.600 870.080 ;
        RECT 4.400 868.680 595.600 868.720 ;
        RECT 4.400 867.320 596.000 868.680 ;
        RECT 4.000 859.880 596.000 867.320 ;
        RECT 4.400 858.480 596.000 859.880 ;
        RECT 4.000 851.040 596.000 858.480 ;
        RECT 4.400 849.640 596.000 851.040 ;
        RECT 4.000 842.200 596.000 849.640 ;
        RECT 4.400 840.800 596.000 842.200 ;
        RECT 4.000 833.360 596.000 840.800 ;
        RECT 4.400 831.960 596.000 833.360 ;
        RECT 4.000 824.520 596.000 831.960 ;
        RECT 4.400 823.120 596.000 824.520 ;
        RECT 4.000 815.680 596.000 823.120 ;
        RECT 4.400 814.280 596.000 815.680 ;
        RECT 4.000 806.840 596.000 814.280 ;
        RECT 4.400 805.440 596.000 806.840 ;
        RECT 4.000 798.000 596.000 805.440 ;
        RECT 4.400 796.600 596.000 798.000 ;
        RECT 4.000 789.160 596.000 796.600 ;
        RECT 4.400 787.760 596.000 789.160 ;
        RECT 4.000 780.320 596.000 787.760 ;
        RECT 4.400 778.920 596.000 780.320 ;
        RECT 4.000 771.480 596.000 778.920 ;
        RECT 4.400 770.080 596.000 771.480 ;
        RECT 4.000 762.640 596.000 770.080 ;
        RECT 4.400 761.240 596.000 762.640 ;
        RECT 4.000 753.800 596.000 761.240 ;
        RECT 4.400 752.400 596.000 753.800 ;
        RECT 4.000 744.960 596.000 752.400 ;
        RECT 4.400 743.560 596.000 744.960 ;
        RECT 4.000 736.120 596.000 743.560 ;
        RECT 4.400 734.720 596.000 736.120 ;
        RECT 4.000 727.280 596.000 734.720 ;
        RECT 4.400 725.880 596.000 727.280 ;
        RECT 4.000 718.440 596.000 725.880 ;
        RECT 4.400 717.040 596.000 718.440 ;
        RECT 4.000 712.320 596.000 717.040 ;
        RECT 4.000 710.920 595.600 712.320 ;
        RECT 4.000 709.600 596.000 710.920 ;
        RECT 4.400 708.200 596.000 709.600 ;
        RECT 4.000 700.760 596.000 708.200 ;
        RECT 4.400 699.360 596.000 700.760 ;
        RECT 4.000 691.920 596.000 699.360 ;
        RECT 4.400 690.520 596.000 691.920 ;
        RECT 4.000 683.080 596.000 690.520 ;
        RECT 4.400 681.680 596.000 683.080 ;
        RECT 4.000 674.240 596.000 681.680 ;
        RECT 4.400 672.840 596.000 674.240 ;
        RECT 4.000 665.400 596.000 672.840 ;
        RECT 4.400 664.000 596.000 665.400 ;
        RECT 4.000 656.560 596.000 664.000 ;
        RECT 4.400 655.160 596.000 656.560 ;
        RECT 4.000 647.720 596.000 655.160 ;
        RECT 4.400 646.320 596.000 647.720 ;
        RECT 4.000 638.880 596.000 646.320 ;
        RECT 4.400 637.480 596.000 638.880 ;
        RECT 4.000 630.040 596.000 637.480 ;
        RECT 4.400 628.640 596.000 630.040 ;
        RECT 4.000 621.200 596.000 628.640 ;
        RECT 4.400 619.800 596.000 621.200 ;
        RECT 4.000 612.360 596.000 619.800 ;
        RECT 4.400 610.960 596.000 612.360 ;
        RECT 4.000 603.520 596.000 610.960 ;
        RECT 4.400 602.120 596.000 603.520 ;
        RECT 4.000 594.680 596.000 602.120 ;
        RECT 4.400 593.280 596.000 594.680 ;
        RECT 4.000 585.840 596.000 593.280 ;
        RECT 4.400 584.440 596.000 585.840 ;
        RECT 4.000 577.000 596.000 584.440 ;
        RECT 4.400 575.600 596.000 577.000 ;
        RECT 4.000 568.160 596.000 575.600 ;
        RECT 4.400 566.760 596.000 568.160 ;
        RECT 4.000 559.320 596.000 566.760 ;
        RECT 4.400 557.920 596.000 559.320 ;
        RECT 4.000 554.560 596.000 557.920 ;
        RECT 4.000 553.160 595.600 554.560 ;
        RECT 4.000 550.480 596.000 553.160 ;
        RECT 4.400 549.080 596.000 550.480 ;
        RECT 4.000 541.640 596.000 549.080 ;
        RECT 4.400 540.240 596.000 541.640 ;
        RECT 4.000 532.800 596.000 540.240 ;
        RECT 4.400 531.400 596.000 532.800 ;
        RECT 4.000 523.960 596.000 531.400 ;
        RECT 4.400 522.560 596.000 523.960 ;
        RECT 4.000 515.120 596.000 522.560 ;
        RECT 4.400 513.720 596.000 515.120 ;
        RECT 4.000 506.280 596.000 513.720 ;
        RECT 4.400 504.880 596.000 506.280 ;
        RECT 4.000 497.440 596.000 504.880 ;
        RECT 4.400 496.040 596.000 497.440 ;
        RECT 4.000 488.600 596.000 496.040 ;
        RECT 4.400 487.200 596.000 488.600 ;
        RECT 4.000 479.760 596.000 487.200 ;
        RECT 4.400 478.360 596.000 479.760 ;
        RECT 4.000 470.920 596.000 478.360 ;
        RECT 4.400 469.520 596.000 470.920 ;
        RECT 4.000 462.080 596.000 469.520 ;
        RECT 4.400 460.680 596.000 462.080 ;
        RECT 4.000 453.240 596.000 460.680 ;
        RECT 4.400 451.840 596.000 453.240 ;
        RECT 4.000 444.400 596.000 451.840 ;
        RECT 4.400 443.000 596.000 444.400 ;
        RECT 4.000 435.560 596.000 443.000 ;
        RECT 4.400 434.160 596.000 435.560 ;
        RECT 4.000 426.720 596.000 434.160 ;
        RECT 4.400 425.320 596.000 426.720 ;
        RECT 4.000 417.880 596.000 425.320 ;
        RECT 4.400 416.480 596.000 417.880 ;
        RECT 4.000 409.040 596.000 416.480 ;
        RECT 4.400 407.640 596.000 409.040 ;
        RECT 4.000 400.200 596.000 407.640 ;
        RECT 4.400 398.800 596.000 400.200 ;
        RECT 4.000 396.800 596.000 398.800 ;
        RECT 4.000 395.400 595.600 396.800 ;
        RECT 4.000 391.360 596.000 395.400 ;
        RECT 4.400 389.960 596.000 391.360 ;
        RECT 4.000 382.520 596.000 389.960 ;
        RECT 4.400 381.120 596.000 382.520 ;
        RECT 4.000 373.680 596.000 381.120 ;
        RECT 4.400 372.280 596.000 373.680 ;
        RECT 4.000 364.840 596.000 372.280 ;
        RECT 4.400 363.440 596.000 364.840 ;
        RECT 4.000 356.000 596.000 363.440 ;
        RECT 4.400 354.600 596.000 356.000 ;
        RECT 4.000 347.160 596.000 354.600 ;
        RECT 4.400 345.760 596.000 347.160 ;
        RECT 4.000 338.320 596.000 345.760 ;
        RECT 4.400 336.920 596.000 338.320 ;
        RECT 4.000 329.480 596.000 336.920 ;
        RECT 4.400 328.080 596.000 329.480 ;
        RECT 4.000 320.640 596.000 328.080 ;
        RECT 4.400 319.240 596.000 320.640 ;
        RECT 4.000 311.800 596.000 319.240 ;
        RECT 4.400 310.400 596.000 311.800 ;
        RECT 4.000 302.960 596.000 310.400 ;
        RECT 4.400 301.560 596.000 302.960 ;
        RECT 4.000 294.120 596.000 301.560 ;
        RECT 4.400 292.720 596.000 294.120 ;
        RECT 4.000 285.280 596.000 292.720 ;
        RECT 4.400 283.880 596.000 285.280 ;
        RECT 4.000 276.440 596.000 283.880 ;
        RECT 4.400 275.040 596.000 276.440 ;
        RECT 4.000 267.600 596.000 275.040 ;
        RECT 4.400 266.200 596.000 267.600 ;
        RECT 4.000 258.760 596.000 266.200 ;
        RECT 4.400 257.360 596.000 258.760 ;
        RECT 4.000 249.920 596.000 257.360 ;
        RECT 4.400 248.520 596.000 249.920 ;
        RECT 4.000 241.080 596.000 248.520 ;
        RECT 4.400 239.680 596.000 241.080 ;
        RECT 4.000 239.040 596.000 239.680 ;
        RECT 4.000 237.640 595.600 239.040 ;
        RECT 4.000 232.240 596.000 237.640 ;
        RECT 4.400 230.840 596.000 232.240 ;
        RECT 4.000 223.400 596.000 230.840 ;
        RECT 4.400 222.000 596.000 223.400 ;
        RECT 4.000 214.560 596.000 222.000 ;
        RECT 4.400 213.160 596.000 214.560 ;
        RECT 4.000 205.720 596.000 213.160 ;
        RECT 4.400 204.320 596.000 205.720 ;
        RECT 4.000 196.880 596.000 204.320 ;
        RECT 4.400 195.480 596.000 196.880 ;
        RECT 4.000 188.040 596.000 195.480 ;
        RECT 4.400 186.640 596.000 188.040 ;
        RECT 4.000 179.200 596.000 186.640 ;
        RECT 4.400 177.800 596.000 179.200 ;
        RECT 4.000 170.360 596.000 177.800 ;
        RECT 4.400 168.960 596.000 170.360 ;
        RECT 4.000 161.520 596.000 168.960 ;
        RECT 4.400 160.120 596.000 161.520 ;
        RECT 4.000 152.680 596.000 160.120 ;
        RECT 4.400 151.280 596.000 152.680 ;
        RECT 4.000 143.840 596.000 151.280 ;
        RECT 4.400 142.440 596.000 143.840 ;
        RECT 4.000 135.000 596.000 142.440 ;
        RECT 4.400 133.600 596.000 135.000 ;
        RECT 4.000 126.160 596.000 133.600 ;
        RECT 4.400 124.760 596.000 126.160 ;
        RECT 4.000 117.320 596.000 124.760 ;
        RECT 4.400 115.920 596.000 117.320 ;
        RECT 4.000 108.480 596.000 115.920 ;
        RECT 4.400 107.080 596.000 108.480 ;
        RECT 4.000 99.640 596.000 107.080 ;
        RECT 4.400 98.240 596.000 99.640 ;
        RECT 4.000 90.800 596.000 98.240 ;
        RECT 4.400 89.400 596.000 90.800 ;
        RECT 4.000 81.960 596.000 89.400 ;
        RECT 4.400 81.280 596.000 81.960 ;
        RECT 4.400 80.560 595.600 81.280 ;
        RECT 4.000 79.880 595.600 80.560 ;
        RECT 4.000 73.120 596.000 79.880 ;
        RECT 4.400 71.720 596.000 73.120 ;
        RECT 4.000 64.280 596.000 71.720 ;
        RECT 4.400 62.880 596.000 64.280 ;
        RECT 4.000 55.440 596.000 62.880 ;
        RECT 4.400 54.040 596.000 55.440 ;
        RECT 4.000 46.600 596.000 54.040 ;
        RECT 4.400 45.200 596.000 46.600 ;
        RECT 4.000 37.760 596.000 45.200 ;
        RECT 4.400 36.360 596.000 37.760 ;
        RECT 4.000 10.715 596.000 36.360 ;
      LAYER met4 ;
        RECT 8.575 11.055 20.640 937.545 ;
        RECT 23.040 11.055 97.440 937.545 ;
        RECT 99.840 11.055 174.240 937.545 ;
        RECT 176.640 11.055 251.040 937.545 ;
        RECT 253.440 11.055 327.840 937.545 ;
        RECT 330.240 11.055 404.640 937.545 ;
        RECT 407.040 11.055 481.440 937.545 ;
        RECT 483.840 11.055 543.425 937.545 ;
  END
END Peripherals
END LIBRARY

