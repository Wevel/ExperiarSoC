VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO IOMultiplexer
  CLASS BLOCK ;
  FOREIGN IOMultiplexer ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END clk
  PIN gpio0_input[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END gpio0_input[0]
  PIN gpio0_input[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END gpio0_input[10]
  PIN gpio0_input[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END gpio0_input[11]
  PIN gpio0_input[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END gpio0_input[12]
  PIN gpio0_input[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END gpio0_input[13]
  PIN gpio0_input[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END gpio0_input[14]
  PIN gpio0_input[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END gpio0_input[15]
  PIN gpio0_input[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END gpio0_input[16]
  PIN gpio0_input[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END gpio0_input[17]
  PIN gpio0_input[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END gpio0_input[18]
  PIN gpio0_input[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END gpio0_input[1]
  PIN gpio0_input[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END gpio0_input[2]
  PIN gpio0_input[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END gpio0_input[3]
  PIN gpio0_input[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END gpio0_input[4]
  PIN gpio0_input[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END gpio0_input[5]
  PIN gpio0_input[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END gpio0_input[6]
  PIN gpio0_input[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END gpio0_input[7]
  PIN gpio0_input[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END gpio0_input[8]
  PIN gpio0_input[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END gpio0_input[9]
  PIN gpio0_oe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END gpio0_oe[0]
  PIN gpio0_oe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END gpio0_oe[10]
  PIN gpio0_oe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END gpio0_oe[11]
  PIN gpio0_oe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END gpio0_oe[12]
  PIN gpio0_oe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END gpio0_oe[13]
  PIN gpio0_oe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END gpio0_oe[14]
  PIN gpio0_oe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END gpio0_oe[15]
  PIN gpio0_oe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END gpio0_oe[16]
  PIN gpio0_oe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END gpio0_oe[17]
  PIN gpio0_oe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END gpio0_oe[18]
  PIN gpio0_oe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END gpio0_oe[1]
  PIN gpio0_oe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END gpio0_oe[2]
  PIN gpio0_oe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END gpio0_oe[3]
  PIN gpio0_oe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END gpio0_oe[4]
  PIN gpio0_oe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END gpio0_oe[5]
  PIN gpio0_oe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END gpio0_oe[6]
  PIN gpio0_oe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END gpio0_oe[7]
  PIN gpio0_oe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END gpio0_oe[8]
  PIN gpio0_oe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END gpio0_oe[9]
  PIN gpio0_output[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END gpio0_output[0]
  PIN gpio0_output[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END gpio0_output[10]
  PIN gpio0_output[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END gpio0_output[11]
  PIN gpio0_output[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END gpio0_output[12]
  PIN gpio0_output[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END gpio0_output[13]
  PIN gpio0_output[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END gpio0_output[14]
  PIN gpio0_output[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END gpio0_output[15]
  PIN gpio0_output[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END gpio0_output[16]
  PIN gpio0_output[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END gpio0_output[17]
  PIN gpio0_output[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END gpio0_output[18]
  PIN gpio0_output[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END gpio0_output[1]
  PIN gpio0_output[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END gpio0_output[2]
  PIN gpio0_output[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END gpio0_output[3]
  PIN gpio0_output[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END gpio0_output[4]
  PIN gpio0_output[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END gpio0_output[5]
  PIN gpio0_output[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END gpio0_output[6]
  PIN gpio0_output[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END gpio0_output[7]
  PIN gpio0_output[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END gpio0_output[8]
  PIN gpio0_output[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END gpio0_output[9]
  PIN gpio1_input[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END gpio1_input[0]
  PIN gpio1_input[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END gpio1_input[10]
  PIN gpio1_input[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END gpio1_input[11]
  PIN gpio1_input[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END gpio1_input[12]
  PIN gpio1_input[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END gpio1_input[13]
  PIN gpio1_input[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END gpio1_input[14]
  PIN gpio1_input[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END gpio1_input[15]
  PIN gpio1_input[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END gpio1_input[16]
  PIN gpio1_input[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END gpio1_input[17]
  PIN gpio1_input[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END gpio1_input[18]
  PIN gpio1_input[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END gpio1_input[1]
  PIN gpio1_input[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END gpio1_input[2]
  PIN gpio1_input[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END gpio1_input[3]
  PIN gpio1_input[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END gpio1_input[4]
  PIN gpio1_input[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END gpio1_input[5]
  PIN gpio1_input[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END gpio1_input[6]
  PIN gpio1_input[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END gpio1_input[7]
  PIN gpio1_input[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END gpio1_input[8]
  PIN gpio1_input[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END gpio1_input[9]
  PIN gpio1_oe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END gpio1_oe[0]
  PIN gpio1_oe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END gpio1_oe[10]
  PIN gpio1_oe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END gpio1_oe[11]
  PIN gpio1_oe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END gpio1_oe[12]
  PIN gpio1_oe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END gpio1_oe[13]
  PIN gpio1_oe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END gpio1_oe[14]
  PIN gpio1_oe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END gpio1_oe[15]
  PIN gpio1_oe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END gpio1_oe[16]
  PIN gpio1_oe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END gpio1_oe[17]
  PIN gpio1_oe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END gpio1_oe[18]
  PIN gpio1_oe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END gpio1_oe[1]
  PIN gpio1_oe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END gpio1_oe[2]
  PIN gpio1_oe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END gpio1_oe[3]
  PIN gpio1_oe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END gpio1_oe[4]
  PIN gpio1_oe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END gpio1_oe[5]
  PIN gpio1_oe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END gpio1_oe[6]
  PIN gpio1_oe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END gpio1_oe[7]
  PIN gpio1_oe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END gpio1_oe[8]
  PIN gpio1_oe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END gpio1_oe[9]
  PIN gpio1_output[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END gpio1_output[0]
  PIN gpio1_output[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END gpio1_output[10]
  PIN gpio1_output[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END gpio1_output[11]
  PIN gpio1_output[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END gpio1_output[12]
  PIN gpio1_output[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END gpio1_output[13]
  PIN gpio1_output[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END gpio1_output[14]
  PIN gpio1_output[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END gpio1_output[15]
  PIN gpio1_output[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END gpio1_output[16]
  PIN gpio1_output[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END gpio1_output[17]
  PIN gpio1_output[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END gpio1_output[18]
  PIN gpio1_output[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END gpio1_output[1]
  PIN gpio1_output[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END gpio1_output[2]
  PIN gpio1_output[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END gpio1_output[3]
  PIN gpio1_output[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END gpio1_output[4]
  PIN gpio1_output[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END gpio1_output[5]
  PIN gpio1_output[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END gpio1_output[6]
  PIN gpio1_output[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END gpio1_output[7]
  PIN gpio1_output[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END gpio1_output[8]
  PIN gpio1_output[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END gpio1_output[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 196.000 0.830 200.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 196.000 53.270 200.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 196.000 58.330 200.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 196.000 63.850 200.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 196.000 68.910 200.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 196.000 74.430 200.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 196.000 79.490 200.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 196.000 85.010 200.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 196.000 90.070 200.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 196.000 95.590 200.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 196.000 100.650 200.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 196.000 5.890 200.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 196.000 105.710 200.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 196.000 111.230 200.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 196.000 116.290 200.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 196.000 121.810 200.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 196.000 126.870 200.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 196.000 132.390 200.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 196.000 137.450 200.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 196.000 142.970 200.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 196.000 148.030 200.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 196.000 153.090 200.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 196.000 10.950 200.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 196.000 158.610 200.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 196.000 163.670 200.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 196.000 169.190 200.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 196.000 174.250 200.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 196.000 179.770 200.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 196.000 184.830 200.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 196.000 190.350 200.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 196.000 195.410 200.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 196.000 16.470 200.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 196.000 21.530 200.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 196.000 27.050 200.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 196.000 32.110 200.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 196.000 37.630 200.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 196.000 42.690 200.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 196.000 48.210 200.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 196.000 2.210 200.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 196.000 55.110 200.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 196.000 60.170 200.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 196.000 65.690 200.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 196.000 70.750 200.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 196.000 76.270 200.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 196.000 81.330 200.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 196.000 86.390 200.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 196.000 91.910 200.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 196.000 96.970 200.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 196.000 102.490 200.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 196.000 7.730 200.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 196.000 107.550 200.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 196.000 113.070 200.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 196.000 118.130 200.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 196.000 123.650 200.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 196.000 128.710 200.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 196.000 134.230 200.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 196.000 139.290 200.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 196.000 144.350 200.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 196.000 149.870 200.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 196.000 154.930 200.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 196.000 12.790 200.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 196.000 160.450 200.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 196.000 165.510 200.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 196.000 171.030 200.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 196.000 176.090 200.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 196.000 181.610 200.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 196.000 186.670 200.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 196.000 191.730 200.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 196.000 197.250 200.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 196.000 18.310 200.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 196.000 23.370 200.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 196.000 28.890 200.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 196.000 33.950 200.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 196.000 39.010 200.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 196.000 44.530 200.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 196.000 49.590 200.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 196.000 4.050 200.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 196.000 56.950 200.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 196.000 62.010 200.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 196.000 67.530 200.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 196.000 72.590 200.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 196.000 77.650 200.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 196.000 83.170 200.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 196.000 88.230 200.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 196.000 93.750 200.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 196.000 98.810 200.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 196.000 104.330 200.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 196.000 9.570 200.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 196.000 109.390 200.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 196.000 114.910 200.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 196.000 119.970 200.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 196.000 125.030 200.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 196.000 130.550 200.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 196.000 135.610 200.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 196.000 141.130 200.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 196.000 146.190 200.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 196.000 151.710 200.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 196.000 156.770 200.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 196.000 14.630 200.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 196.000 162.290 200.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 196.000 167.350 200.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 196.000 172.410 200.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 196.000 177.930 200.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 196.000 182.990 200.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 196.000 188.510 200.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 196.000 193.570 200.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 196.000 199.090 200.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 196.000 19.690 200.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 196.000 25.210 200.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 196.000 30.270 200.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 196.000 35.790 200.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 196.000 40.850 200.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 196.000 46.370 200.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 196.000 51.430 200.000 ;
    END
  END io_out[9]
  PIN la_blink[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 187.040 200.000 187.640 ;
    END
  END la_blink[0]
  PIN la_blink[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 195.200 200.000 195.800 ;
    END
  END la_blink[1]
  PIN pwm_en[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 4.000 ;
    END
  END pwm_en[0]
  PIN pwm_en[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END pwm_en[10]
  PIN pwm_en[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END pwm_en[11]
  PIN pwm_en[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END pwm_en[12]
  PIN pwm_en[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END pwm_en[13]
  PIN pwm_en[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END pwm_en[14]
  PIN pwm_en[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END pwm_en[15]
  PIN pwm_en[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END pwm_en[1]
  PIN pwm_en[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END pwm_en[2]
  PIN pwm_en[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END pwm_en[3]
  PIN pwm_en[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END pwm_en[4]
  PIN pwm_en[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END pwm_en[5]
  PIN pwm_en[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END pwm_en[6]
  PIN pwm_en[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END pwm_en[7]
  PIN pwm_en[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END pwm_en[8]
  PIN pwm_en[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END pwm_en[9]
  PIN pwm_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END pwm_out[0]
  PIN pwm_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END pwm_out[10]
  PIN pwm_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END pwm_out[11]
  PIN pwm_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END pwm_out[12]
  PIN pwm_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END pwm_out[13]
  PIN pwm_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END pwm_out[14]
  PIN pwm_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END pwm_out[15]
  PIN pwm_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END pwm_out[1]
  PIN pwm_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END pwm_out[2]
  PIN pwm_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END pwm_out[3]
  PIN pwm_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END pwm_out[4]
  PIN pwm_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END pwm_out[5]
  PIN pwm_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END pwm_out[6]
  PIN pwm_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END pwm_out[7]
  PIN pwm_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END pwm_out[8]
  PIN pwm_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END pwm_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END rst
  PIN spi_clk[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 104.080 200.000 104.680 ;
    END
  END spi_clk[0]
  PIN spi_clk[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 145.560 200.000 146.160 ;
    END
  END spi_clk[1]
  PIN spi_cs[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 112.240 200.000 112.840 ;
    END
  END spi_cs[0]
  PIN spi_cs[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 153.720 200.000 154.320 ;
    END
  END spi_cs[1]
  PIN spi_en[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 120.400 200.000 121.000 ;
    END
  END spi_en[0]
  PIN spi_en[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 161.880 200.000 162.480 ;
    END
  END spi_en[1]
  PIN spi_miso[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 128.560 200.000 129.160 ;
    END
  END spi_miso[0]
  PIN spi_miso[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 170.720 200.000 171.320 ;
    END
  END spi_miso[1]
  PIN spi_mosi[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 137.400 200.000 138.000 ;
    END
  END spi_mosi[0]
  PIN spi_mosi[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 178.880 200.000 179.480 ;
    END
  END spi_mosi[1]
  PIN uart_en[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 4.120 200.000 4.720 ;
    END
  END uart_en[0]
  PIN uart_en[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 28.600 200.000 29.200 ;
    END
  END uart_en[1]
  PIN uart_en[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 53.760 200.000 54.360 ;
    END
  END uart_en[2]
  PIN uart_en[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 78.920 200.000 79.520 ;
    END
  END uart_en[3]
  PIN uart_rx[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 12.280 200.000 12.880 ;
    END
  END uart_rx[0]
  PIN uart_rx[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 37.440 200.000 38.040 ;
    END
  END uart_rx[1]
  PIN uart_rx[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 61.920 200.000 62.520 ;
    END
  END uart_rx[2]
  PIN uart_rx[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 87.080 200.000 87.680 ;
    END
  END uart_rx[3]
  PIN uart_tx[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 20.440 200.000 21.040 ;
    END
  END uart_tx[0]
  PIN uart_tx[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 45.600 200.000 46.200 ;
    END
  END uart_tx[1]
  PIN uart_tx[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 70.760 200.000 71.360 ;
    END
  END uart_tx[2]
  PIN uart_tx[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 95.240 200.000 95.840 ;
    END
  END uart_tx[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 0.530 8.540 199.570 189.340 ;
      LAYER met2 ;
        RECT 1.110 195.720 1.650 196.250 ;
        RECT 2.490 195.720 3.490 196.250 ;
        RECT 4.330 195.720 5.330 196.250 ;
        RECT 6.170 195.720 7.170 196.250 ;
        RECT 8.010 195.720 9.010 196.250 ;
        RECT 9.850 195.720 10.390 196.250 ;
        RECT 11.230 195.720 12.230 196.250 ;
        RECT 13.070 195.720 14.070 196.250 ;
        RECT 14.910 195.720 15.910 196.250 ;
        RECT 16.750 195.720 17.750 196.250 ;
        RECT 18.590 195.720 19.130 196.250 ;
        RECT 19.970 195.720 20.970 196.250 ;
        RECT 21.810 195.720 22.810 196.250 ;
        RECT 23.650 195.720 24.650 196.250 ;
        RECT 25.490 195.720 26.490 196.250 ;
        RECT 27.330 195.720 28.330 196.250 ;
        RECT 29.170 195.720 29.710 196.250 ;
        RECT 30.550 195.720 31.550 196.250 ;
        RECT 32.390 195.720 33.390 196.250 ;
        RECT 34.230 195.720 35.230 196.250 ;
        RECT 36.070 195.720 37.070 196.250 ;
        RECT 37.910 195.720 38.450 196.250 ;
        RECT 39.290 195.720 40.290 196.250 ;
        RECT 41.130 195.720 42.130 196.250 ;
        RECT 42.970 195.720 43.970 196.250 ;
        RECT 44.810 195.720 45.810 196.250 ;
        RECT 46.650 195.720 47.650 196.250 ;
        RECT 48.490 195.720 49.030 196.250 ;
        RECT 49.870 195.720 50.870 196.250 ;
        RECT 51.710 195.720 52.710 196.250 ;
        RECT 53.550 195.720 54.550 196.250 ;
        RECT 55.390 195.720 56.390 196.250 ;
        RECT 57.230 195.720 57.770 196.250 ;
        RECT 58.610 195.720 59.610 196.250 ;
        RECT 60.450 195.720 61.450 196.250 ;
        RECT 62.290 195.720 63.290 196.250 ;
        RECT 64.130 195.720 65.130 196.250 ;
        RECT 65.970 195.720 66.970 196.250 ;
        RECT 67.810 195.720 68.350 196.250 ;
        RECT 69.190 195.720 70.190 196.250 ;
        RECT 71.030 195.720 72.030 196.250 ;
        RECT 72.870 195.720 73.870 196.250 ;
        RECT 74.710 195.720 75.710 196.250 ;
        RECT 76.550 195.720 77.090 196.250 ;
        RECT 77.930 195.720 78.930 196.250 ;
        RECT 79.770 195.720 80.770 196.250 ;
        RECT 81.610 195.720 82.610 196.250 ;
        RECT 83.450 195.720 84.450 196.250 ;
        RECT 85.290 195.720 85.830 196.250 ;
        RECT 86.670 195.720 87.670 196.250 ;
        RECT 88.510 195.720 89.510 196.250 ;
        RECT 90.350 195.720 91.350 196.250 ;
        RECT 92.190 195.720 93.190 196.250 ;
        RECT 94.030 195.720 95.030 196.250 ;
        RECT 95.870 195.720 96.410 196.250 ;
        RECT 97.250 195.720 98.250 196.250 ;
        RECT 99.090 195.720 100.090 196.250 ;
        RECT 100.930 195.720 101.930 196.250 ;
        RECT 102.770 195.720 103.770 196.250 ;
        RECT 104.610 195.720 105.150 196.250 ;
        RECT 105.990 195.720 106.990 196.250 ;
        RECT 107.830 195.720 108.830 196.250 ;
        RECT 109.670 195.720 110.670 196.250 ;
        RECT 111.510 195.720 112.510 196.250 ;
        RECT 113.350 195.720 114.350 196.250 ;
        RECT 115.190 195.720 115.730 196.250 ;
        RECT 116.570 195.720 117.570 196.250 ;
        RECT 118.410 195.720 119.410 196.250 ;
        RECT 120.250 195.720 121.250 196.250 ;
        RECT 122.090 195.720 123.090 196.250 ;
        RECT 123.930 195.720 124.470 196.250 ;
        RECT 125.310 195.720 126.310 196.250 ;
        RECT 127.150 195.720 128.150 196.250 ;
        RECT 128.990 195.720 129.990 196.250 ;
        RECT 130.830 195.720 131.830 196.250 ;
        RECT 132.670 195.720 133.670 196.250 ;
        RECT 134.510 195.720 135.050 196.250 ;
        RECT 135.890 195.720 136.890 196.250 ;
        RECT 137.730 195.720 138.730 196.250 ;
        RECT 139.570 195.720 140.570 196.250 ;
        RECT 141.410 195.720 142.410 196.250 ;
        RECT 143.250 195.720 143.790 196.250 ;
        RECT 144.630 195.720 145.630 196.250 ;
        RECT 146.470 195.720 147.470 196.250 ;
        RECT 148.310 195.720 149.310 196.250 ;
        RECT 150.150 195.720 151.150 196.250 ;
        RECT 151.990 195.720 152.530 196.250 ;
        RECT 153.370 195.720 154.370 196.250 ;
        RECT 155.210 195.720 156.210 196.250 ;
        RECT 157.050 195.720 158.050 196.250 ;
        RECT 158.890 195.720 159.890 196.250 ;
        RECT 160.730 195.720 161.730 196.250 ;
        RECT 162.570 195.720 163.110 196.250 ;
        RECT 163.950 195.720 164.950 196.250 ;
        RECT 165.790 195.720 166.790 196.250 ;
        RECT 167.630 195.720 168.630 196.250 ;
        RECT 169.470 195.720 170.470 196.250 ;
        RECT 171.310 195.720 171.850 196.250 ;
        RECT 172.690 195.720 173.690 196.250 ;
        RECT 174.530 195.720 175.530 196.250 ;
        RECT 176.370 195.720 177.370 196.250 ;
        RECT 178.210 195.720 179.210 196.250 ;
        RECT 180.050 195.720 181.050 196.250 ;
        RECT 181.890 195.720 182.430 196.250 ;
        RECT 183.270 195.720 184.270 196.250 ;
        RECT 185.110 195.720 186.110 196.250 ;
        RECT 186.950 195.720 187.950 196.250 ;
        RECT 188.790 195.720 189.790 196.250 ;
        RECT 190.630 195.720 191.170 196.250 ;
        RECT 192.010 195.720 193.010 196.250 ;
        RECT 193.850 195.720 194.850 196.250 ;
        RECT 195.690 195.720 196.690 196.250 ;
        RECT 197.530 195.720 198.530 196.250 ;
        RECT 199.370 195.720 199.540 196.250 ;
        RECT 0.560 4.280 199.540 195.720 ;
        RECT 1.110 4.000 1.190 4.280 ;
        RECT 2.030 4.000 2.570 4.280 ;
        RECT 3.410 4.000 3.950 4.280 ;
        RECT 4.790 4.000 5.330 4.280 ;
        RECT 6.170 4.000 6.710 4.280 ;
        RECT 7.550 4.000 8.090 4.280 ;
        RECT 8.930 4.000 9.470 4.280 ;
        RECT 10.310 4.000 10.850 4.280 ;
        RECT 11.690 4.000 12.230 4.280 ;
        RECT 13.070 4.000 13.610 4.280 ;
        RECT 14.450 4.000 14.990 4.280 ;
        RECT 15.830 4.000 16.370 4.280 ;
        RECT 17.210 4.000 17.750 4.280 ;
        RECT 18.590 4.000 19.130 4.280 ;
        RECT 19.970 4.000 20.510 4.280 ;
        RECT 21.350 4.000 21.890 4.280 ;
        RECT 22.730 4.000 23.270 4.280 ;
        RECT 24.110 4.000 24.650 4.280 ;
        RECT 25.490 4.000 26.030 4.280 ;
        RECT 26.870 4.000 27.410 4.280 ;
        RECT 28.250 4.000 28.790 4.280 ;
        RECT 29.630 4.000 30.170 4.280 ;
        RECT 31.010 4.000 31.550 4.280 ;
        RECT 32.390 4.000 32.930 4.280 ;
        RECT 33.770 4.000 34.310 4.280 ;
        RECT 35.150 4.000 35.690 4.280 ;
        RECT 36.530 4.000 37.070 4.280 ;
        RECT 37.910 4.000 38.450 4.280 ;
        RECT 39.290 4.000 39.830 4.280 ;
        RECT 40.670 4.000 41.210 4.280 ;
        RECT 42.050 4.000 42.590 4.280 ;
        RECT 43.430 4.000 43.970 4.280 ;
        RECT 44.810 4.000 45.350 4.280 ;
        RECT 46.190 4.000 46.730 4.280 ;
        RECT 47.570 4.000 48.110 4.280 ;
        RECT 48.950 4.000 49.490 4.280 ;
        RECT 50.330 4.000 50.870 4.280 ;
        RECT 51.710 4.000 52.250 4.280 ;
        RECT 53.090 4.000 53.630 4.280 ;
        RECT 54.470 4.000 55.010 4.280 ;
        RECT 55.850 4.000 56.390 4.280 ;
        RECT 57.230 4.000 57.770 4.280 ;
        RECT 58.610 4.000 59.150 4.280 ;
        RECT 59.990 4.000 60.530 4.280 ;
        RECT 61.370 4.000 61.910 4.280 ;
        RECT 62.750 4.000 63.290 4.280 ;
        RECT 64.130 4.000 64.670 4.280 ;
        RECT 65.510 4.000 66.050 4.280 ;
        RECT 66.890 4.000 66.970 4.280 ;
        RECT 67.810 4.000 68.350 4.280 ;
        RECT 69.190 4.000 69.730 4.280 ;
        RECT 70.570 4.000 71.110 4.280 ;
        RECT 71.950 4.000 72.490 4.280 ;
        RECT 73.330 4.000 73.870 4.280 ;
        RECT 74.710 4.000 75.250 4.280 ;
        RECT 76.090 4.000 76.630 4.280 ;
        RECT 77.470 4.000 78.010 4.280 ;
        RECT 78.850 4.000 79.390 4.280 ;
        RECT 80.230 4.000 80.770 4.280 ;
        RECT 81.610 4.000 82.150 4.280 ;
        RECT 82.990 4.000 83.530 4.280 ;
        RECT 84.370 4.000 84.910 4.280 ;
        RECT 85.750 4.000 86.290 4.280 ;
        RECT 87.130 4.000 87.670 4.280 ;
        RECT 88.510 4.000 89.050 4.280 ;
        RECT 89.890 4.000 90.430 4.280 ;
        RECT 91.270 4.000 91.810 4.280 ;
        RECT 92.650 4.000 93.190 4.280 ;
        RECT 94.030 4.000 94.570 4.280 ;
        RECT 95.410 4.000 95.950 4.280 ;
        RECT 96.790 4.000 97.330 4.280 ;
        RECT 98.170 4.000 98.710 4.280 ;
        RECT 99.550 4.000 100.090 4.280 ;
        RECT 100.930 4.000 101.470 4.280 ;
        RECT 102.310 4.000 102.850 4.280 ;
        RECT 103.690 4.000 104.230 4.280 ;
        RECT 105.070 4.000 105.610 4.280 ;
        RECT 106.450 4.000 106.990 4.280 ;
        RECT 107.830 4.000 108.370 4.280 ;
        RECT 109.210 4.000 109.750 4.280 ;
        RECT 110.590 4.000 111.130 4.280 ;
        RECT 111.970 4.000 112.510 4.280 ;
        RECT 113.350 4.000 113.890 4.280 ;
        RECT 114.730 4.000 115.270 4.280 ;
        RECT 116.110 4.000 116.650 4.280 ;
        RECT 117.490 4.000 118.030 4.280 ;
        RECT 118.870 4.000 119.410 4.280 ;
        RECT 120.250 4.000 120.790 4.280 ;
        RECT 121.630 4.000 122.170 4.280 ;
        RECT 123.010 4.000 123.550 4.280 ;
        RECT 124.390 4.000 124.930 4.280 ;
        RECT 125.770 4.000 126.310 4.280 ;
        RECT 127.150 4.000 127.690 4.280 ;
        RECT 128.530 4.000 129.070 4.280 ;
        RECT 129.910 4.000 130.450 4.280 ;
        RECT 131.290 4.000 131.830 4.280 ;
        RECT 132.670 4.000 133.210 4.280 ;
        RECT 134.050 4.000 134.130 4.280 ;
        RECT 134.970 4.000 135.510 4.280 ;
        RECT 136.350 4.000 136.890 4.280 ;
        RECT 137.730 4.000 138.270 4.280 ;
        RECT 139.110 4.000 139.650 4.280 ;
        RECT 140.490 4.000 141.030 4.280 ;
        RECT 141.870 4.000 142.410 4.280 ;
        RECT 143.250 4.000 143.790 4.280 ;
        RECT 144.630 4.000 145.170 4.280 ;
        RECT 146.010 4.000 146.550 4.280 ;
        RECT 147.390 4.000 147.930 4.280 ;
        RECT 148.770 4.000 149.310 4.280 ;
        RECT 150.150 4.000 150.690 4.280 ;
        RECT 151.530 4.000 152.070 4.280 ;
        RECT 152.910 4.000 153.450 4.280 ;
        RECT 154.290 4.000 154.830 4.280 ;
        RECT 155.670 4.000 156.210 4.280 ;
        RECT 157.050 4.000 157.590 4.280 ;
        RECT 158.430 4.000 158.970 4.280 ;
        RECT 159.810 4.000 160.350 4.280 ;
        RECT 161.190 4.000 161.730 4.280 ;
        RECT 162.570 4.000 163.110 4.280 ;
        RECT 163.950 4.000 164.490 4.280 ;
        RECT 165.330 4.000 165.870 4.280 ;
        RECT 166.710 4.000 167.250 4.280 ;
        RECT 168.090 4.000 168.630 4.280 ;
        RECT 169.470 4.000 170.010 4.280 ;
        RECT 170.850 4.000 171.390 4.280 ;
        RECT 172.230 4.000 172.770 4.280 ;
        RECT 173.610 4.000 174.150 4.280 ;
        RECT 174.990 4.000 175.530 4.280 ;
        RECT 176.370 4.000 176.910 4.280 ;
        RECT 177.750 4.000 178.290 4.280 ;
        RECT 179.130 4.000 179.670 4.280 ;
        RECT 180.510 4.000 181.050 4.280 ;
        RECT 181.890 4.000 182.430 4.280 ;
        RECT 183.270 4.000 183.810 4.280 ;
        RECT 184.650 4.000 185.190 4.280 ;
        RECT 186.030 4.000 186.570 4.280 ;
        RECT 187.410 4.000 187.950 4.280 ;
        RECT 188.790 4.000 189.330 4.280 ;
        RECT 190.170 4.000 190.710 4.280 ;
        RECT 191.550 4.000 192.090 4.280 ;
        RECT 192.930 4.000 193.470 4.280 ;
        RECT 194.310 4.000 194.850 4.280 ;
        RECT 195.690 4.000 196.230 4.280 ;
        RECT 197.070 4.000 197.610 4.280 ;
        RECT 198.450 4.000 198.990 4.280 ;
      LAYER met3 ;
        RECT 4.000 194.800 195.600 195.665 ;
        RECT 4.000 188.040 196.000 194.800 ;
        RECT 4.000 186.640 195.600 188.040 ;
        RECT 4.000 179.880 196.000 186.640 ;
        RECT 4.000 178.480 195.600 179.880 ;
        RECT 4.000 171.720 196.000 178.480 ;
        RECT 4.000 170.320 195.600 171.720 ;
        RECT 4.000 162.880 196.000 170.320 ;
        RECT 4.000 161.480 195.600 162.880 ;
        RECT 4.000 154.720 196.000 161.480 ;
        RECT 4.000 153.320 195.600 154.720 ;
        RECT 4.000 150.640 196.000 153.320 ;
        RECT 4.400 149.240 196.000 150.640 ;
        RECT 4.000 146.560 196.000 149.240 ;
        RECT 4.000 145.160 195.600 146.560 ;
        RECT 4.000 138.400 196.000 145.160 ;
        RECT 4.000 137.000 195.600 138.400 ;
        RECT 4.000 129.560 196.000 137.000 ;
        RECT 4.000 128.160 195.600 129.560 ;
        RECT 4.000 121.400 196.000 128.160 ;
        RECT 4.000 120.000 195.600 121.400 ;
        RECT 4.000 113.240 196.000 120.000 ;
        RECT 4.000 111.840 195.600 113.240 ;
        RECT 4.000 105.080 196.000 111.840 ;
        RECT 4.000 103.680 195.600 105.080 ;
        RECT 4.000 96.240 196.000 103.680 ;
        RECT 4.000 94.840 195.600 96.240 ;
        RECT 4.000 88.080 196.000 94.840 ;
        RECT 4.000 86.680 195.600 88.080 ;
        RECT 4.000 79.920 196.000 86.680 ;
        RECT 4.000 78.520 195.600 79.920 ;
        RECT 4.000 71.760 196.000 78.520 ;
        RECT 4.000 70.360 195.600 71.760 ;
        RECT 4.000 62.920 196.000 70.360 ;
        RECT 4.000 61.520 195.600 62.920 ;
        RECT 4.000 54.760 196.000 61.520 ;
        RECT 4.000 53.360 195.600 54.760 ;
        RECT 4.000 50.680 196.000 53.360 ;
        RECT 4.400 49.280 196.000 50.680 ;
        RECT 4.000 46.600 196.000 49.280 ;
        RECT 4.000 45.200 195.600 46.600 ;
        RECT 4.000 38.440 196.000 45.200 ;
        RECT 4.000 37.040 195.600 38.440 ;
        RECT 4.000 29.600 196.000 37.040 ;
        RECT 4.000 28.200 195.600 29.600 ;
        RECT 4.000 21.440 196.000 28.200 ;
        RECT 4.000 20.040 195.600 21.440 ;
        RECT 4.000 13.280 196.000 20.040 ;
        RECT 4.000 11.880 195.600 13.280 ;
        RECT 4.000 5.120 196.000 11.880 ;
        RECT 4.000 4.255 195.600 5.120 ;
  END
END IOMultiplexer
END LIBRARY

