magic
tech sky130A
magscale 1 2
timestamp 1653063340
<< obsli1 >>
rect 1104 2159 118864 137649
<< obsm1 >>
rect 1104 2128 119402 137896
<< metal2 >>
rect 478 139200 534 140000
rect 1490 139200 1546 140000
rect 2502 139200 2558 140000
rect 3606 139200 3662 140000
rect 4618 139200 4674 140000
rect 5722 139200 5778 140000
rect 6734 139200 6790 140000
rect 7838 139200 7894 140000
rect 8850 139200 8906 140000
rect 9862 139200 9918 140000
rect 10966 139200 11022 140000
rect 11978 139200 12034 140000
rect 13082 139200 13138 140000
rect 14094 139200 14150 140000
rect 15198 139200 15254 140000
rect 16210 139200 16266 140000
rect 17314 139200 17370 140000
rect 18326 139200 18382 140000
rect 19338 139200 19394 140000
rect 20442 139200 20498 140000
rect 21454 139200 21510 140000
rect 22558 139200 22614 140000
rect 23570 139200 23626 140000
rect 24674 139200 24730 140000
rect 25686 139200 25742 140000
rect 26698 139200 26754 140000
rect 27802 139200 27858 140000
rect 28814 139200 28870 140000
rect 29918 139200 29974 140000
rect 30930 139200 30986 140000
rect 32034 139200 32090 140000
rect 33046 139200 33102 140000
rect 34150 139200 34206 140000
rect 35162 139200 35218 140000
rect 36174 139200 36230 140000
rect 37278 139200 37334 140000
rect 38290 139200 38346 140000
rect 39394 139200 39450 140000
rect 40406 139200 40462 140000
rect 41510 139200 41566 140000
rect 42522 139200 42578 140000
rect 43534 139200 43590 140000
rect 44638 139200 44694 140000
rect 45650 139200 45706 140000
rect 46754 139200 46810 140000
rect 47766 139200 47822 140000
rect 48870 139200 48926 140000
rect 49882 139200 49938 140000
rect 50986 139200 51042 140000
rect 51998 139200 52054 140000
rect 53010 139200 53066 140000
rect 54114 139200 54170 140000
rect 55126 139200 55182 140000
rect 56230 139200 56286 140000
rect 57242 139200 57298 140000
rect 58346 139200 58402 140000
rect 59358 139200 59414 140000
rect 60462 139200 60518 140000
rect 61474 139200 61530 140000
rect 62486 139200 62542 140000
rect 63590 139200 63646 140000
rect 64602 139200 64658 140000
rect 65706 139200 65762 140000
rect 66718 139200 66774 140000
rect 67822 139200 67878 140000
rect 68834 139200 68890 140000
rect 69846 139200 69902 140000
rect 70950 139200 71006 140000
rect 71962 139200 72018 140000
rect 73066 139200 73122 140000
rect 74078 139200 74134 140000
rect 75182 139200 75238 140000
rect 76194 139200 76250 140000
rect 77298 139200 77354 140000
rect 78310 139200 78366 140000
rect 79322 139200 79378 140000
rect 80426 139200 80482 140000
rect 81438 139200 81494 140000
rect 82542 139200 82598 140000
rect 83554 139200 83610 140000
rect 84658 139200 84714 140000
rect 85670 139200 85726 140000
rect 86682 139200 86738 140000
rect 87786 139200 87842 140000
rect 88798 139200 88854 140000
rect 89902 139200 89958 140000
rect 90914 139200 90970 140000
rect 92018 139200 92074 140000
rect 93030 139200 93086 140000
rect 94134 139200 94190 140000
rect 95146 139200 95202 140000
rect 96158 139200 96214 140000
rect 97262 139200 97318 140000
rect 98274 139200 98330 140000
rect 99378 139200 99434 140000
rect 100390 139200 100446 140000
rect 101494 139200 101550 140000
rect 102506 139200 102562 140000
rect 103518 139200 103574 140000
rect 104622 139200 104678 140000
rect 105634 139200 105690 140000
rect 106738 139200 106794 140000
rect 107750 139200 107806 140000
rect 108854 139200 108910 140000
rect 109866 139200 109922 140000
rect 110970 139200 111026 140000
rect 111982 139200 112038 140000
rect 112994 139200 113050 140000
rect 114098 139200 114154 140000
rect 115110 139200 115166 140000
rect 116214 139200 116270 140000
rect 117226 139200 117282 140000
rect 118330 139200 118386 140000
rect 119342 139200 119398 140000
rect 3330 0 3386 800
rect 9954 0 10010 800
rect 16578 0 16634 800
rect 23294 0 23350 800
rect 29918 0 29974 800
rect 36634 0 36690 800
rect 43258 0 43314 800
rect 49974 0 50030 800
rect 56598 0 56654 800
rect 63314 0 63370 800
rect 69938 0 69994 800
rect 76562 0 76618 800
rect 83278 0 83334 800
rect 89902 0 89958 800
rect 96618 0 96674 800
rect 103242 0 103298 800
rect 109958 0 110014 800
rect 116582 0 116638 800
<< obsm2 >>
rect 1320 139144 1434 139346
rect 1602 139144 2446 139346
rect 2614 139144 3550 139346
rect 3718 139144 4562 139346
rect 4730 139144 5666 139346
rect 5834 139144 6678 139346
rect 6846 139144 7782 139346
rect 7950 139144 8794 139346
rect 8962 139144 9806 139346
rect 9974 139144 10910 139346
rect 11078 139144 11922 139346
rect 12090 139144 13026 139346
rect 13194 139144 14038 139346
rect 14206 139144 15142 139346
rect 15310 139144 16154 139346
rect 16322 139144 17258 139346
rect 17426 139144 18270 139346
rect 18438 139144 19282 139346
rect 19450 139144 20386 139346
rect 20554 139144 21398 139346
rect 21566 139144 22502 139346
rect 22670 139144 23514 139346
rect 23682 139144 24618 139346
rect 24786 139144 25630 139346
rect 25798 139144 26642 139346
rect 26810 139144 27746 139346
rect 27914 139144 28758 139346
rect 28926 139144 29862 139346
rect 30030 139144 30874 139346
rect 31042 139144 31978 139346
rect 32146 139144 32990 139346
rect 33158 139144 34094 139346
rect 34262 139144 35106 139346
rect 35274 139144 36118 139346
rect 36286 139144 37222 139346
rect 37390 139144 38234 139346
rect 38402 139144 39338 139346
rect 39506 139144 40350 139346
rect 40518 139144 41454 139346
rect 41622 139144 42466 139346
rect 42634 139144 43478 139346
rect 43646 139144 44582 139346
rect 44750 139144 45594 139346
rect 45762 139144 46698 139346
rect 46866 139144 47710 139346
rect 47878 139144 48814 139346
rect 48982 139144 49826 139346
rect 49994 139144 50930 139346
rect 51098 139144 51942 139346
rect 52110 139144 52954 139346
rect 53122 139144 54058 139346
rect 54226 139144 55070 139346
rect 55238 139144 56174 139346
rect 56342 139144 57186 139346
rect 57354 139144 58290 139346
rect 58458 139144 59302 139346
rect 59470 139144 60406 139346
rect 60574 139144 61418 139346
rect 61586 139144 62430 139346
rect 62598 139144 63534 139346
rect 63702 139144 64546 139346
rect 64714 139144 65650 139346
rect 65818 139144 66662 139346
rect 66830 139144 67766 139346
rect 67934 139144 68778 139346
rect 68946 139144 69790 139346
rect 69958 139144 70894 139346
rect 71062 139144 71906 139346
rect 72074 139144 73010 139346
rect 73178 139144 74022 139346
rect 74190 139144 75126 139346
rect 75294 139144 76138 139346
rect 76306 139144 77242 139346
rect 77410 139144 78254 139346
rect 78422 139144 79266 139346
rect 79434 139144 80370 139346
rect 80538 139144 81382 139346
rect 81550 139144 82486 139346
rect 82654 139144 83498 139346
rect 83666 139144 84602 139346
rect 84770 139144 85614 139346
rect 85782 139144 86626 139346
rect 86794 139144 87730 139346
rect 87898 139144 88742 139346
rect 88910 139144 89846 139346
rect 90014 139144 90858 139346
rect 91026 139144 91962 139346
rect 92130 139144 92974 139346
rect 93142 139144 94078 139346
rect 94246 139144 95090 139346
rect 95258 139144 96102 139346
rect 96270 139144 97206 139346
rect 97374 139144 98218 139346
rect 98386 139144 99322 139346
rect 99490 139144 100334 139346
rect 100502 139144 101438 139346
rect 101606 139144 102450 139346
rect 102618 139144 103462 139346
rect 103630 139144 104566 139346
rect 104734 139144 105578 139346
rect 105746 139144 106682 139346
rect 106850 139144 107694 139346
rect 107862 139144 108798 139346
rect 108966 139144 109810 139346
rect 109978 139144 110914 139346
rect 111082 139144 111926 139346
rect 112094 139144 112938 139346
rect 113106 139144 114042 139346
rect 114210 139144 115054 139346
rect 115222 139144 116158 139346
rect 116326 139144 117170 139346
rect 117338 139144 118274 139346
rect 118442 139144 119286 139346
rect 1320 856 119396 139144
rect 1320 711 3274 856
rect 3442 711 9898 856
rect 10066 711 16522 856
rect 16690 711 23238 856
rect 23406 711 29862 856
rect 30030 711 36578 856
rect 36746 711 43202 856
rect 43370 711 49918 856
rect 50086 711 56542 856
rect 56710 711 63258 856
rect 63426 711 69882 856
rect 70050 711 76506 856
rect 76674 711 83222 856
rect 83390 711 89846 856
rect 90014 711 96562 856
rect 96730 711 103186 856
rect 103354 711 109902 856
rect 110070 711 116526 856
rect 116694 711 119396 856
<< metal3 >>
rect 0 139136 800 139256
rect 0 137776 800 137896
rect 0 136416 800 136536
rect 0 134920 800 135040
rect 0 133560 800 133680
rect 0 132200 800 132320
rect 0 130704 800 130824
rect 0 129344 800 129464
rect 0 127984 800 128104
rect 119200 128120 120000 128240
rect 0 126624 800 126744
rect 0 125128 800 125248
rect 0 123768 800 123888
rect 0 122408 800 122528
rect 0 120912 800 121032
rect 0 119552 800 119672
rect 0 118192 800 118312
rect 0 116832 800 116952
rect 0 115336 800 115456
rect 0 113976 800 114096
rect 0 112616 800 112736
rect 0 111120 800 111240
rect 0 109760 800 109880
rect 0 108400 800 108520
rect 0 107040 800 107160
rect 0 105544 800 105664
rect 119200 104864 120000 104984
rect 0 104184 800 104304
rect 0 102824 800 102944
rect 0 101328 800 101448
rect 0 99968 800 100088
rect 0 98608 800 98728
rect 0 97248 800 97368
rect 0 95752 800 95872
rect 0 94392 800 94512
rect 0 93032 800 93152
rect 0 91536 800 91656
rect 0 90176 800 90296
rect 0 88816 800 88936
rect 0 87320 800 87440
rect 0 85960 800 86080
rect 0 84600 800 84720
rect 0 83240 800 83360
rect 0 81744 800 81864
rect 119200 81472 120000 81592
rect 0 80384 800 80504
rect 0 79024 800 79144
rect 0 77528 800 77648
rect 0 76168 800 76288
rect 0 74808 800 74928
rect 0 73448 800 73568
rect 0 71952 800 72072
rect 0 70592 800 70712
rect 0 69232 800 69352
rect 0 67736 800 67856
rect 0 66376 800 66496
rect 0 65016 800 65136
rect 0 63656 800 63776
rect 0 62160 800 62280
rect 0 60800 800 60920
rect 0 59440 800 59560
rect 119200 58216 120000 58336
rect 0 57944 800 58064
rect 0 56584 800 56704
rect 0 55224 800 55344
rect 0 53864 800 53984
rect 0 52368 800 52488
rect 0 51008 800 51128
rect 0 49648 800 49768
rect 0 48152 800 48272
rect 0 46792 800 46912
rect 0 45432 800 45552
rect 0 43936 800 44056
rect 0 42576 800 42696
rect 0 41216 800 41336
rect 0 39856 800 39976
rect 0 38360 800 38480
rect 0 37000 800 37120
rect 0 35640 800 35760
rect 119200 34824 120000 34944
rect 0 34144 800 34264
rect 0 32784 800 32904
rect 0 31424 800 31544
rect 0 30064 800 30184
rect 0 28568 800 28688
rect 0 27208 800 27328
rect 0 25848 800 25968
rect 0 24352 800 24472
rect 0 22992 800 23112
rect 0 21632 800 21752
rect 0 20272 800 20392
rect 0 18776 800 18896
rect 0 17416 800 17536
rect 0 16056 800 16176
rect 0 14560 800 14680
rect 0 13200 800 13320
rect 0 11840 800 11960
rect 119200 11568 120000 11688
rect 0 10480 800 10600
rect 0 8984 800 9104
rect 0 7624 800 7744
rect 0 6264 800 6384
rect 0 4768 800 4888
rect 0 3408 800 3528
rect 0 2048 800 2168
rect 0 688 800 808
<< obsm3 >>
rect 880 139056 119200 139229
rect 800 137976 119200 139056
rect 880 137696 119200 137976
rect 800 136616 119200 137696
rect 880 136336 119200 136616
rect 800 135120 119200 136336
rect 880 134840 119200 135120
rect 800 133760 119200 134840
rect 880 133480 119200 133760
rect 800 132400 119200 133480
rect 880 132120 119200 132400
rect 800 130904 119200 132120
rect 880 130624 119200 130904
rect 800 129544 119200 130624
rect 880 129264 119200 129544
rect 800 128320 119200 129264
rect 800 128184 119120 128320
rect 880 128040 119120 128184
rect 880 127904 119200 128040
rect 800 126824 119200 127904
rect 880 126544 119200 126824
rect 800 125328 119200 126544
rect 880 125048 119200 125328
rect 800 123968 119200 125048
rect 880 123688 119200 123968
rect 800 122608 119200 123688
rect 880 122328 119200 122608
rect 800 121112 119200 122328
rect 880 120832 119200 121112
rect 800 119752 119200 120832
rect 880 119472 119200 119752
rect 800 118392 119200 119472
rect 880 118112 119200 118392
rect 800 117032 119200 118112
rect 880 116752 119200 117032
rect 800 115536 119200 116752
rect 880 115256 119200 115536
rect 800 114176 119200 115256
rect 880 113896 119200 114176
rect 800 112816 119200 113896
rect 880 112536 119200 112816
rect 800 111320 119200 112536
rect 880 111040 119200 111320
rect 800 109960 119200 111040
rect 880 109680 119200 109960
rect 800 108600 119200 109680
rect 880 108320 119200 108600
rect 800 107240 119200 108320
rect 880 106960 119200 107240
rect 800 105744 119200 106960
rect 880 105464 119200 105744
rect 800 105064 119200 105464
rect 800 104784 119120 105064
rect 800 104384 119200 104784
rect 880 104104 119200 104384
rect 800 103024 119200 104104
rect 880 102744 119200 103024
rect 800 101528 119200 102744
rect 880 101248 119200 101528
rect 800 100168 119200 101248
rect 880 99888 119200 100168
rect 800 98808 119200 99888
rect 880 98528 119200 98808
rect 800 97448 119200 98528
rect 880 97168 119200 97448
rect 800 95952 119200 97168
rect 880 95672 119200 95952
rect 800 94592 119200 95672
rect 880 94312 119200 94592
rect 800 93232 119200 94312
rect 880 92952 119200 93232
rect 800 91736 119200 92952
rect 880 91456 119200 91736
rect 800 90376 119200 91456
rect 880 90096 119200 90376
rect 800 89016 119200 90096
rect 880 88736 119200 89016
rect 800 87520 119200 88736
rect 880 87240 119200 87520
rect 800 86160 119200 87240
rect 880 85880 119200 86160
rect 800 84800 119200 85880
rect 880 84520 119200 84800
rect 800 83440 119200 84520
rect 880 83160 119200 83440
rect 800 81944 119200 83160
rect 880 81672 119200 81944
rect 880 81664 119120 81672
rect 800 81392 119120 81664
rect 800 80584 119200 81392
rect 880 80304 119200 80584
rect 800 79224 119200 80304
rect 880 78944 119200 79224
rect 800 77728 119200 78944
rect 880 77448 119200 77728
rect 800 76368 119200 77448
rect 880 76088 119200 76368
rect 800 75008 119200 76088
rect 880 74728 119200 75008
rect 800 73648 119200 74728
rect 880 73368 119200 73648
rect 800 72152 119200 73368
rect 880 71872 119200 72152
rect 800 70792 119200 71872
rect 880 70512 119200 70792
rect 800 69432 119200 70512
rect 880 69152 119200 69432
rect 800 67936 119200 69152
rect 880 67656 119200 67936
rect 800 66576 119200 67656
rect 880 66296 119200 66576
rect 800 65216 119200 66296
rect 880 64936 119200 65216
rect 800 63856 119200 64936
rect 880 63576 119200 63856
rect 800 62360 119200 63576
rect 880 62080 119200 62360
rect 800 61000 119200 62080
rect 880 60720 119200 61000
rect 800 59640 119200 60720
rect 880 59360 119200 59640
rect 800 58416 119200 59360
rect 800 58144 119120 58416
rect 880 58136 119120 58144
rect 880 57864 119200 58136
rect 800 56784 119200 57864
rect 880 56504 119200 56784
rect 800 55424 119200 56504
rect 880 55144 119200 55424
rect 800 54064 119200 55144
rect 880 53784 119200 54064
rect 800 52568 119200 53784
rect 880 52288 119200 52568
rect 800 51208 119200 52288
rect 880 50928 119200 51208
rect 800 49848 119200 50928
rect 880 49568 119200 49848
rect 800 48352 119200 49568
rect 880 48072 119200 48352
rect 800 46992 119200 48072
rect 880 46712 119200 46992
rect 800 45632 119200 46712
rect 880 45352 119200 45632
rect 800 44136 119200 45352
rect 880 43856 119200 44136
rect 800 42776 119200 43856
rect 880 42496 119200 42776
rect 800 41416 119200 42496
rect 880 41136 119200 41416
rect 800 40056 119200 41136
rect 880 39776 119200 40056
rect 800 38560 119200 39776
rect 880 38280 119200 38560
rect 800 37200 119200 38280
rect 880 36920 119200 37200
rect 800 35840 119200 36920
rect 880 35560 119200 35840
rect 800 35024 119200 35560
rect 800 34744 119120 35024
rect 800 34344 119200 34744
rect 880 34064 119200 34344
rect 800 32984 119200 34064
rect 880 32704 119200 32984
rect 800 31624 119200 32704
rect 880 31344 119200 31624
rect 800 30264 119200 31344
rect 880 29984 119200 30264
rect 800 28768 119200 29984
rect 880 28488 119200 28768
rect 800 27408 119200 28488
rect 880 27128 119200 27408
rect 800 26048 119200 27128
rect 880 25768 119200 26048
rect 800 24552 119200 25768
rect 880 24272 119200 24552
rect 800 23192 119200 24272
rect 880 22912 119200 23192
rect 800 21832 119200 22912
rect 880 21552 119200 21832
rect 800 20472 119200 21552
rect 880 20192 119200 20472
rect 800 18976 119200 20192
rect 880 18696 119200 18976
rect 800 17616 119200 18696
rect 880 17336 119200 17616
rect 800 16256 119200 17336
rect 880 15976 119200 16256
rect 800 14760 119200 15976
rect 880 14480 119200 14760
rect 800 13400 119200 14480
rect 880 13120 119200 13400
rect 800 12040 119200 13120
rect 880 11768 119200 12040
rect 880 11760 119120 11768
rect 800 11488 119120 11760
rect 800 10680 119200 11488
rect 880 10400 119200 10680
rect 800 9184 119200 10400
rect 880 8904 119200 9184
rect 800 7824 119200 8904
rect 880 7544 119200 7824
rect 800 6464 119200 7544
rect 880 6184 119200 6464
rect 800 4968 119200 6184
rect 880 4688 119200 4968
rect 800 3608 119200 4688
rect 880 3328 119200 3608
rect 800 2248 119200 3328
rect 880 1968 119200 2248
rect 800 888 119200 1968
rect 880 715 119200 888
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
rect 111728 2128 112048 137680
<< obsm4 >>
rect 4843 6835 19488 122229
rect 19968 6835 34848 122229
rect 35328 6835 50208 122229
rect 50688 6835 65568 122229
rect 66048 6835 80928 122229
rect 81408 6835 96288 122229
rect 96768 6835 108685 122229
<< labels >>
rlabel metal2 s 16578 0 16634 800 6 flash_csb
port 1 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 flash_io0_read
port 2 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 flash_io0_we
port 3 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 flash_io0_write
port 4 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 flash_io1_read
port 5 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 flash_io1_we
port 6 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 flash_io1_write
port 7 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 flash_sck
port 8 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 internal_uart_rx
port 9 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 internal_uart_tx
port 10 nsew signal output
rlabel metal2 s 478 139200 534 140000 6 io_in[0]
port 11 nsew signal input
rlabel metal2 s 32034 139200 32090 140000 6 io_in[10]
port 12 nsew signal input
rlabel metal2 s 35162 139200 35218 140000 6 io_in[11]
port 13 nsew signal input
rlabel metal2 s 38290 139200 38346 140000 6 io_in[12]
port 14 nsew signal input
rlabel metal2 s 41510 139200 41566 140000 6 io_in[13]
port 15 nsew signal input
rlabel metal2 s 44638 139200 44694 140000 6 io_in[14]
port 16 nsew signal input
rlabel metal2 s 47766 139200 47822 140000 6 io_in[15]
port 17 nsew signal input
rlabel metal2 s 50986 139200 51042 140000 6 io_in[16]
port 18 nsew signal input
rlabel metal2 s 54114 139200 54170 140000 6 io_in[17]
port 19 nsew signal input
rlabel metal2 s 57242 139200 57298 140000 6 io_in[18]
port 20 nsew signal input
rlabel metal2 s 60462 139200 60518 140000 6 io_in[19]
port 21 nsew signal input
rlabel metal2 s 3606 139200 3662 140000 6 io_in[1]
port 22 nsew signal input
rlabel metal2 s 63590 139200 63646 140000 6 io_in[20]
port 23 nsew signal input
rlabel metal2 s 66718 139200 66774 140000 6 io_in[21]
port 24 nsew signal input
rlabel metal2 s 69846 139200 69902 140000 6 io_in[22]
port 25 nsew signal input
rlabel metal2 s 73066 139200 73122 140000 6 io_in[23]
port 26 nsew signal input
rlabel metal2 s 76194 139200 76250 140000 6 io_in[24]
port 27 nsew signal input
rlabel metal2 s 79322 139200 79378 140000 6 io_in[25]
port 28 nsew signal input
rlabel metal2 s 82542 139200 82598 140000 6 io_in[26]
port 29 nsew signal input
rlabel metal2 s 85670 139200 85726 140000 6 io_in[27]
port 30 nsew signal input
rlabel metal2 s 88798 139200 88854 140000 6 io_in[28]
port 31 nsew signal input
rlabel metal2 s 92018 139200 92074 140000 6 io_in[29]
port 32 nsew signal input
rlabel metal2 s 6734 139200 6790 140000 6 io_in[2]
port 33 nsew signal input
rlabel metal2 s 95146 139200 95202 140000 6 io_in[30]
port 34 nsew signal input
rlabel metal2 s 98274 139200 98330 140000 6 io_in[31]
port 35 nsew signal input
rlabel metal2 s 101494 139200 101550 140000 6 io_in[32]
port 36 nsew signal input
rlabel metal2 s 104622 139200 104678 140000 6 io_in[33]
port 37 nsew signal input
rlabel metal2 s 107750 139200 107806 140000 6 io_in[34]
port 38 nsew signal input
rlabel metal2 s 110970 139200 111026 140000 6 io_in[35]
port 39 nsew signal input
rlabel metal2 s 114098 139200 114154 140000 6 io_in[36]
port 40 nsew signal input
rlabel metal2 s 117226 139200 117282 140000 6 io_in[37]
port 41 nsew signal input
rlabel metal2 s 9862 139200 9918 140000 6 io_in[3]
port 42 nsew signal input
rlabel metal2 s 13082 139200 13138 140000 6 io_in[4]
port 43 nsew signal input
rlabel metal2 s 16210 139200 16266 140000 6 io_in[5]
port 44 nsew signal input
rlabel metal2 s 19338 139200 19394 140000 6 io_in[6]
port 45 nsew signal input
rlabel metal2 s 22558 139200 22614 140000 6 io_in[7]
port 46 nsew signal input
rlabel metal2 s 25686 139200 25742 140000 6 io_in[8]
port 47 nsew signal input
rlabel metal2 s 28814 139200 28870 140000 6 io_in[9]
port 48 nsew signal input
rlabel metal2 s 1490 139200 1546 140000 6 io_oeb[0]
port 49 nsew signal output
rlabel metal2 s 33046 139200 33102 140000 6 io_oeb[10]
port 50 nsew signal output
rlabel metal2 s 36174 139200 36230 140000 6 io_oeb[11]
port 51 nsew signal output
rlabel metal2 s 39394 139200 39450 140000 6 io_oeb[12]
port 52 nsew signal output
rlabel metal2 s 42522 139200 42578 140000 6 io_oeb[13]
port 53 nsew signal output
rlabel metal2 s 45650 139200 45706 140000 6 io_oeb[14]
port 54 nsew signal output
rlabel metal2 s 48870 139200 48926 140000 6 io_oeb[15]
port 55 nsew signal output
rlabel metal2 s 51998 139200 52054 140000 6 io_oeb[16]
port 56 nsew signal output
rlabel metal2 s 55126 139200 55182 140000 6 io_oeb[17]
port 57 nsew signal output
rlabel metal2 s 58346 139200 58402 140000 6 io_oeb[18]
port 58 nsew signal output
rlabel metal2 s 61474 139200 61530 140000 6 io_oeb[19]
port 59 nsew signal output
rlabel metal2 s 4618 139200 4674 140000 6 io_oeb[1]
port 60 nsew signal output
rlabel metal2 s 64602 139200 64658 140000 6 io_oeb[20]
port 61 nsew signal output
rlabel metal2 s 67822 139200 67878 140000 6 io_oeb[21]
port 62 nsew signal output
rlabel metal2 s 70950 139200 71006 140000 6 io_oeb[22]
port 63 nsew signal output
rlabel metal2 s 74078 139200 74134 140000 6 io_oeb[23]
port 64 nsew signal output
rlabel metal2 s 77298 139200 77354 140000 6 io_oeb[24]
port 65 nsew signal output
rlabel metal2 s 80426 139200 80482 140000 6 io_oeb[25]
port 66 nsew signal output
rlabel metal2 s 83554 139200 83610 140000 6 io_oeb[26]
port 67 nsew signal output
rlabel metal2 s 86682 139200 86738 140000 6 io_oeb[27]
port 68 nsew signal output
rlabel metal2 s 89902 139200 89958 140000 6 io_oeb[28]
port 69 nsew signal output
rlabel metal2 s 93030 139200 93086 140000 6 io_oeb[29]
port 70 nsew signal output
rlabel metal2 s 7838 139200 7894 140000 6 io_oeb[2]
port 71 nsew signal output
rlabel metal2 s 96158 139200 96214 140000 6 io_oeb[30]
port 72 nsew signal output
rlabel metal2 s 99378 139200 99434 140000 6 io_oeb[31]
port 73 nsew signal output
rlabel metal2 s 102506 139200 102562 140000 6 io_oeb[32]
port 74 nsew signal output
rlabel metal2 s 105634 139200 105690 140000 6 io_oeb[33]
port 75 nsew signal output
rlabel metal2 s 108854 139200 108910 140000 6 io_oeb[34]
port 76 nsew signal output
rlabel metal2 s 111982 139200 112038 140000 6 io_oeb[35]
port 77 nsew signal output
rlabel metal2 s 115110 139200 115166 140000 6 io_oeb[36]
port 78 nsew signal output
rlabel metal2 s 118330 139200 118386 140000 6 io_oeb[37]
port 79 nsew signal output
rlabel metal2 s 10966 139200 11022 140000 6 io_oeb[3]
port 80 nsew signal output
rlabel metal2 s 14094 139200 14150 140000 6 io_oeb[4]
port 81 nsew signal output
rlabel metal2 s 17314 139200 17370 140000 6 io_oeb[5]
port 82 nsew signal output
rlabel metal2 s 20442 139200 20498 140000 6 io_oeb[6]
port 83 nsew signal output
rlabel metal2 s 23570 139200 23626 140000 6 io_oeb[7]
port 84 nsew signal output
rlabel metal2 s 26698 139200 26754 140000 6 io_oeb[8]
port 85 nsew signal output
rlabel metal2 s 29918 139200 29974 140000 6 io_oeb[9]
port 86 nsew signal output
rlabel metal2 s 2502 139200 2558 140000 6 io_out[0]
port 87 nsew signal output
rlabel metal2 s 34150 139200 34206 140000 6 io_out[10]
port 88 nsew signal output
rlabel metal2 s 37278 139200 37334 140000 6 io_out[11]
port 89 nsew signal output
rlabel metal2 s 40406 139200 40462 140000 6 io_out[12]
port 90 nsew signal output
rlabel metal2 s 43534 139200 43590 140000 6 io_out[13]
port 91 nsew signal output
rlabel metal2 s 46754 139200 46810 140000 6 io_out[14]
port 92 nsew signal output
rlabel metal2 s 49882 139200 49938 140000 6 io_out[15]
port 93 nsew signal output
rlabel metal2 s 53010 139200 53066 140000 6 io_out[16]
port 94 nsew signal output
rlabel metal2 s 56230 139200 56286 140000 6 io_out[17]
port 95 nsew signal output
rlabel metal2 s 59358 139200 59414 140000 6 io_out[18]
port 96 nsew signal output
rlabel metal2 s 62486 139200 62542 140000 6 io_out[19]
port 97 nsew signal output
rlabel metal2 s 5722 139200 5778 140000 6 io_out[1]
port 98 nsew signal output
rlabel metal2 s 65706 139200 65762 140000 6 io_out[20]
port 99 nsew signal output
rlabel metal2 s 68834 139200 68890 140000 6 io_out[21]
port 100 nsew signal output
rlabel metal2 s 71962 139200 72018 140000 6 io_out[22]
port 101 nsew signal output
rlabel metal2 s 75182 139200 75238 140000 6 io_out[23]
port 102 nsew signal output
rlabel metal2 s 78310 139200 78366 140000 6 io_out[24]
port 103 nsew signal output
rlabel metal2 s 81438 139200 81494 140000 6 io_out[25]
port 104 nsew signal output
rlabel metal2 s 84658 139200 84714 140000 6 io_out[26]
port 105 nsew signal output
rlabel metal2 s 87786 139200 87842 140000 6 io_out[27]
port 106 nsew signal output
rlabel metal2 s 90914 139200 90970 140000 6 io_out[28]
port 107 nsew signal output
rlabel metal2 s 94134 139200 94190 140000 6 io_out[29]
port 108 nsew signal output
rlabel metal2 s 8850 139200 8906 140000 6 io_out[2]
port 109 nsew signal output
rlabel metal2 s 97262 139200 97318 140000 6 io_out[30]
port 110 nsew signal output
rlabel metal2 s 100390 139200 100446 140000 6 io_out[31]
port 111 nsew signal output
rlabel metal2 s 103518 139200 103574 140000 6 io_out[32]
port 112 nsew signal output
rlabel metal2 s 106738 139200 106794 140000 6 io_out[33]
port 113 nsew signal output
rlabel metal2 s 109866 139200 109922 140000 6 io_out[34]
port 114 nsew signal output
rlabel metal2 s 112994 139200 113050 140000 6 io_out[35]
port 115 nsew signal output
rlabel metal2 s 116214 139200 116270 140000 6 io_out[36]
port 116 nsew signal output
rlabel metal2 s 119342 139200 119398 140000 6 io_out[37]
port 117 nsew signal output
rlabel metal2 s 11978 139200 12034 140000 6 io_out[3]
port 118 nsew signal output
rlabel metal2 s 15198 139200 15254 140000 6 io_out[4]
port 119 nsew signal output
rlabel metal2 s 18326 139200 18382 140000 6 io_out[5]
port 120 nsew signal output
rlabel metal2 s 21454 139200 21510 140000 6 io_out[6]
port 121 nsew signal output
rlabel metal2 s 24674 139200 24730 140000 6 io_out[7]
port 122 nsew signal output
rlabel metal2 s 27802 139200 27858 140000 6 io_out[8]
port 123 nsew signal output
rlabel metal2 s 30930 139200 30986 140000 6 io_out[9]
port 124 nsew signal output
rlabel metal3 s 119200 58216 120000 58336 6 jtag_tck
port 125 nsew signal output
rlabel metal3 s 119200 81472 120000 81592 6 jtag_tdi
port 126 nsew signal output
rlabel metal3 s 119200 104864 120000 104984 6 jtag_tdo
port 127 nsew signal input
rlabel metal3 s 119200 128120 120000 128240 6 jtag_tms
port 128 nsew signal output
rlabel metal3 s 119200 11568 120000 11688 6 probe_blink[0]
port 129 nsew signal output
rlabel metal3 s 119200 34824 120000 34944 6 probe_blink[1]
port 130 nsew signal output
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 131 nsew power bidirectional
rlabel metal2 s 83278 0 83334 800 6 vga_b[0]
port 132 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 vga_b[1]
port 133 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 vga_g[0]
port 134 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 vga_g[1]
port 135 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 vga_hsync
port 136 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 vga_r[0]
port 137 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 vga_r[1]
port 138 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 vga_vsync
port 139 nsew signal input
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 140 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 140 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 140 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 140 nsew ground bidirectional
rlabel metal3 s 0 688 800 808 6 wb_ack_o
port 141 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 wb_adr_i[0]
port 142 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 wb_adr_i[10]
port 143 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 wb_adr_i[11]
port 144 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 wb_adr_i[12]
port 145 nsew signal input
rlabel metal3 s 0 71952 800 72072 6 wb_adr_i[13]
port 146 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 wb_adr_i[14]
port 147 nsew signal input
rlabel metal3 s 0 80384 800 80504 6 wb_adr_i[15]
port 148 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 wb_adr_i[16]
port 149 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 wb_adr_i[17]
port 150 nsew signal input
rlabel metal3 s 0 93032 800 93152 6 wb_adr_i[18]
port 151 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 wb_adr_i[19]
port 152 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 wb_adr_i[1]
port 153 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 wb_adr_i[20]
port 154 nsew signal input
rlabel metal3 s 0 105544 800 105664 6 wb_adr_i[21]
port 155 nsew signal input
rlabel metal3 s 0 109760 800 109880 6 wb_adr_i[22]
port 156 nsew signal input
rlabel metal3 s 0 113976 800 114096 6 wb_adr_i[23]
port 157 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 wb_adr_i[2]
port 158 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 wb_adr_i[3]
port 159 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 wb_adr_i[4]
port 160 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 wb_adr_i[5]
port 161 nsew signal input
rlabel metal3 s 0 42576 800 42696 6 wb_adr_i[6]
port 162 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 wb_adr_i[7]
port 163 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 wb_adr_i[8]
port 164 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 wb_adr_i[9]
port 165 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 wb_clk_i
port 166 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 wb_cyc_i
port 167 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 wb_data_i[0]
port 168 nsew signal input
rlabel metal3 s 0 60800 800 60920 6 wb_data_i[10]
port 169 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 wb_data_i[11]
port 170 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 wb_data_i[12]
port 171 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 wb_data_i[13]
port 172 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 wb_data_i[14]
port 173 nsew signal input
rlabel metal3 s 0 81744 800 81864 6 wb_data_i[15]
port 174 nsew signal input
rlabel metal3 s 0 85960 800 86080 6 wb_data_i[16]
port 175 nsew signal input
rlabel metal3 s 0 90176 800 90296 6 wb_data_i[17]
port 176 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 wb_data_i[18]
port 177 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 wb_data_i[19]
port 178 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 wb_data_i[1]
port 179 nsew signal input
rlabel metal3 s 0 102824 800 102944 6 wb_data_i[20]
port 180 nsew signal input
rlabel metal3 s 0 107040 800 107160 6 wb_data_i[21]
port 181 nsew signal input
rlabel metal3 s 0 111120 800 111240 6 wb_data_i[22]
port 182 nsew signal input
rlabel metal3 s 0 115336 800 115456 6 wb_data_i[23]
port 183 nsew signal input
rlabel metal3 s 0 118192 800 118312 6 wb_data_i[24]
port 184 nsew signal input
rlabel metal3 s 0 120912 800 121032 6 wb_data_i[25]
port 185 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 wb_data_i[26]
port 186 nsew signal input
rlabel metal3 s 0 126624 800 126744 6 wb_data_i[27]
port 187 nsew signal input
rlabel metal3 s 0 129344 800 129464 6 wb_data_i[28]
port 188 nsew signal input
rlabel metal3 s 0 132200 800 132320 6 wb_data_i[29]
port 189 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 wb_data_i[2]
port 190 nsew signal input
rlabel metal3 s 0 134920 800 135040 6 wb_data_i[30]
port 191 nsew signal input
rlabel metal3 s 0 137776 800 137896 6 wb_data_i[31]
port 192 nsew signal input
rlabel metal3 s 0 30064 800 30184 6 wb_data_i[3]
port 193 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 wb_data_i[4]
port 194 nsew signal input
rlabel metal3 s 0 39856 800 39976 6 wb_data_i[5]
port 195 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 wb_data_i[6]
port 196 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 wb_data_i[7]
port 197 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 wb_data_i[8]
port 198 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 wb_data_i[9]
port 199 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 wb_data_o[0]
port 200 nsew signal output
rlabel metal3 s 0 62160 800 62280 6 wb_data_o[10]
port 201 nsew signal output
rlabel metal3 s 0 66376 800 66496 6 wb_data_o[11]
port 202 nsew signal output
rlabel metal3 s 0 70592 800 70712 6 wb_data_o[12]
port 203 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 wb_data_o[13]
port 204 nsew signal output
rlabel metal3 s 0 79024 800 79144 6 wb_data_o[14]
port 205 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 wb_data_o[15]
port 206 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 wb_data_o[16]
port 207 nsew signal output
rlabel metal3 s 0 91536 800 91656 6 wb_data_o[17]
port 208 nsew signal output
rlabel metal3 s 0 95752 800 95872 6 wb_data_o[18]
port 209 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 wb_data_o[19]
port 210 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 wb_data_o[1]
port 211 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 wb_data_o[20]
port 212 nsew signal output
rlabel metal3 s 0 108400 800 108520 6 wb_data_o[21]
port 213 nsew signal output
rlabel metal3 s 0 112616 800 112736 6 wb_data_o[22]
port 214 nsew signal output
rlabel metal3 s 0 116832 800 116952 6 wb_data_o[23]
port 215 nsew signal output
rlabel metal3 s 0 119552 800 119672 6 wb_data_o[24]
port 216 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 wb_data_o[25]
port 217 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 wb_data_o[26]
port 218 nsew signal output
rlabel metal3 s 0 127984 800 128104 6 wb_data_o[27]
port 219 nsew signal output
rlabel metal3 s 0 130704 800 130824 6 wb_data_o[28]
port 220 nsew signal output
rlabel metal3 s 0 133560 800 133680 6 wb_data_o[29]
port 221 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 wb_data_o[2]
port 222 nsew signal output
rlabel metal3 s 0 136416 800 136536 6 wb_data_o[30]
port 223 nsew signal output
rlabel metal3 s 0 139136 800 139256 6 wb_data_o[31]
port 224 nsew signal output
rlabel metal3 s 0 31424 800 31544 6 wb_data_o[3]
port 225 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 wb_data_o[4]
port 226 nsew signal output
rlabel metal3 s 0 41216 800 41336 6 wb_data_o[5]
port 227 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 wb_data_o[6]
port 228 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 wb_data_o[7]
port 229 nsew signal output
rlabel metal3 s 0 53864 800 53984 6 wb_data_o[8]
port 230 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 wb_data_o[9]
port 231 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 wb_error_o
port 232 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 wb_rst_i
port 233 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 wb_sel_i[0]
port 234 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 wb_sel_i[1]
port 235 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 wb_sel_i[2]
port 236 nsew signal input
rlabel metal3 s 0 32784 800 32904 6 wb_sel_i[3]
port 237 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 wb_stall_o
port 238 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 wb_stb_i
port 239 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 wb_we_i
port 240 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 29573842
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripherals_Flat/runs/Peripherals_Flat/results/signoff/Peripherals.magic.gds
string GDS_START 1009082
<< end >>

